library ieee;use ieee.std_logic_1164.all;entity memblock is	port (				clk : in std_logic;				aqa,aqb,aqc,aqd : out std_logic_vector(32*3-1 downto 0);		ada,adb,adc,add : in std_logic_vector(32*3-1 downto 0);		aaa,aab,aac,aad : in std_logic_vector(7*3-1 downto 0);		awa,awb,awc,awd : in std_logic_vector(2 downto 0);				q			: out std_logic_vector(31 downto 0);		d			: in std_logic_vector(31 downto 0);		a			: in std_logic_vector(11 downto 0);		w			: in std_logic	);end entity;architecture memblock_arch of memblock is	component altsyncram		generic (			address_reg_b		: string;			clock_enable_input_a		: string;			clock_enable_input_b		: string;			clock_enable_output_a		: string;			clock_enable_output_b		: string;			indata_reg_b		: string;			intended_device_family		: string;			lpm_type		: string;			numwords_a		: natural;			numwords_b		: natural;			operation_mode		: string;			outdata_aclr_a		: string;			outdata_aclr_b		: string;			outdata_reg_a		: string;			outdata_reg_b		: string;			power_up_uninitialized		: string;			ram_block_type		: string;			read_during_write_mode_mixed_ports		: string;			read_during_write_mode_port_a		: string;			read_during_write_mode_port_b		: string;			widthad_a		: natural;			widthad_b		: natural;			width_a		: natural;			width_b		: natural;			width_byteena_a		: natural;			width_byteena_b		: natural;			wrcontrol_wraddress_reg_b		: string		);		port (			wren_a	: in std_logic ;			clock0	: in std_logic ;			wren_b	: in std_logic ;			address_a : in std_logic_vector (6 downto 0);			address_b : in std_logic_vector (6 downto 0);			q_a	: out std_logic_vector (31 downto 0);			q_b	: out std_logic_vector (31 downto 0);			data_a	: in std_logic_vector (31 downto 0);			data_b	: in std_logic_vector (31 downto 0)		);	end component;		signal bqa,bqb,bqc,bqd : std_logic_vector(32*3-1 downto 0);	signal bda,bdb,bdc,bdd : std_logic_vector(32*3-1 downto 0);	signal baa,bab,bac,bad : std_logic_vector(7*3-1 downto 0);	signal bwa,bwb,bwc,bwd : std_logic_vector(2 downto 0);	beginend memblock_arch;	begin	ax : altsyncram	generic map ("CLOCK0","BYPASS","BYPASS","BYPASS","BYPASS","CLOCK0","Cyclone III","altsyncram",256,256,"BIDIR_DUAL_PORT","NONE","NONE","CLOCK0","CLOCK0","FALSE","M9K","OLD_DATA","OLD_DATA","OLD_DATA",8,8,32,32,1,1,"CLOCK0");	port map (wren_a,clock,wren_b,address_a,		address_b => address_b,		data_a => data_a,		data_b => data_b,		q_a => sub_wire0,		q_b => sub_wire1	);