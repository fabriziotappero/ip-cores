-- ------------------------------------------------------------------------
-- Copyright (C) 2004 Arif Endro Nugroho
-- All rights reserved.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY ARIF ENDRO NUGROHO "AS IS" AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL ARIF ENDRO NUGROHO BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
-- ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
-- 
-- End Of License.
-- ------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity input_fm is
   port (
   clock              : in  bit;
   clear              : in  bit;
   test_signal_fm     : out bit_vector (07 downto 0);
   test_signal_fmTri  : out bit_vector (07 downto 0)
   );
end input_fm;

architecture input_data of input_fm is
component adder_10bit
	port (
	addend_10bit          : in  bit_vector (09 downto 0);
	augend_10bit          : in  bit_vector (09 downto 0);
	adder10_output        : out bit_vector (10 downto 0)
	);
end component;

signal test_signal_fm_int    : bit_vector (07 downto 0);
signal test_signal_fmTri_int : bit_vector (07 downto 0);
signal counter               : bit_vector (09 downto 0);
signal counter_tmp           : bit_vector (10 downto 0);
signal one_increment         : bit_vector (09 downto 0);

begin


    one_increment (00) <= '1';
    one_increment (01) <= '0';
    one_increment (02) <= '0';
    one_increment (03) <= '0';
    one_increment (04) <= '0';
    one_increment (05) <= '0';
    one_increment (06) <= '0';
    one_increment (07) <= '0';
    one_increment (08) <= '0';
    one_increment (09) <= '0';

counter_one : adder_10bit
    port map (
    addend_10bit   => counter,
    augend_10bit   => one_increment,
    adder10_output => counter_tmp
    );
    
process (clock, clear)
begin

    if (clear = '1') then
    		counter              <= (others => '0');
		test_signal_fm       <= (others => '0');
		test_signal_fmTri    <= (others => '0');
    elsif (((clock = '1') and (not( clear = '1'))) and clock'event) then
		counter(09 downto 0) <= counter_tmp(09 downto 0);
		test_signal_fm       <= test_signal_fm_int;
		test_signal_fmTri    <= test_signal_fmTri_int;
    end if;

end process;

	with counter (09 downto 0) select

	test_signal_fm_int <=

-- START INPUT FM SIGNAL

	B"01111111" when B"0000000000",  -- INDEX 0
	B"01110110" when B"0000000001",  -- INDEX 1
	B"01011010" when B"0000000010",  -- INDEX 2
	B"00110000" when B"0000000011",  -- INDEX 3
	B"11111110" when B"0000000100",  -- INDEX 4
	B"11001101" when B"0000000101",  -- INDEX 5
	B"10100011" when B"0000000110",  -- INDEX 6
	B"10001000" when B"0000000111",  -- INDEX 7
	B"10000000" when B"0000001000",  -- INDEX 8
	B"10001100" when B"0000001001",  -- INDEX 9
	B"10101001" when B"0000001010",  -- INDEX 10
	B"11010100" when B"0000001011",  -- INDEX 11
	B"00000110" when B"0000001100",  -- INDEX 12
	B"00110111" when B"0000001101",  -- INDEX 13
	B"01011111" when B"0000001110",  -- INDEX 14
	B"01111001" when B"0000001111",  -- INDEX 15
	B"01111111" when B"0000010000",  -- INDEX 16
	B"01110011" when B"0000010001",  -- INDEX 17
	B"01010100" when B"0000010010",  -- INDEX 18
	B"00101000" when B"0000010011",  -- INDEX 19
	B"11110110" when B"0000010100",  -- INDEX 20
	B"11000101" when B"0000010101",  -- INDEX 21
	B"10011110" when B"0000010110",  -- INDEX 22
	B"10000110" when B"0000010111",  -- INDEX 23
	B"10000001" when B"0000011000",  -- INDEX 24
	B"10001111" when B"0000011001",  -- INDEX 25
	B"10101111" when B"0000011010",  -- INDEX 26
	B"11011100" when B"0000011011",  -- INDEX 27
	B"00001110" when B"0000011100",  -- INDEX 28
	B"00111110" when B"0000011101",  -- INDEX 29
	B"01100101" when B"0000011110",  -- INDEX 30
	B"01111011" when B"0000011111",  -- INDEX 31
	B"01111111" when B"0000100000",  -- INDEX 32
	B"01101111" when B"0000100001",  -- INDEX 33
	B"01001110" when B"0000100010",  -- INDEX 34
	B"00100000" when B"0000100011",  -- INDEX 35
	B"11101110" when B"0000100100",  -- INDEX 36
	B"10111110" when B"0000100101",  -- INDEX 37
	B"10011001" when B"0000100110",  -- INDEX 38
	B"10000100" when B"0000100111",  -- INDEX 39
	B"10000010" when B"0000101000",  -- INDEX 40
	B"10010011" when B"0000101001",  -- INDEX 41
	B"10110110" when B"0000101010",  -- INDEX 42
	B"11100100" when B"0000101011",  -- INDEX 43
	B"00010110" when B"0000101100",  -- INDEX 44
	B"01000101" when B"0000101101",  -- INDEX 45
	B"01101001" when B"0000101110",  -- INDEX 46
	B"01111101" when B"0000101111",  -- INDEX 47
	B"01111110" when B"0000110000",  -- INDEX 48
	B"01101011" when B"0000110001",  -- INDEX 49
	B"01000111" when B"0000110010",  -- INDEX 50
	B"00011000" when B"0000110011",  -- INDEX 51
	B"11100110" when B"0000110100",  -- INDEX 52
	B"10111000" when B"0000110101",  -- INDEX 53
	B"10010100" when B"0000110110",  -- INDEX 54
	B"10000010" when B"0000110111",  -- INDEX 55
	B"10000011" when B"0000111000",  -- INDEX 56
	B"10011000" when B"0000111001",  -- INDEX 57
	B"10111100" when B"0000111010",  -- INDEX 58
	B"11101011" when B"0000111011",  -- INDEX 59
	B"00011110" when B"0000111100",  -- INDEX 60
	B"01001100" when B"0000111101",  -- INDEX 61
	B"01101110" when B"0000111110",  -- INDEX 62
	B"01111111" when B"0000111111",  -- INDEX 63
	B"01111100" when B"0001000000",  -- INDEX 64
	B"01100110" when B"0001000001",  -- INDEX 65
	B"01000000" when B"0001000010",  -- INDEX 66
	B"00010001" when B"0001000011",  -- INDEX 67
	B"11011110" when B"0001000100",  -- INDEX 68
	B"10110001" when B"0001000101",  -- INDEX 69
	B"10010000" when B"0001000110",  -- INDEX 70
	B"10000001" when B"0001000111",  -- INDEX 71
	B"10000101" when B"0001001000",  -- INDEX 72
	B"10011100" when B"0001001001",  -- INDEX 73
	B"11000011" when B"0001001010",  -- INDEX 74
	B"11110011" when B"0001001011",  -- INDEX 75
	B"00100110" when B"0001001100",  -- INDEX 76
	B"01010010" when B"0001001101",  -- INDEX 77
	B"01110010" when B"0001001110",  -- INDEX 78
	B"01111111" when B"0001001111",  -- INDEX 79
	B"01111010" when B"0001010000",  -- INDEX 80
	B"01100001" when B"0001010001",  -- INDEX 81
	B"00111001" when B"0001010010",  -- INDEX 82
	B"00001001" when B"0001010011",  -- INDEX 83
	B"11010111" when B"0001010100",  -- INDEX 84
	B"10101011" when B"0001010101",  -- INDEX 85
	B"10001101" when B"0001010110",  -- INDEX 86
	B"10000000" when B"0001010111",  -- INDEX 87
	B"10001000" when B"0001011000",  -- INDEX 88
	B"10100010" when B"0001011001",  -- INDEX 89
	B"11001010" when B"0001011010",  -- INDEX 90
	B"11111011" when B"0001011011",  -- INDEX 91
	B"00101101" when B"0001011100",  -- INDEX 92
	B"01011000" when B"0001011101",  -- INDEX 93
	B"01110101" when B"0001011110",  -- INDEX 94
	B"01111111" when B"0001011111",  -- INDEX 95
	B"01110111" when B"0001100000",  -- INDEX 96
	B"01011100" when B"0001100001",  -- INDEX 97
	B"00110010" when B"0001100010",  -- INDEX 98
	B"00000001" when B"0001100011",  -- INDEX 99
	B"11001111" when B"0001100100",  -- INDEX 100
	B"10100101" when B"0001100101",  -- INDEX 101
	B"10001001" when B"0001100110",  -- INDEX 102
	B"10000000" when B"0001100111",  -- INDEX 103
	B"10001011" when B"0001101000",  -- INDEX 104
	B"10100111" when B"0001101001",  -- INDEX 105
	B"11010010" when B"0001101010",  -- INDEX 106
	B"00000100" when B"0001101011",  -- INDEX 107
	B"00110101" when B"0001101100",  -- INDEX 108
	B"01011110" when B"0001101101",  -- INDEX 109
	B"01111000" when B"0001101110",  -- INDEX 110
	B"01111111" when B"0001101111",  -- INDEX 111
	B"01110100" when B"0001110000",  -- INDEX 112
	B"01010110" when B"0001110001",  -- INDEX 113
	B"00101010" when B"0001110010",  -- INDEX 114
	B"11111000" when B"0001110011",  -- INDEX 115
	B"11001000" when B"0001110100",  -- INDEX 116
	B"10100000" when B"0001110101",  -- INDEX 117
	B"10000111" when B"0001110110",  -- INDEX 118
	B"10000000" when B"0001110111",  -- INDEX 119
	B"10001110" when B"0001111000",  -- INDEX 120
	B"10101101" when B"0001111001",  -- INDEX 121
	B"11011001" when B"0001111010",  -- INDEX 122
	B"00001100" when B"0001111011",  -- INDEX 123
	B"00111100" when B"0001111100",  -- INDEX 124
	B"01100011" when B"0001111101",  -- INDEX 125
	B"01111011" when B"0001111110",  -- INDEX 126
	B"01111111" when B"0001111111",  -- INDEX 127
	B"01110000" when B"0010000000",  -- INDEX 128
	B"01010000" when B"0010000001",  -- INDEX 129
	B"00100011" when B"0010000010",  -- INDEX 130
	B"11110000" when B"0010000011",  -- INDEX 131
	B"11000001" when B"0010000100",  -- INDEX 132
	B"10011011" when B"0010000101",  -- INDEX 133
	B"10000100" when B"0010000110",  -- INDEX 134
	B"10000001" when B"0010000111",  -- INDEX 135
	B"10010010" when B"0010001000",  -- INDEX 136
	B"10110100" when B"0010001001",  -- INDEX 137
	B"11100001" when B"0010001010",  -- INDEX 138
	B"00010100" when B"0010001011",  -- INDEX 139
	B"01000011" when B"0010001100",  -- INDEX 140
	B"01101000" when B"0010001101",  -- INDEX 141
	B"01111101" when B"0010001110",  -- INDEX 142
	B"01111110" when B"0010001111",  -- INDEX 143
	B"01101100" when B"0010010000",  -- INDEX 144
	B"01001001" when B"0010010001",  -- INDEX 145
	B"00011011" when B"0010010010",  -- INDEX 146
	B"11101001" when B"0010010011",  -- INDEX 147
	B"10111010" when B"0010010100",  -- INDEX 148
	B"10010110" when B"0010010101",  -- INDEX 149
	B"10000010" when B"0010010110",  -- INDEX 150
	B"10000011" when B"0010010111",  -- INDEX 151
	B"10010110" when B"0010011000",  -- INDEX 152
	B"10111010" when B"0010011001",  -- INDEX 153
	B"11101001" when B"0010011010",  -- INDEX 154
	B"00011011" when B"0010011011",  -- INDEX 155
	B"01001010" when B"0010011100",  -- INDEX 156
	B"01101100" when B"0010011101",  -- INDEX 157
	B"01111110" when B"0010011110",  -- INDEX 158
	B"01111101" when B"0010011111",  -- INDEX 159
	B"01101000" when B"0010100000",  -- INDEX 160
	B"01000010" when B"0010100001",  -- INDEX 161
	B"00010011" when B"0010100010",  -- INDEX 162
	B"11100001" when B"0010100011",  -- INDEX 163
	B"10110011" when B"0010100100",  -- INDEX 164
	B"10010010" when B"0010100101",  -- INDEX 165
	B"10000001" when B"0010100110",  -- INDEX 166
	B"10000100" when B"0010100111",  -- INDEX 167
	B"10011011" when B"0010101000",  -- INDEX 168
	B"11000001" when B"0010101001",  -- INDEX 169
	B"11110001" when B"0010101010",  -- INDEX 170
	B"00100011" when B"0010101011",  -- INDEX 171
	B"01010000" when B"0010101100",  -- INDEX 172
	B"01110000" when B"0010101101",  -- INDEX 173
	B"01111111" when B"0010101110",  -- INDEX 174
	B"01111010" when B"0010101111",  -- INDEX 175
	B"01100011" when B"0010110000",  -- INDEX 176
	B"00111011" when B"0010110001",  -- INDEX 177
	B"00001011" when B"0010110010",  -- INDEX 178
	B"11011001" when B"0010110011",  -- INDEX 179
	B"10101101" when B"0010110100",  -- INDEX 180
	B"10001110" when B"0010110101",  -- INDEX 181
	B"10000000" when B"0010110110",  -- INDEX 182
	B"10000111" when B"0010110111",  -- INDEX 183
	B"10100000" when B"0010111000",  -- INDEX 184
	B"11001000" when B"0010111001",  -- INDEX 185
	B"11111001" when B"0010111010",  -- INDEX 186
	B"00101011" when B"0010111011",  -- INDEX 187
	B"01010110" when B"0010111100",  -- INDEX 188
	B"01110100" when B"0010111101",  -- INDEX 189
	B"01111111" when B"0010111110",  -- INDEX 190
	B"01111000" when B"0010111111",  -- INDEX 191
	B"01011101" when B"0011000000",  -- INDEX 192
	B"00110100" when B"0011000001",  -- INDEX 193
	B"00000011" when B"0011000010",  -- INDEX 194
	B"11010001" when B"0011000011",  -- INDEX 195
	B"10100111" when B"0011000100",  -- INDEX 196
	B"10001010" when B"0011000101",  -- INDEX 197
	B"10000000" when B"0011000110",  -- INDEX 198
	B"10001010" when B"0011000111",  -- INDEX 199
	B"10100101" when B"0011001000",  -- INDEX 200
	B"11001111" when B"0011001001",  -- INDEX 201
	B"11111111" when B"0011001010",  -- INDEX 202
	B"00110000" when B"0011001011",  -- INDEX 203
	B"01011001" when B"0011001100",  -- INDEX 204
	B"01110101" when B"0011001101",  -- INDEX 205
	B"01111111" when B"0011001110",  -- INDEX 206
	B"01111000" when B"0011001111",  -- INDEX 207
	B"01011101" when B"0011010000",  -- INDEX 208
	B"00110101" when B"0011010001",  -- INDEX 209
	B"00000101" when B"0011010010",  -- INDEX 210
	B"11010100" when B"0011010011",  -- INDEX 211
	B"10101010" when B"0011010100",  -- INDEX 212
	B"10001100" when B"0011010101",  -- INDEX 213
	B"10000000" when B"0011010110",  -- INDEX 214
	B"10000111" when B"0011010111",  -- INDEX 215
	B"10100000" when B"0011011000",  -- INDEX 216
	B"11000111" when B"0011011001",  -- INDEX 217
	B"11110111" when B"0011011010",  -- INDEX 218
	B"00101000" when B"0011011011",  -- INDEX 219
	B"01010011" when B"0011011100",  -- INDEX 220
	B"01110010" when B"0011011101",  -- INDEX 221
	B"01111111" when B"0011011110",  -- INDEX 222
	B"01111010" when B"0011011111",  -- INDEX 223
	B"01100011" when B"0011100000",  -- INDEX 224
	B"00111100" when B"0011100001",  -- INDEX 225
	B"00001101" when B"0011100010",  -- INDEX 226
	B"11011100" when B"0011100011",  -- INDEX 227
	B"10110000" when B"0011100100",  -- INDEX 228
	B"10010000" when B"0011100101",  -- INDEX 229
	B"10000001" when B"0011100110",  -- INDEX 230
	B"10000101" when B"0011100111",  -- INDEX 231
	B"10011011" when B"0011101000",  -- INDEX 232
	B"11000000" when B"0011101001",  -- INDEX 233
	B"11101111" when B"0011101010",  -- INDEX 234
	B"00100000" when B"0011101011",  -- INDEX 235
	B"01001101" when B"0011101100",  -- INDEX 236
	B"01101110" when B"0011101101",  -- INDEX 237
	B"01111111" when B"0011101110",  -- INDEX 238
	B"01111100" when B"0011101111",  -- INDEX 239
	B"01101000" when B"0011110000",  -- INDEX 240
	B"01000011" when B"0011110001",  -- INDEX 241
	B"00010101" when B"0011110010",  -- INDEX 242
	B"11100100" when B"0011110011",  -- INDEX 243
	B"10110110" when B"0011110100",  -- INDEX 244
	B"10010100" when B"0011110101",  -- INDEX 245
	B"10000010" when B"0011110110",  -- INDEX 246
	B"10000011" when B"0011110111",  -- INDEX 247
	B"10010110" when B"0011111000",  -- INDEX 248
	B"10111001" when B"0011111001",  -- INDEX 249
	B"11100111" when B"0011111010",  -- INDEX 250
	B"00011000" when B"0011111011",  -- INDEX 251
	B"01000110" when B"0011111100",  -- INDEX 252
	B"01101010" when B"0011111101",  -- INDEX 253
	B"01111101" when B"0011111110",  -- INDEX 254
	B"01111110" when B"0011111111",  -- INDEX 255
	B"01101100" when B"0100000000",  -- INDEX 256
	B"01001010" when B"0100000001",  -- INDEX 257
	B"00011101" when B"0100000010",  -- INDEX 258
	B"11101011" when B"0100000011",  -- INDEX 259
	B"10111101" when B"0100000100",  -- INDEX 260
	B"10011001" when B"0100000101",  -- INDEX 261
	B"10000100" when B"0100000110",  -- INDEX 262
	B"10000001" when B"0100000111",  -- INDEX 263
	B"10010010" when B"0100001000",  -- INDEX 264
	B"10110011" when B"0100001001",  -- INDEX 265
	B"11011111" when B"0100001010",  -- INDEX 266
	B"00010001" when B"0100001011",  -- INDEX 267
	B"00111111" when B"0100001100",  -- INDEX 268
	B"01100101" when B"0100001101",  -- INDEX 269
	B"01111011" when B"0100001110",  -- INDEX 270
	B"01111111" when B"0100001111",  -- INDEX 271
	B"01110000" when B"0100010000",  -- INDEX 272
	B"01010000" when B"0100010001",  -- INDEX 273
	B"00100101" when B"0100010010",  -- INDEX 274
	B"11110011" when B"0100010011",  -- INDEX 275
	B"11000100" when B"0100010100",  -- INDEX 276
	B"10011110" when B"0100010101",  -- INDEX 277
	B"10000110" when B"0100010110",  -- INDEX 278
	B"10000000" when B"0100010111",  -- INDEX 279
	B"10001110" when B"0100011000",  -- INDEX 280
	B"10101100" when B"0100011001",  -- INDEX 281
	B"11010111" when B"0100011010",  -- INDEX 282
	B"00001001" when B"0100011011",  -- INDEX 283
	B"00111000" when B"0100011100",  -- INDEX 284
	B"01100000" when B"0100011101",  -- INDEX 285
	B"01111001" when B"0100011110",  -- INDEX 286
	B"01111111" when B"0100011111",  -- INDEX 287
	B"01110100" when B"0100100000",  -- INDEX 288
	B"01010111" when B"0100100001",  -- INDEX 289
	B"00101100" when B"0100100010",  -- INDEX 290
	B"11111011" when B"0100100011",  -- INDEX 291
	B"11001011" when B"0100100100",  -- INDEX 292
	B"10100011" when B"0100100101",  -- INDEX 293
	B"10001001" when B"0100100110",  -- INDEX 294
	B"10000000" when B"0100100111",  -- INDEX 295
	B"10001011" when B"0100101000",  -- INDEX 296
	B"10100111" when B"0100101001",  -- INDEX 297
	B"11010000" when B"0100101010",  -- INDEX 298
	B"00000001" when B"0100101011",  -- INDEX 299
	B"00110001" when B"0100101100",  -- INDEX 300
	B"01011010" when B"0100101101",  -- INDEX 301
	B"01110110" when B"0100101110",  -- INDEX 302
	B"01111111" when B"0100101111",  -- INDEX 303
	B"01110111" when B"0100110000",  -- INDEX 304
	B"01011100" when B"0100110001",  -- INDEX 305
	B"00110100" when B"0100110010",  -- INDEX 306
	B"00000100" when B"0100110011",  -- INDEX 307
	B"11010011" when B"0100110100",  -- INDEX 308
	B"10101001" when B"0100110101",  -- INDEX 309
	B"10001100" when B"0100110110",  -- INDEX 310
	B"10000000" when B"0100110111",  -- INDEX 311
	B"10001000" when B"0100111000",  -- INDEX 312
	B"10100001" when B"0100111001",  -- INDEX 313
	B"11001001" when B"0100111010",  -- INDEX 314
	B"11111000" when B"0100111011",  -- INDEX 315
	B"00101001" when B"0100111100",  -- INDEX 316
	B"01010100" when B"0100111101",  -- INDEX 317
	B"01110011" when B"0100111110",  -- INDEX 318
	B"01111111" when B"0100111111",  -- INDEX 319
	B"01111010" when B"0101000000",  -- INDEX 320
	B"01100010" when B"0101000001",  -- INDEX 321
	B"00111011" when B"0101000010",  -- INDEX 322
	B"00001100" when B"0101000011",  -- INDEX 323
	B"11011010" when B"0101000100",  -- INDEX 324
	B"10101111" when B"0101000101",  -- INDEX 325
	B"10001111" when B"0101000110",  -- INDEX 326
	B"10000001" when B"0101000111",  -- INDEX 327
	B"10000101" when B"0101001000",  -- INDEX 328
	B"10011100" when B"0101001001",  -- INDEX 329
	B"11000001" when B"0101001010",  -- INDEX 330
	B"11110000" when B"0101001011",  -- INDEX 331
	B"00100010" when B"0101001100",  -- INDEX 332
	B"01001110" when B"0101001101",  -- INDEX 333
	B"01101111" when B"0101001110",  -- INDEX 334
	B"01111111" when B"0101001111",  -- INDEX 335
	B"01111100" when B"0101010000",  -- INDEX 336
	B"01100111" when B"0101010001",  -- INDEX 337
	B"01000010" when B"0101010010",  -- INDEX 338
	B"00010100" when B"0101010011",  -- INDEX 339
	B"11100010" when B"0101010100",  -- INDEX 340
	B"10110101" when B"0101010101",  -- INDEX 341
	B"10010011" when B"0101010110",  -- INDEX 342
	B"10000010" when B"0101010111",  -- INDEX 343
	B"10000011" when B"0101011000",  -- INDEX 344
	B"10010111" when B"0101011001",  -- INDEX 345
	B"10111011" when B"0101011010",  -- INDEX 346
	B"11101001" when B"0101011011",  -- INDEX 347
	B"00011010" when B"0101011100",  -- INDEX 348
	B"01001000" when B"0101011101",  -- INDEX 349
	B"01101010" when B"0101011110",  -- INDEX 350
	B"01111101" when B"0101011111",  -- INDEX 351
	B"01111110" when B"0101100000",  -- INDEX 352
	B"01101011" when B"0101100001",  -- INDEX 353
	B"01001001" when B"0101100010",  -- INDEX 354
	B"00011011" when B"0101100011",  -- INDEX 355
	B"11101010" when B"0101100100",  -- INDEX 356
	B"10111100" when B"0101100101",  -- INDEX 357
	B"10011000" when B"0101100110",  -- INDEX 358
	B"10000011" when B"0101100111",  -- INDEX 359
	B"10000010" when B"0101101000",  -- INDEX 360
	B"10010011" when B"0101101001",  -- INDEX 361
	B"10110100" when B"0101101010",  -- INDEX 362
	B"11100001" when B"0101101011",  -- INDEX 363
	B"00010010" when B"0101101100",  -- INDEX 364
	B"01000001" when B"0101101101",  -- INDEX 365
	B"01100110" when B"0101101110",  -- INDEX 366
	B"01111100" when B"0101101111",  -- INDEX 367
	B"01111111" when B"0101110000",  -- INDEX 368
	B"01101111" when B"0101110001",  -- INDEX 369
	B"01001111" when B"0101110010",  -- INDEX 370
	B"00100011" when B"0101110011",  -- INDEX 371
	B"11110010" when B"0101110100",  -- INDEX 372
	B"11000011" when B"0101110101",  -- INDEX 373
	B"10011101" when B"0101110110",  -- INDEX 374
	B"10000110" when B"0101110111",  -- INDEX 375
	B"10000001" when B"0101111000",  -- INDEX 376
	B"10001111" when B"0101111001",  -- INDEX 377
	B"10101110" when B"0101111010",  -- INDEX 378
	B"11011001" when B"0101111011",  -- INDEX 379
	B"00001010" when B"0101111100",  -- INDEX 380
	B"00111010" when B"0101111101",  -- INDEX 381
	B"01100001" when B"0101111110",  -- INDEX 382
	B"01111001" when B"0101111111",  -- INDEX 383
	B"01111111" when B"0110000000",  -- INDEX 384
	B"01110011" when B"0110000001",  -- INDEX 385
	B"01010101" when B"0110000010",  -- INDEX 386
	B"00101011" when B"0110000011",  -- INDEX 387
	B"11111010" when B"0110000100",  -- INDEX 388
	B"11001010" when B"0110000101",  -- INDEX 389
	B"10100010" when B"0110000110",  -- INDEX 390
	B"10001000" when B"0110000111",  -- INDEX 391
	B"10000000" when B"0110001000",  -- INDEX 392
	B"10001011" when B"0110001001",  -- INDEX 393
	B"10101000" when B"0110001010",  -- INDEX 394
	B"11010001" when B"0110001011",  -- INDEX 395
	B"00000010" when B"0110001100",  -- INDEX 396
	B"00110010" when B"0110001101",  -- INDEX 397
	B"01011011" when B"0110001110",  -- INDEX 398
	B"01110110" when B"0110001111",  -- INDEX 399
	B"01111111" when B"0110010000",  -- INDEX 400
	B"01110110" when B"0110010001",  -- INDEX 401
	B"01011010" when B"0110010010",  -- INDEX 402
	B"00110000" when B"0110010011",  -- INDEX 403
	B"11111110" when B"0110010100",  -- INDEX 404
	B"11001101" when B"0110010101",  -- INDEX 405
	B"10100011" when B"0110010110",  -- INDEX 406
	B"10001000" when B"0110010111",  -- INDEX 407
	B"10000000" when B"0110011000",  -- INDEX 408
	B"10001100" when B"0110011001",  -- INDEX 409
	B"10101001" when B"0110011010",  -- INDEX 410
	B"11010100" when B"0110011011",  -- INDEX 411
	B"00000110" when B"0110011100",  -- INDEX 412
	B"00110111" when B"0110011101",  -- INDEX 413
	B"01011111" when B"0110011110",  -- INDEX 414
	B"01111001" when B"0110011111",  -- INDEX 415
	B"01111111" when B"0110100000",  -- INDEX 416
	B"01110011" when B"0110100001",  -- INDEX 417
	B"01010100" when B"0110100010",  -- INDEX 418
	B"00101000" when B"0110100011",  -- INDEX 419
	B"11110110" when B"0110100100",  -- INDEX 420
	B"11000101" when B"0110100101",  -- INDEX 421
	B"10011110" when B"0110100110",  -- INDEX 422
	B"10000110" when B"0110100111",  -- INDEX 423
	B"10000001" when B"0110101000",  -- INDEX 424
	B"10001111" when B"0110101001",  -- INDEX 425
	B"10101111" when B"0110101010",  -- INDEX 426
	B"11011100" when B"0110101011",  -- INDEX 427
	B"00001110" when B"0110101100",  -- INDEX 428
	B"00111110" when B"0110101101",  -- INDEX 429
	B"01100101" when B"0110101110",  -- INDEX 430
	B"01111011" when B"0110101111",  -- INDEX 431
	B"01111111" when B"0110110000",  -- INDEX 432
	B"01101111" when B"0110110001",  -- INDEX 433
	B"01001110" when B"0110110010",  -- INDEX 434
	B"00100000" when B"0110110011",  -- INDEX 435
	B"11101110" when B"0110110100",  -- INDEX 436
	B"10111110" when B"0110110101",  -- INDEX 437
	B"10011001" when B"0110110110",  -- INDEX 438
	B"10000100" when B"0110110111",  -- INDEX 439
	B"10000010" when B"0110111000",  -- INDEX 440
	B"10010011" when B"0110111001",  -- INDEX 441
	B"10110110" when B"0110111010",  -- INDEX 442
	B"11100100" when B"0110111011",  -- INDEX 443
	B"00010110" when B"0110111100",  -- INDEX 444
	B"01000101" when B"0110111101",  -- INDEX 445
	B"01101001" when B"0110111110",  -- INDEX 446
	B"01111101" when B"0110111111",  -- INDEX 447
	B"01111110" when B"0111000000",  -- INDEX 448
	B"01101011" when B"0111000001",  -- INDEX 449
	B"01000111" when B"0111000010",  -- INDEX 450
	B"00011000" when B"0111000011",  -- INDEX 451
	B"11100110" when B"0111000100",  -- INDEX 452
	B"10111000" when B"0111000101",  -- INDEX 453
	B"10010100" when B"0111000110",  -- INDEX 454
	B"10000010" when B"0111000111",  -- INDEX 455
	B"10000011" when B"0111001000",  -- INDEX 456
	B"10011000" when B"0111001001",  -- INDEX 457
	B"10111100" when B"0111001010",  -- INDEX 458
	B"11101011" when B"0111001011",  -- INDEX 459
	B"00011110" when B"0111001100",  -- INDEX 460
	B"01001100" when B"0111001101",  -- INDEX 461
	B"01101110" when B"0111001110",  -- INDEX 462
	B"01111111" when B"0111001111",  -- INDEX 463
	B"01111100" when B"0111010000",  -- INDEX 464
	B"01100110" when B"0111010001",  -- INDEX 465
	B"01000000" when B"0111010010",  -- INDEX 466
	B"00010001" when B"0111010011",  -- INDEX 467
	B"11011110" when B"0111010100",  -- INDEX 468
	B"10110001" when B"0111010101",  -- INDEX 469
	B"10010000" when B"0111010110",  -- INDEX 470
	B"10000001" when B"0111010111",  -- INDEX 471
	B"10000101" when B"0111011000",  -- INDEX 472
	B"10011100" when B"0111011001",  -- INDEX 473
	B"11000011" when B"0111011010",  -- INDEX 474
	B"11110011" when B"0111011011",  -- INDEX 475
	B"00100110" when B"0111011100",  -- INDEX 476
	B"01010010" when B"0111011101",  -- INDEX 477
	B"01110010" when B"0111011110",  -- INDEX 478
	B"01111111" when B"0111011111",  -- INDEX 479
	B"01111010" when B"0111100000",  -- INDEX 480
	B"01100001" when B"0111100001",  -- INDEX 481
	B"00111001" when B"0111100010",  -- INDEX 482
	B"00001001" when B"0111100011",  -- INDEX 483
	B"11010111" when B"0111100100",  -- INDEX 484
	B"10101011" when B"0111100101",  -- INDEX 485
	B"10001101" when B"0111100110",  -- INDEX 486
	B"10000000" when B"0111100111",  -- INDEX 487
	B"10001000" when B"0111101000",  -- INDEX 488
	B"10100010" when B"0111101001",  -- INDEX 489
	B"11001010" when B"0111101010",  -- INDEX 490
	B"11111011" when B"0111101011",  -- INDEX 491
	B"00101101" when B"0111101100",  -- INDEX 492
	B"01011000" when B"0111101101",  -- INDEX 493
	B"01110101" when B"0111101110",  -- INDEX 494
	B"01111111" when B"0111101111",  -- INDEX 495
	B"01110111" when B"0111110000",  -- INDEX 496
	B"01011100" when B"0111110001",  -- INDEX 497
	B"00110010" when B"0111110010",  -- INDEX 498
	B"00000001" when B"0111110011",  -- INDEX 499
	B"11001111" when B"0111110100",  -- INDEX 500
	B"10100101" when B"0111110101",  -- INDEX 501
	B"10001001" when B"0111110110",  -- INDEX 502
	B"10000000" when B"0111110111",  -- INDEX 503
	B"10001011" when B"0111111000",  -- INDEX 504
	B"10100111" when B"0111111001",  -- INDEX 505
	B"11010010" when B"0111111010",  -- INDEX 506
	B"00000100" when B"0111111011",  -- INDEX 507
	B"00110101" when B"0111111100",  -- INDEX 508
	B"01011110" when B"0111111101",  -- INDEX 509
	B"01111000" when B"0111111110",  -- INDEX 510
	B"01111111" when B"0111111111",  -- INDEX 511
	B"01110100" when B"1000000000",  -- INDEX 512
	B"01010110" when B"1000000001",  -- INDEX 513
	B"00101010" when B"1000000010",  -- INDEX 514
	B"11111000" when B"1000000011",  -- INDEX 515
	B"11001000" when B"1000000100",  -- INDEX 516
	B"10100000" when B"1000000101",  -- INDEX 517
	B"10000111" when B"1000000110",  -- INDEX 518
	B"10000000" when B"1000000111",  -- INDEX 519
	B"10001110" when B"1000001000",  -- INDEX 520
	B"10101101" when B"1000001001",  -- INDEX 521
	B"11011001" when B"1000001010",  -- INDEX 522
	B"00001100" when B"1000001011",  -- INDEX 523
	B"00111100" when B"1000001100",  -- INDEX 524
	B"01100011" when B"1000001101",  -- INDEX 525
	B"01111011" when B"1000001110",  -- INDEX 526
	B"01111111" when B"1000001111",  -- INDEX 527
	B"01110000" when B"1000010000",  -- INDEX 528
	B"01010000" when B"1000010001",  -- INDEX 529
	B"00100011" when B"1000010010",  -- INDEX 530
	B"11110000" when B"1000010011",  -- INDEX 531
	B"11000001" when B"1000010100",  -- INDEX 532
	B"10011011" when B"1000010101",  -- INDEX 533
	B"10000100" when B"1000010110",  -- INDEX 534
	B"10000001" when B"1000010111",  -- INDEX 535
	B"10010010" when B"1000011000",  -- INDEX 536
	B"10110100" when B"1000011001",  -- INDEX 537
	B"11100001" when B"1000011010",  -- INDEX 538
	B"00010100" when B"1000011011",  -- INDEX 539
	B"01000011" when B"1000011100",  -- INDEX 540
	B"01101000" when B"1000011101",  -- INDEX 541
	B"01111101" when B"1000011110",  -- INDEX 542
	B"01111110" when B"1000011111",  -- INDEX 543
	B"01101100" when B"1000100000",  -- INDEX 544
	B"01001001" when B"1000100001",  -- INDEX 545
	B"00011011" when B"1000100010",  -- INDEX 546
	B"11101001" when B"1000100011",  -- INDEX 547
	B"10111010" when B"1000100100",  -- INDEX 548
	B"10010110" when B"1000100101",  -- INDEX 549
	B"10000010" when B"1000100110",  -- INDEX 550
	B"10000011" when B"1000100111",  -- INDEX 551
	B"10010110" when B"1000101000",  -- INDEX 552
	B"10111010" when B"1000101001",  -- INDEX 553
	B"11101001" when B"1000101010",  -- INDEX 554
	B"00011011" when B"1000101011",  -- INDEX 555
	B"01001010" when B"1000101100",  -- INDEX 556
	B"01101100" when B"1000101101",  -- INDEX 557
	B"01111110" when B"1000101110",  -- INDEX 558
	B"01111101" when B"1000101111",  -- INDEX 559
	B"01101000" when B"1000110000",  -- INDEX 560
	B"01000010" when B"1000110001",  -- INDEX 561
	B"00010011" when B"1000110010",  -- INDEX 562
	B"11100001" when B"1000110011",  -- INDEX 563
	B"10110011" when B"1000110100",  -- INDEX 564
	B"10010010" when B"1000110101",  -- INDEX 565
	B"10000001" when B"1000110110",  -- INDEX 566
	B"10000100" when B"1000110111",  -- INDEX 567
	B"10011011" when B"1000111000",  -- INDEX 568
	B"11000001" when B"1000111001",  -- INDEX 569
	B"11110001" when B"1000111010",  -- INDEX 570
	B"00100011" when B"1000111011",  -- INDEX 571
	B"01010000" when B"1000111100",  -- INDEX 572
	B"01110000" when B"1000111101",  -- INDEX 573
	B"01111111" when B"1000111110",  -- INDEX 574
	B"01111010" when B"1000111111",  -- INDEX 575
	B"01100011" when B"1001000000",  -- INDEX 576
	B"00111011" when B"1001000001",  -- INDEX 577
	B"00001011" when B"1001000010",  -- INDEX 578
	B"11011001" when B"1001000011",  -- INDEX 579
	B"10101101" when B"1001000100",  -- INDEX 580
	B"10001110" when B"1001000101",  -- INDEX 581
	B"10000000" when B"1001000110",  -- INDEX 582
	B"10000111" when B"1001000111",  -- INDEX 583
	B"10100000" when B"1001001000",  -- INDEX 584
	B"11001000" when B"1001001001",  -- INDEX 585
	B"11111001" when B"1001001010",  -- INDEX 586
	B"00101011" when B"1001001011",  -- INDEX 587
	B"01010110" when B"1001001100",  -- INDEX 588
	B"01110100" when B"1001001101",  -- INDEX 589
	B"01111111" when B"1001001110",  -- INDEX 590
	B"01111000" when B"1001001111",  -- INDEX 591
	B"01011101" when B"1001010000",  -- INDEX 592
	B"00110100" when B"1001010001",  -- INDEX 593
	B"00000011" when B"1001010010",  -- INDEX 594
	B"11010001" when B"1001010011",  -- INDEX 595
	B"10100111" when B"1001010100",  -- INDEX 596
	B"10001010" when B"1001010101",  -- INDEX 597
	B"10000000" when B"1001010110",  -- INDEX 598
	B"10001010" when B"1001010111",  -- INDEX 599
	B"10100101" when B"1001011000",  -- INDEX 600
	B"11001111" when B"1001011001",  -- INDEX 601
	B"11111111" when B"1001011010",  -- INDEX 602
	B"00110000" when B"1001011011",  -- INDEX 603
	B"01011001" when B"1001011100",  -- INDEX 604
	B"01110101" when B"1001011101",  -- INDEX 605
	B"01111111" when B"1001011110",  -- INDEX 606
	B"01111000" when B"1001011111",  -- INDEX 607
	B"01011101" when B"1001100000",  -- INDEX 608
	B"00110101" when B"1001100001",  -- INDEX 609
	B"00000101" when B"1001100010",  -- INDEX 610
	B"11010100" when B"1001100011",  -- INDEX 611
	B"10101010" when B"1001100100",  -- INDEX 612
	B"10001100" when B"1001100101",  -- INDEX 613
	B"10000000" when B"1001100110",  -- INDEX 614
	B"10000111" when B"1001100111",  -- INDEX 615
	B"10100000" when B"1001101000",  -- INDEX 616
	B"11000111" when B"1001101001",  -- INDEX 617
	B"11110111" when B"1001101010",  -- INDEX 618
	B"00101000" when B"1001101011",  -- INDEX 619
	B"01010011" when B"1001101100",  -- INDEX 620
	B"01110010" when B"1001101101",  -- INDEX 621
	B"01111111" when B"1001101110",  -- INDEX 622
	B"01111010" when B"1001101111",  -- INDEX 623
	B"01100011" when B"1001110000",  -- INDEX 624
	B"00111100" when B"1001110001",  -- INDEX 625
	B"00001101" when B"1001110010",  -- INDEX 626
	B"11011100" when B"1001110011",  -- INDEX 627
	B"10110000" when B"1001110100",  -- INDEX 628
	B"10010000" when B"1001110101",  -- INDEX 629
	B"10000001" when B"1001110110",  -- INDEX 630
	B"10000101" when B"1001110111",  -- INDEX 631
	B"10011011" when B"1001111000",  -- INDEX 632
	B"11000000" when B"1001111001",  -- INDEX 633
	B"11101111" when B"1001111010",  -- INDEX 634
	B"00100000" when B"1001111011",  -- INDEX 635
	B"01001101" when B"1001111100",  -- INDEX 636
	B"01101110" when B"1001111101",  -- INDEX 637
	B"01111111" when B"1001111110",  -- INDEX 638
	B"01111100" when B"1001111111",  -- INDEX 639
	B"01101000" when B"1010000000",  -- INDEX 640
	B"01000011" when B"1010000001",  -- INDEX 641
	B"00010101" when B"1010000010",  -- INDEX 642
	B"11100100" when B"1010000011",  -- INDEX 643
	B"10110110" when B"1010000100",  -- INDEX 644
	B"10010100" when B"1010000101",  -- INDEX 645
	B"10000010" when B"1010000110",  -- INDEX 646
	B"10000011" when B"1010000111",  -- INDEX 647
	B"10010110" when B"1010001000",  -- INDEX 648
	B"10111001" when B"1010001001",  -- INDEX 649
	B"11100111" when B"1010001010",  -- INDEX 650
	B"00011000" when B"1010001011",  -- INDEX 651
	B"01000110" when B"1010001100",  -- INDEX 652
	B"01101010" when B"1010001101",  -- INDEX 653
	B"01111101" when B"1010001110",  -- INDEX 654
	B"01111110" when B"1010001111",  -- INDEX 655
	B"01101100" when B"1010010000",  -- INDEX 656
	B"01001010" when B"1010010001",  -- INDEX 657
	B"00011101" when B"1010010010",  -- INDEX 658
	B"11101011" when B"1010010011",  -- INDEX 659
	B"10111101" when B"1010010100",  -- INDEX 660
	B"10011001" when B"1010010101",  -- INDEX 661
	B"10000100" when B"1010010110",  -- INDEX 662
	B"10000001" when B"1010010111",  -- INDEX 663
	B"10010010" when B"1010011000",  -- INDEX 664
	B"10110011" when B"1010011001",  -- INDEX 665
	B"11011111" when B"1010011010",  -- INDEX 666
	B"00010001" when B"1010011011",  -- INDEX 667
	B"00111111" when B"1010011100",  -- INDEX 668
	B"01100101" when B"1010011101",  -- INDEX 669
	B"01111011" when B"1010011110",  -- INDEX 670
	B"01111111" when B"1010011111",  -- INDEX 671
	B"01110000" when B"1010100000",  -- INDEX 672
	B"01010000" when B"1010100001",  -- INDEX 673
	B"00100101" when B"1010100010",  -- INDEX 674
	B"11110011" when B"1010100011",  -- INDEX 675
	B"11000100" when B"1010100100",  -- INDEX 676
	B"10011110" when B"1010100101",  -- INDEX 677
	B"10000110" when B"1010100110",  -- INDEX 678
	B"10000000" when B"1010100111",  -- INDEX 679
	B"10001110" when B"1010101000",  -- INDEX 680
	B"10101100" when B"1010101001",  -- INDEX 681
	B"11010111" when B"1010101010",  -- INDEX 682
	B"00001001" when B"1010101011",  -- INDEX 683
	B"00111000" when B"1010101100",  -- INDEX 684
	B"01100000" when B"1010101101",  -- INDEX 685
	B"01111001" when B"1010101110",  -- INDEX 686
	B"01111111" when B"1010101111",  -- INDEX 687
	B"01110100" when B"1010110000",  -- INDEX 688
	B"01010111" when B"1010110001",  -- INDEX 689
	B"00101100" when B"1010110010",  -- INDEX 690
	B"11111011" when B"1010110011",  -- INDEX 691
	B"11001011" when B"1010110100",  -- INDEX 692
	B"10100011" when B"1010110101",  -- INDEX 693
	B"10001001" when B"1010110110",  -- INDEX 694
	B"10000000" when B"1010110111",  -- INDEX 695
	B"10001011" when B"1010111000",  -- INDEX 696
	B"10100111" when B"1010111001",  -- INDEX 697
	B"11010000" when B"1010111010",  -- INDEX 698
	B"00000001" when B"1010111011",  -- INDEX 699
	B"00110001" when B"1010111100",  -- INDEX 700
	B"01011010" when B"1010111101",  -- INDEX 701
	B"01110110" when B"1010111110",  -- INDEX 702
	B"01111111" when B"1010111111",  -- INDEX 703
	B"01110111" when B"1011000000",  -- INDEX 704
	B"01011100" when B"1011000001",  -- INDEX 705
	B"00110100" when B"1011000010",  -- INDEX 706
	B"00000100" when B"1011000011",  -- INDEX 707
	B"11010011" when B"1011000100",  -- INDEX 708
	B"10101001" when B"1011000101",  -- INDEX 709
	B"10001100" when B"1011000110",  -- INDEX 710
	B"10000000" when B"1011000111",  -- INDEX 711
	B"10001000" when B"1011001000",  -- INDEX 712
	B"10100001" when B"1011001001",  -- INDEX 713
	B"11001001" when B"1011001010",  -- INDEX 714
	B"11111000" when B"1011001011",  -- INDEX 715
	B"00101001" when B"1011001100",  -- INDEX 716
	B"01010100" when B"1011001101",  -- INDEX 717
	B"01110011" when B"1011001110",  -- INDEX 718
	B"01111111" when B"1011001111",  -- INDEX 719
	B"01111010" when B"1011010000",  -- INDEX 720
	B"01100010" when B"1011010001",  -- INDEX 721
	B"00111011" when B"1011010010",  -- INDEX 722
	B"00001100" when B"1011010011",  -- INDEX 723
	B"11011010" when B"1011010100",  -- INDEX 724
	B"10101111" when B"1011010101",  -- INDEX 725
	B"10001111" when B"1011010110",  -- INDEX 726
	B"10000001" when B"1011010111",  -- INDEX 727
	B"10000101" when B"1011011000",  -- INDEX 728
	B"10011100" when B"1011011001",  -- INDEX 729
	B"11000001" when B"1011011010",  -- INDEX 730
	B"11110000" when B"1011011011",  -- INDEX 731
	B"00100010" when B"1011011100",  -- INDEX 732
	B"01001110" when B"1011011101",  -- INDEX 733
	B"01101111" when B"1011011110",  -- INDEX 734
	B"01111111" when B"1011011111",  -- INDEX 735
	B"01111100" when B"1011100000",  -- INDEX 736
	B"01100111" when B"1011100001",  -- INDEX 737
	B"01000010" when B"1011100010",  -- INDEX 738
	B"00010100" when B"1011100011",  -- INDEX 739
	B"11100010" when B"1011100100",  -- INDEX 740
	B"10110101" when B"1011100101",  -- INDEX 741
	B"10010011" when B"1011100110",  -- INDEX 742
	B"10000010" when B"1011100111",  -- INDEX 743
	B"10000011" when B"1011101000",  -- INDEX 744
	B"10010111" when B"1011101001",  -- INDEX 745
	B"10111011" when B"1011101010",  -- INDEX 746
	B"11101001" when B"1011101011",  -- INDEX 747
	B"00011010" when B"1011101100",  -- INDEX 748
	B"01001000" when B"1011101101",  -- INDEX 749
	B"01101010" when B"1011101110",  -- INDEX 750
	B"01111101" when B"1011101111",  -- INDEX 751
	B"01111110" when B"1011110000",  -- INDEX 752
	B"01101011" when B"1011110001",  -- INDEX 753
	B"01001001" when B"1011110010",  -- INDEX 754
	B"00011011" when B"1011110011",  -- INDEX 755
	B"11101010" when B"1011110100",  -- INDEX 756
	B"10111100" when B"1011110101",  -- INDEX 757
	B"10011000" when B"1011110110",  -- INDEX 758
	B"10000011" when B"1011110111",  -- INDEX 759
	B"10000010" when B"1011111000",  -- INDEX 760
	B"10010011" when B"1011111001",  -- INDEX 761
	B"10110100" when B"1011111010",  -- INDEX 762
	B"11100001" when B"1011111011",  -- INDEX 763
	B"00010010" when B"1011111100",  -- INDEX 764
	B"01000001" when B"1011111101",  -- INDEX 765
	B"01100110" when B"1011111110",  -- INDEX 766
	B"01111100" when B"1011111111",  -- INDEX 767
	B"01111111" when B"1100000000",  -- INDEX 768
	B"01101111" when B"1100000001",  -- INDEX 769
	B"01001111" when B"1100000010",  -- INDEX 770
	B"00100011" when B"1100000011",  -- INDEX 771
	B"11110010" when B"1100000100",  -- INDEX 772
	B"11000011" when B"1100000101",  -- INDEX 773
	B"10011101" when B"1100000110",  -- INDEX 774
	B"10000110" when B"1100000111",  -- INDEX 775
	B"10000001" when B"1100001000",  -- INDEX 776
	B"10001111" when B"1100001001",  -- INDEX 777
	B"10101110" when B"1100001010",  -- INDEX 778
	B"11011001" when B"1100001011",  -- INDEX 779
	B"00001010" when B"1100001100",  -- INDEX 780
	B"00111010" when B"1100001101",  -- INDEX 781
	B"01100001" when B"1100001110",  -- INDEX 782
	B"01111001" when B"1100001111",  -- INDEX 783
	B"01111111" when B"1100010000",  -- INDEX 784
	B"01110011" when B"1100010001",  -- INDEX 785
	B"01010101" when B"1100010010",  -- INDEX 786
	B"00101011" when B"1100010011",  -- INDEX 787
	B"11111010" when B"1100010100",  -- INDEX 788
	B"11001010" when B"1100010101",  -- INDEX 789
	B"10100010" when B"1100010110",  -- INDEX 790
	B"10001000" when B"1100010111",  -- INDEX 791
	B"10000000" when B"1100011000",  -- INDEX 792
	B"10001011" when B"1100011001",  -- INDEX 793
	B"10101000" when B"1100011010",  -- INDEX 794
	B"11010001" when B"1100011011",  -- INDEX 795
	B"00000010" when B"1100011100",  -- INDEX 796
	B"00110010" when B"1100011101",  -- INDEX 797
	B"01011011" when B"1100011110",  -- INDEX 798
	B"01110110" when B"1100011111",  -- INDEX 799
	B"01111111" when B"1100100000",  -- INDEX 800
	B"01110110" when B"1100100001",  -- INDEX 801
	B"01011010" when B"1100100010",  -- INDEX 802
	B"00110000" when B"1100100011",  -- INDEX 803
	B"11111110" when B"1100100100",  -- INDEX 804
	B"11001101" when B"1100100101",  -- INDEX 805
	B"10100011" when B"1100100110",  -- INDEX 806
	B"10001000" when B"1100100111",  -- INDEX 807
	B"10000000" when B"1100101000",  -- INDEX 808
	B"10001100" when B"1100101001",  -- INDEX 809
	B"10101001" when B"1100101010",  -- INDEX 810
	B"11010100" when B"1100101011",  -- INDEX 811
	B"00000110" when B"1100101100",  -- INDEX 812
	B"00110111" when B"1100101101",  -- INDEX 813
	B"01011111" when B"1100101110",  -- INDEX 814
	B"01111001" when B"1100101111",  -- INDEX 815
	B"01111111" when B"1100110000",  -- INDEX 816
	B"01110011" when B"1100110001",  -- INDEX 817
	B"01010100" when B"1100110010",  -- INDEX 818
	B"00101000" when B"1100110011",  -- INDEX 819
	B"11110110" when B"1100110100",  -- INDEX 820
	B"11000101" when B"1100110101",  -- INDEX 821
	B"10011110" when B"1100110110",  -- INDEX 822
	B"10000110" when B"1100110111",  -- INDEX 823
	B"10000001" when B"1100111000",  -- INDEX 824
	B"10001111" when B"1100111001",  -- INDEX 825
	B"10101111" when B"1100111010",  -- INDEX 826
	B"11011100" when B"1100111011",  -- INDEX 827
	B"00001110" when B"1100111100",  -- INDEX 828
	B"00111110" when B"1100111101",  -- INDEX 829
	B"01100101" when B"1100111110",  -- INDEX 830
	B"01111011" when B"1100111111",  -- INDEX 831
	B"01111111" when B"1101000000",  -- INDEX 832
	B"01101111" when B"1101000001",  -- INDEX 833
	B"01001110" when B"1101000010",  -- INDEX 834
	B"00100000" when B"1101000011",  -- INDEX 835
	B"11101110" when B"1101000100",  -- INDEX 836
	B"10111110" when B"1101000101",  -- INDEX 837
	B"10011001" when B"1101000110",  -- INDEX 838
	B"10000100" when B"1101000111",  -- INDEX 839
	B"10000010" when B"1101001000",  -- INDEX 840
	B"10010011" when B"1101001001",  -- INDEX 841
	B"10110110" when B"1101001010",  -- INDEX 842
	B"11100100" when B"1101001011",  -- INDEX 843
	B"00010110" when B"1101001100",  -- INDEX 844
	B"01000101" when B"1101001101",  -- INDEX 845
	B"01101001" when B"1101001110",  -- INDEX 846
	B"01111101" when B"1101001111",  -- INDEX 847
	B"01111110" when B"1101010000",  -- INDEX 848
	B"01101011" when B"1101010001",  -- INDEX 849
	B"01000111" when B"1101010010",  -- INDEX 850
	B"00011000" when B"1101010011",  -- INDEX 851
	B"11100110" when B"1101010100",  -- INDEX 852
	B"10111000" when B"1101010101",  -- INDEX 853
	B"10010100" when B"1101010110",  -- INDEX 854
	B"10000010" when B"1101010111",  -- INDEX 855
	B"10000011" when B"1101011000",  -- INDEX 856
	B"10011000" when B"1101011001",  -- INDEX 857
	B"10111100" when B"1101011010",  -- INDEX 858
	B"11101011" when B"1101011011",  -- INDEX 859
	B"00011110" when B"1101011100",  -- INDEX 860
	B"01001100" when B"1101011101",  -- INDEX 861
	B"01101110" when B"1101011110",  -- INDEX 862
	B"01111111" when B"1101011111",  -- INDEX 863
	B"01111100" when B"1101100000",  -- INDEX 864
	B"01100110" when B"1101100001",  -- INDEX 865
	B"01000000" when B"1101100010",  -- INDEX 866
	B"00010001" when B"1101100011",  -- INDEX 867
	B"11011110" when B"1101100100",  -- INDEX 868
	B"10110001" when B"1101100101",  -- INDEX 869
	B"10010000" when B"1101100110",  -- INDEX 870
	B"10000001" when B"1101100111",  -- INDEX 871
	B"10000101" when B"1101101000",  -- INDEX 872
	B"10011100" when B"1101101001",  -- INDEX 873
	B"11000011" when B"1101101010",  -- INDEX 874
	B"11110011" when B"1101101011",  -- INDEX 875
	B"00100110" when B"1101101100",  -- INDEX 876
	B"01010010" when B"1101101101",  -- INDEX 877
	B"01110010" when B"1101101110",  -- INDEX 878
	B"01111111" when B"1101101111",  -- INDEX 879
	B"01111010" when B"1101110000",  -- INDEX 880
	B"01100001" when B"1101110001",  -- INDEX 881
	B"00111001" when B"1101110010",  -- INDEX 882
	B"00001001" when B"1101110011",  -- INDEX 883
	B"11010111" when B"1101110100",  -- INDEX 884
	B"10101011" when B"1101110101",  -- INDEX 885
	B"10001101" when B"1101110110",  -- INDEX 886
	B"10000000" when B"1101110111",  -- INDEX 887
	B"10001000" when B"1101111000",  -- INDEX 888
	B"10100010" when B"1101111001",  -- INDEX 889
	B"11001010" when B"1101111010",  -- INDEX 890
	B"11111011" when B"1101111011",  -- INDEX 891
	B"00101101" when B"1101111100",  -- INDEX 892
	B"01011000" when B"1101111101",  -- INDEX 893
	B"01110101" when B"1101111110",  -- INDEX 894
	B"01111111" when B"1101111111",  -- INDEX 895
	B"01110111" when B"1110000000",  -- INDEX 896
	B"01011100" when B"1110000001",  -- INDEX 897
	B"00110010" when B"1110000010",  -- INDEX 898
	B"00000001" when B"1110000011",  -- INDEX 899
	B"11001111" when B"1110000100",  -- INDEX 900
	B"10100101" when B"1110000101",  -- INDEX 901
	B"10001001" when B"1110000110",  -- INDEX 902
	B"10000000" when B"1110000111",  -- INDEX 903
	B"10001011" when B"1110001000",  -- INDEX 904
	B"10100111" when B"1110001001",  -- INDEX 905
	B"11010010" when B"1110001010",  -- INDEX 906
	B"00000100" when B"1110001011",  -- INDEX 907
	B"00110101" when B"1110001100",  -- INDEX 908
	B"01011110" when B"1110001101",  -- INDEX 909
	B"01111000" when B"1110001110",  -- INDEX 910
	B"01111111" when B"1110001111",  -- INDEX 911
	B"01110100" when B"1110010000",  -- INDEX 912
	B"01010110" when B"1110010001",  -- INDEX 913
	B"00101010" when B"1110010010",  -- INDEX 914
	B"11111000" when B"1110010011",  -- INDEX 915
	B"11001000" when B"1110010100",  -- INDEX 916
	B"10100000" when B"1110010101",  -- INDEX 917
	B"10000111" when B"1110010110",  -- INDEX 918
	B"10000000" when B"1110010111",  -- INDEX 919
	B"10001110" when B"1110011000",  -- INDEX 920
	B"10101101" when B"1110011001",  -- INDEX 921
	B"11011001" when B"1110011010",  -- INDEX 922
	B"00001100" when B"1110011011",  -- INDEX 923
	B"00111100" when B"1110011100",  -- INDEX 924
	B"01100011" when B"1110011101",  -- INDEX 925
	B"01111011" when B"1110011110",  -- INDEX 926
	B"01111111" when B"1110011111",  -- INDEX 927
	B"01110000" when B"1110100000",  -- INDEX 928
	B"01010000" when B"1110100001",  -- INDEX 929
	B"00100011" when B"1110100010",  -- INDEX 930
	B"11110000" when B"1110100011",  -- INDEX 931
	B"11000001" when B"1110100100",  -- INDEX 932
	B"10011011" when B"1110100101",  -- INDEX 933
	B"10000100" when B"1110100110",  -- INDEX 934
	B"10000001" when B"1110100111",  -- INDEX 935
	B"10010010" when B"1110101000",  -- INDEX 936
	B"10110100" when B"1110101001",  -- INDEX 937
	B"11100001" when B"1110101010",  -- INDEX 938
	B"00010100" when B"1110101011",  -- INDEX 939
	B"01000011" when B"1110101100",  -- INDEX 940
	B"01101000" when B"1110101101",  -- INDEX 941
	B"01111101" when B"1110101110",  -- INDEX 942
	B"01111110" when B"1110101111",  -- INDEX 943
	B"01101100" when B"1110110000",  -- INDEX 944
	B"01001001" when B"1110110001",  -- INDEX 945
	B"00011011" when B"1110110010",  -- INDEX 946
	B"11101001" when B"1110110011",  -- INDEX 947
	B"10111010" when B"1110110100",  -- INDEX 948
	B"10010110" when B"1110110101",  -- INDEX 949
	B"10000010" when B"1110110110",  -- INDEX 950
	B"10000011" when B"1110110111",  -- INDEX 951
	B"10010110" when B"1110111000",  -- INDEX 952
	B"10111010" when B"1110111001",  -- INDEX 953
	B"11101001" when B"1110111010",  -- INDEX 954
	B"00011011" when B"1110111011",  -- INDEX 955
	B"01001010" when B"1110111100",  -- INDEX 956
	B"01101100" when B"1110111101",  -- INDEX 957
	B"01111110" when B"1110111110",  -- INDEX 958
	B"01111101" when B"1110111111",  -- INDEX 959
	B"01101000" when B"1111000000",  -- INDEX 960
	B"01000010" when B"1111000001",  -- INDEX 961
	B"00010011" when B"1111000010",  -- INDEX 962
	B"11100001" when B"1111000011",  -- INDEX 963
	B"10110011" when B"1111000100",  -- INDEX 964
	B"10010010" when B"1111000101",  -- INDEX 965
	B"10000001" when B"1111000110",  -- INDEX 966
	B"10000100" when B"1111000111",  -- INDEX 967
	B"10011011" when B"1111001000",  -- INDEX 968
	B"11000001" when B"1111001001",  -- INDEX 969
	B"11110001" when B"1111001010",  -- INDEX 970
	B"00100011" when B"1111001011",  -- INDEX 971
	B"01010000" when B"1111001100",  -- INDEX 972
	B"01110000" when B"1111001101",  -- INDEX 973
	B"01111111" when B"1111001110",  -- INDEX 974
	B"01111010" when B"1111001111",  -- INDEX 975
	B"01100011" when B"1111010000",  -- INDEX 976
	B"00111011" when B"1111010001",  -- INDEX 977
	B"00001011" when B"1111010010",  -- INDEX 978
	B"11011001" when B"1111010011",  -- INDEX 979
	B"10101101" when B"1111010100",  -- INDEX 980
	B"10001110" when B"1111010101",  -- INDEX 981
	B"10000000" when B"1111010110",  -- INDEX 982
	B"10000111" when B"1111010111",  -- INDEX 983
	B"10100000" when B"1111011000",  -- INDEX 984
	B"11001000" when B"1111011001",  -- INDEX 985
	B"11111001" when B"1111011010",  -- INDEX 986
	B"00101011" when B"1111011011",  -- INDEX 987
	B"01010110" when B"1111011100",  -- INDEX 988
	B"01110100" when B"1111011101",  -- INDEX 989
	B"01111111" when B"1111011110",  -- INDEX 990
	B"01111000" when B"1111011111",  -- INDEX 991
	B"01011101" when B"1111100000",  -- INDEX 992
	B"00110100" when B"1111100001",  -- INDEX 993
	B"00000011" when B"1111100010",  -- INDEX 994
	B"11010001" when B"1111100011",  -- INDEX 995
	B"10100111" when B"1111100100",  -- INDEX 996
	B"10001010" when B"1111100101",  -- INDEX 997
	B"10000000" when B"1111100110",  -- INDEX 998
	B"10001010" when B"1111100111",  -- INDEX 999

-- END INPUT FM SIGNAL
	B"00000000" when others;
	
	with counter (09 downto 0) select
	test_signal_fmTri_int <=
-- START INPUT FM-TRI SIGNAL

	B"01111111" when B"0000000000",  -- INDEX 0
	B"01110110" when B"0000000001",  -- INDEX 1
	B"01011011" when B"0000000010",  -- INDEX 2
	B"00110010" when B"0000000011",  -- INDEX 3
	B"00000010" when B"0000000100",  -- INDEX 4
	B"11010001" when B"0000000101",  -- INDEX 5
	B"10101000" when B"0000000110",  -- INDEX 6
	B"10001011" when B"0000000111",  -- INDEX 7
	B"10000000" when B"0000001000",  -- INDEX 8
	B"10001000" when B"0000001001",  -- INDEX 9
	B"10100010" when B"0000001010",  -- INDEX 10
	B"11001010" when B"0000001011",  -- INDEX 11
	B"11111010" when B"0000001100",  -- INDEX 12
	B"00101011" when B"0000001101",  -- INDEX 13
	B"01010110" when B"0000001110",  -- INDEX 14
	B"01110011" when B"0000001111",  -- INDEX 15
	B"01111111" when B"0000010000",  -- INDEX 16
	B"01111001" when B"0000010001",  -- INDEX 17
	B"01100000" when B"0000010010",  -- INDEX 18
	B"00111001" when B"0000010011",  -- INDEX 19
	B"00001001" when B"0000010100",  -- INDEX 20
	B"11011000" when B"0000010101",  -- INDEX 21
	B"10101101" when B"0000010110",  -- INDEX 22
	B"10001110" when B"0000010111",  -- INDEX 23
	B"10000000" when B"0000011000",  -- INDEX 24
	B"10000110" when B"0000011001",  -- INDEX 25
	B"10011110" when B"0000011010",  -- INDEX 26
	B"11000100" when B"0000011011",  -- INDEX 27
	B"11110100" when B"0000011100",  -- INDEX 28
	B"00100101" when B"0000011101",  -- INDEX 29
	B"01010001" when B"0000011110",  -- INDEX 30
	B"01110001" when B"0000011111",  -- INDEX 31
	B"01111111" when B"0000100000",  -- INDEX 32
	B"01111011" when B"0000100001",  -- INDEX 33
	B"01100100" when B"0000100010",  -- INDEX 34
	B"00111110" when B"0000100011",  -- INDEX 35
	B"00001111" when B"0000100100",  -- INDEX 36
	B"11011101" when B"0000100101",  -- INDEX 37
	B"10110001" when B"0000100110",  -- INDEX 38
	B"10010001" when B"0000100111",  -- INDEX 39
	B"10000001" when B"0000101000",  -- INDEX 40
	B"10000100" when B"0000101001",  -- INDEX 41
	B"10011010" when B"0000101010",  -- INDEX 42
	B"11000000" when B"0000101011",  -- INDEX 43
	B"11101111" when B"0000101100",  -- INDEX 44
	B"00100000" when B"0000101101",  -- INDEX 45
	B"01001101" when B"0000101110",  -- INDEX 46
	B"01101110" when B"0000101111",  -- INDEX 47
	B"01111111" when B"0000110000",  -- INDEX 48
	B"01111100" when B"0000110001",  -- INDEX 49
	B"01100111" when B"0000110010",  -- INDEX 50
	B"01000010" when B"0000110011",  -- INDEX 51
	B"00010011" when B"0000110100",  -- INDEX 52
	B"11100010" when B"0000110101",  -- INDEX 53
	B"10110101" when B"0000110110",  -- INDEX 54
	B"10010011" when B"0000110111",  -- INDEX 55
	B"10000010" when B"0000111000",  -- INDEX 56
	B"10000011" when B"0000111001",  -- INDEX 57
	B"10011000" when B"0000111010",  -- INDEX 58
	B"10111100" when B"0000111011",  -- INDEX 59
	B"11101011" when B"0000111100",  -- INDEX 60
	B"00011101" when B"0000111101",  -- INDEX 61
	B"01001010" when B"0000111110",  -- INDEX 62
	B"01101100" when B"0000111111",  -- INDEX 63
	B"01111110" when B"0001000000",  -- INDEX 64
	B"01111101" when B"0001000001",  -- INDEX 65
	B"01101001" when B"0001000010",  -- INDEX 66
	B"01000101" when B"0001000011",  -- INDEX 67
	B"00010111" when B"0001000100",  -- INDEX 68
	B"11100101" when B"0001000101",  -- INDEX 69
	B"10110111" when B"0001000110",  -- INDEX 70
	B"10010101" when B"0001000111",  -- INDEX 71
	B"10000010" when B"0001001000",  -- INDEX 72
	B"10000011" when B"0001001001",  -- INDEX 73
	B"10010110" when B"0001001010",  -- INDEX 74
	B"10111010" when B"0001001011",  -- INDEX 75
	B"11101000" when B"0001001100",  -- INDEX 76
	B"00011010" when B"0001001101",  -- INDEX 77
	B"01001000" when B"0001001110",  -- INDEX 78
	B"01101011" when B"0001001111",  -- INDEX 79
	B"01111110" when B"0001010000",  -- INDEX 80
	B"01111101" when B"0001010001",  -- INDEX 81
	B"01101010" when B"0001010010",  -- INDEX 82
	B"01000111" when B"0001010011",  -- INDEX 83
	B"00011001" when B"0001010100",  -- INDEX 84
	B"11100111" when B"0001010101",  -- INDEX 85
	B"10111001" when B"0001010110",  -- INDEX 86
	B"10010101" when B"0001010111",  -- INDEX 87
	B"10000010" when B"0001011000",  -- INDEX 88
	B"10000010" when B"0001011001",  -- INDEX 89
	B"10010110" when B"0001011010",  -- INDEX 90
	B"10111001" when B"0001011011",  -- INDEX 91
	B"11100111" when B"0001011100",  -- INDEX 92
	B"00011001" when B"0001011101",  -- INDEX 93
	B"01000111" when B"0001011110",  -- INDEX 94
	B"01101010" when B"0001011111",  -- INDEX 95
	B"01111110" when B"0001100000",  -- INDEX 96
	B"01111110" when B"0001100001",  -- INDEX 97
	B"01101011" when B"0001100010",  -- INDEX 98
	B"01000111" when B"0001100011",  -- INDEX 99
	B"00011001" when B"0001100100",  -- INDEX 100
	B"11100111" when B"0001100101",  -- INDEX 101
	B"10111001" when B"0001100110",  -- INDEX 102
	B"10010110" when B"0001100111",  -- INDEX 103
	B"10000011" when B"0001101000",  -- INDEX 104
	B"10000010" when B"0001101001",  -- INDEX 105
	B"10010101" when B"0001101010",  -- INDEX 106
	B"10111001" when B"0001101011",  -- INDEX 107
	B"11100111" when B"0001101100",  -- INDEX 108
	B"00011001" when B"0001101101",  -- INDEX 109
	B"01000111" when B"0001101110",  -- INDEX 110
	B"01101010" when B"0001101111",  -- INDEX 111
	B"01111110" when B"0001110000",  -- INDEX 112
	B"01111110" when B"0001110001",  -- INDEX 113
	B"01101010" when B"0001110010",  -- INDEX 114
	B"01000111" when B"0001110011",  -- INDEX 115
	B"00011001" when B"0001110100",  -- INDEX 116
	B"11100111" when B"0001110101",  -- INDEX 117
	B"10111000" when B"0001110110",  -- INDEX 118
	B"10010101" when B"0001110111",  -- INDEX 119
	B"10000010" when B"0001111000",  -- INDEX 120
	B"10000011" when B"0001111001",  -- INDEX 121
	B"10010110" when B"0001111010",  -- INDEX 122
	B"10111010" when B"0001111011",  -- INDEX 123
	B"11101000" when B"0001111100",  -- INDEX 124
	B"00011010" when B"0001111101",  -- INDEX 125
	B"01001000" when B"0001111110",  -- INDEX 126
	B"01101011" when B"0001111111",  -- INDEX 127
	B"01111110" when B"0010000000",  -- INDEX 128
	B"01111101" when B"0010000001",  -- INDEX 129
	B"01101001" when B"0010000010",  -- INDEX 130
	B"01000101" when B"0010000011",  -- INDEX 131
	B"00010111" when B"0010000100",  -- INDEX 132
	B"11100101" when B"0010000101",  -- INDEX 133
	B"10110111" when B"0010000110",  -- INDEX 134
	B"10010100" when B"0010000111",  -- INDEX 135
	B"10000010" when B"0010001000",  -- INDEX 136
	B"10000011" when B"0010001001",  -- INDEX 137
	B"10010111" when B"0010001010",  -- INDEX 138
	B"10111100" when B"0010001011",  -- INDEX 139
	B"11101011" when B"0010001100",  -- INDEX 140
	B"00011101" when B"0010001101",  -- INDEX 141
	B"01001010" when B"0010001110",  -- INDEX 142
	B"01101101" when B"0010001111",  -- INDEX 143
	B"01111110" when B"0010010000",  -- INDEX 144
	B"01111101" when B"0010010001",  -- INDEX 145
	B"01101000" when B"0010010010",  -- INDEX 146
	B"01000011" when B"0010010011",  -- INDEX 147
	B"00010100" when B"0010010100",  -- INDEX 148
	B"11100010" when B"0010010101",  -- INDEX 149
	B"10110100" when B"0010010110",  -- INDEX 150
	B"10010010" when B"0010010111",  -- INDEX 151
	B"10000001" when B"0010011000",  -- INDEX 152
	B"10000100" when B"0010011001",  -- INDEX 153
	B"10011010" when B"0010011010",  -- INDEX 154
	B"10111111" when B"0010011011",  -- INDEX 155
	B"11101110" when B"0010011100",  -- INDEX 156
	B"00100001" when B"0010011101",  -- INDEX 157
	B"01001110" when B"0010011110",  -- INDEX 158
	B"01101111" when B"0010011111",  -- INDEX 159
	B"01111111" when B"0010100000",  -- INDEX 160
	B"01111011" when B"0010100001",  -- INDEX 161
	B"01100101" when B"0010100010",  -- INDEX 162
	B"00111111" when B"0010100011",  -- INDEX 163
	B"00001111" when B"0010100100",  -- INDEX 164
	B"11011101" when B"0010100101",  -- INDEX 165
	B"10110000" when B"0010100110",  -- INDEX 166
	B"10010000" when B"0010100111",  -- INDEX 167
	B"10000001" when B"0010101000",  -- INDEX 168
	B"10000101" when B"0010101001",  -- INDEX 169
	B"10011101" when B"0010101010",  -- INDEX 170
	B"11000011" when B"0010101011",  -- INDEX 171
	B"11110011" when B"0010101100",  -- INDEX 172
	B"00100110" when B"0010101101",  -- INDEX 173
	B"01010010" when B"0010101110",  -- INDEX 174
	B"01110001" when B"0010101111",  -- INDEX 175
	B"01111111" when B"0010110000",  -- INDEX 176
	B"01111010" when B"0010110001",  -- INDEX 177
	B"01100001" when B"0010110010",  -- INDEX 178
	B"00111010" when B"0010110011",  -- INDEX 179
	B"00001001" when B"0010110100",  -- INDEX 180
	B"11011000" when B"0010110101",  -- INDEX 181
	B"10101100" when B"0010110110",  -- INDEX 182
	B"10001101" when B"0010110111",  -- INDEX 183
	B"10000000" when B"0010111000",  -- INDEX 184
	B"10000111" when B"0010111001",  -- INDEX 185
	B"10100001" when B"0010111010",  -- INDEX 186
	B"11001001" when B"0010111011",  -- INDEX 187
	B"11111010" when B"0010111100",  -- INDEX 188
	B"00101100" when B"0010111101",  -- INDEX 189
	B"01010111" when B"0010111110",  -- INDEX 190
	B"01110100" when B"0010111111",  -- INDEX 191
	B"01111111" when B"0011000000",  -- INDEX 192
	B"01111000" when B"0011000001",  -- INDEX 193
	B"01011101" when B"0011000010",  -- INDEX 194
	B"00110100" when B"0011000011",  -- INDEX 195
	B"00000010" when B"0011000100",  -- INDEX 196
	B"11010001" when B"0011000101",  -- INDEX 197
	B"10100111" when B"0011000110",  -- INDEX 198
	B"10001010" when B"0011000111",  -- INDEX 199
	B"10000000" when B"0011001000",  -- INDEX 200
	B"10001010" when B"0011001001",  -- INDEX 201
	B"10100110" when B"0011001010",  -- INDEX 202
	B"11010000" when B"0011001011",  -- INDEX 203
	B"00000001" when B"0011001100",  -- INDEX 204
	B"00110011" when B"0011001101",  -- INDEX 205
	B"01011100" when B"0011001110",  -- INDEX 206
	B"01110111" when B"0011001111",  -- INDEX 207
	B"01111111" when B"0011010000",  -- INDEX 208
	B"01110101" when B"0011010001",  -- INDEX 209
	B"01010111" when B"0011010010",  -- INDEX 210
	B"00101101" when B"0011010011",  -- INDEX 211
	B"11111011" when B"0011010100",  -- INDEX 212
	B"11001010" when B"0011010101",  -- INDEX 213
	B"10100001" when B"0011010110",  -- INDEX 214
	B"10000111" when B"0011010111",  -- INDEX 215
	B"10000000" when B"0011011000",  -- INDEX 216
	B"10001101" when B"0011011001",  -- INDEX 217
	B"10101011" when B"0011011010",  -- INDEX 218
	B"11010111" when B"0011011011",  -- INDEX 219
	B"00001001" when B"0011011100",  -- INDEX 220
	B"00111001" when B"0011011101",  -- INDEX 221
	B"01100001" when B"0011011110",  -- INDEX 222
	B"01111010" when B"0011011111",  -- INDEX 223
	B"01111111" when B"0011100000",  -- INDEX 224
	B"01110010" when B"0011100001",  -- INDEX 225
	B"01010010" when B"0011100010",  -- INDEX 226
	B"00100110" when B"0011100011",  -- INDEX 227
	B"11110100" when B"0011100100",  -- INDEX 228
	B"11000100" when B"0011100101",  -- INDEX 229
	B"10011101" when B"0011100110",  -- INDEX 230
	B"10000101" when B"0011100111",  -- INDEX 231
	B"10000001" when B"0011101000",  -- INDEX 232
	B"10010000" when B"0011101001",  -- INDEX 233
	B"10110000" when B"0011101010",  -- INDEX 234
	B"11011100" when B"0011101011",  -- INDEX 235
	B"00001110" when B"0011101100",  -- INDEX 236
	B"00111110" when B"0011101101",  -- INDEX 237
	B"01100101" when B"0011101110",  -- INDEX 238
	B"01111011" when B"0011101111",  -- INDEX 239
	B"01111111" when B"0011110000",  -- INDEX 240
	B"01101111" when B"0011110001",  -- INDEX 241
	B"01001110" when B"0011110010",  -- INDEX 242
	B"00100001" when B"0011110011",  -- INDEX 243
	B"11101111" when B"0011110100",  -- INDEX 244
	B"11000000" when B"0011110101",  -- INDEX 245
	B"10011010" when B"0011110110",  -- INDEX 246
	B"10000100" when B"0011110111",  -- INDEX 247
	B"10000001" when B"0011111000",  -- INDEX 248
	B"10010010" when B"0011111001",  -- INDEX 249
	B"10110011" when B"0011111010",  -- INDEX 250
	B"11100001" when B"0011111011",  -- INDEX 251
	B"00010011" when B"0011111100",  -- INDEX 252
	B"01000010" when B"0011111101",  -- INDEX 253
	B"01100111" when B"0011111110",  -- INDEX 254
	B"01111100" when B"0011111111",  -- INDEX 255
	B"01111110" when B"0100000000",  -- INDEX 256
	B"01101101" when B"0100000001",  -- INDEX 257
	B"01001011" when B"0100000010",  -- INDEX 258
	B"00011101" when B"0100000011",  -- INDEX 259
	B"11101011" when B"0100000100",  -- INDEX 260
	B"10111100" when B"0100000101",  -- INDEX 261
	B"10011000" when B"0100000110",  -- INDEX 262
	B"10000011" when B"0100000111",  -- INDEX 263
	B"10000010" when B"0100001000",  -- INDEX 264
	B"10010100" when B"0100001001",  -- INDEX 265
	B"10110110" when B"0100001010",  -- INDEX 266
	B"11100100" when B"0100001011",  -- INDEX 267
	B"00010110" when B"0100001100",  -- INDEX 268
	B"01000101" when B"0100001101",  -- INDEX 269
	B"01101001" when B"0100001110",  -- INDEX 270
	B"01111101" when B"0100001111",  -- INDEX 271
	B"01111110" when B"0100010000",  -- INDEX 272
	B"01101100" when B"0100010001",  -- INDEX 273
	B"01001001" when B"0100010010",  -- INDEX 274
	B"00011011" when B"0100010011",  -- INDEX 275
	B"11101001" when B"0100010100",  -- INDEX 276
	B"10111010" when B"0100010101",  -- INDEX 277
	B"10010110" when B"0100010110",  -- INDEX 278
	B"10000011" when B"0100010111",  -- INDEX 279
	B"10000010" when B"0100011000",  -- INDEX 280
	B"10010101" when B"0100011001",  -- INDEX 281
	B"10111000" when B"0100011010",  -- INDEX 282
	B"11100110" when B"0100011011",  -- INDEX 283
	B"00011000" when B"0100011100",  -- INDEX 284
	B"01000110" when B"0100011101",  -- INDEX 285
	B"01101010" when B"0100011110",  -- INDEX 286
	B"01111101" when B"0100011111",  -- INDEX 287
	B"01111110" when B"0100100000",  -- INDEX 288
	B"01101011" when B"0100100001",  -- INDEX 289
	B"01001000" when B"0100100010",  -- INDEX 290
	B"00011001" when B"0100100011",  -- INDEX 291
	B"11100111" when B"0100100100",  -- INDEX 292
	B"10111001" when B"0100100101",  -- INDEX 293
	B"10010110" when B"0100100110",  -- INDEX 294
	B"10000011" when B"0100100111",  -- INDEX 295
	B"10000010" when B"0100101000",  -- INDEX 296
	B"10010101" when B"0100101001",  -- INDEX 297
	B"10111001" when B"0100101010",  -- INDEX 298
	B"11100111" when B"0100101011",  -- INDEX 299
	B"00011001" when B"0100101100",  -- INDEX 300
	B"01000111" when B"0100101101",  -- INDEX 301
	B"01101010" when B"0100101110",  -- INDEX 302
	B"01111101" when B"0100101111",  -- INDEX 303
	B"01111110" when B"0100110000",  -- INDEX 304
	B"01101011" when B"0100110001",  -- INDEX 305
	B"01000111" when B"0100110010",  -- INDEX 306
	B"00011001" when B"0100110011",  -- INDEX 307
	B"11100111" when B"0100110100",  -- INDEX 308
	B"10111001" when B"0100110101",  -- INDEX 309
	B"10010110" when B"0100110110",  -- INDEX 310
	B"10000011" when B"0100110111",  -- INDEX 311
	B"10000010" when B"0100111000",  -- INDEX 312
	B"10010101" when B"0100111001",  -- INDEX 313
	B"10111000" when B"0100111010",  -- INDEX 314
	B"11100110" when B"0100111011",  -- INDEX 315
	B"00011000" when B"0100111100",  -- INDEX 316
	B"01000110" when B"0100111101",  -- INDEX 317
	B"01101010" when B"0100111110",  -- INDEX 318
	B"01111101" when B"0100111111",  -- INDEX 319
	B"01111110" when B"0101000000",  -- INDEX 320
	B"01101011" when B"0101000001",  -- INDEX 321
	B"01001000" when B"0101000010",  -- INDEX 322
	B"00011010" when B"0101000011",  -- INDEX 323
	B"11101001" when B"0101000100",  -- INDEX 324
	B"10111010" when B"0101000101",  -- INDEX 325
	B"10010111" when B"0101000110",  -- INDEX 326
	B"10000011" when B"0101000111",  -- INDEX 327
	B"10000010" when B"0101001000",  -- INDEX 328
	B"10010100" when B"0101001001",  -- INDEX 329
	B"10110111" when B"0101001010",  -- INDEX 330
	B"11100100" when B"0101001011",  -- INDEX 331
	B"00010110" when B"0101001100",  -- INDEX 332
	B"01000101" when B"0101001101",  -- INDEX 333
	B"01101001" when B"0101001110",  -- INDEX 334
	B"01111101" when B"0101001111",  -- INDEX 335
	B"01111110" when B"0101010000",  -- INDEX 336
	B"01101100" when B"0101010001",  -- INDEX 337
	B"01001010" when B"0101010010",  -- INDEX 338
	B"00011101" when B"0101010011",  -- INDEX 339
	B"11101011" when B"0101010100",  -- INDEX 340
	B"10111101" when B"0101010101",  -- INDEX 341
	B"10011000" when B"0101010110",  -- INDEX 342
	B"10000011" when B"0101010111",  -- INDEX 343
	B"10000010" when B"0101011000",  -- INDEX 344
	B"10010011" when B"0101011001",  -- INDEX 345
	B"10110100" when B"0101011010",  -- INDEX 346
	B"11100001" when B"0101011011",  -- INDEX 347
	B"00010011" when B"0101011100",  -- INDEX 348
	B"01000010" when B"0101011101",  -- INDEX 349
	B"01100111" when B"0101011110",  -- INDEX 350
	B"01111100" when B"0101011111",  -- INDEX 351
	B"01111111" when B"0101100000",  -- INDEX 352
	B"01101110" when B"0101100001",  -- INDEX 353
	B"01001101" when B"0101100010",  -- INDEX 354
	B"00100000" when B"0101100011",  -- INDEX 355
	B"11101111" when B"0101100100",  -- INDEX 356
	B"11000000" when B"0101100101",  -- INDEX 357
	B"10011011" when B"0101100110",  -- INDEX 358
	B"10000100" when B"0101100111",  -- INDEX 359
	B"10000001" when B"0101101000",  -- INDEX 360
	B"10010001" when B"0101101001",  -- INDEX 361
	B"10110001" when B"0101101010",  -- INDEX 362
	B"11011101" when B"0101101011",  -- INDEX 363
	B"00001111" when B"0101101100",  -- INDEX 364
	B"00111110" when B"0101101101",  -- INDEX 365
	B"01100100" when B"0101101110",  -- INDEX 366
	B"01111011" when B"0101101111",  -- INDEX 367
	B"01111111" when B"0101110000",  -- INDEX 368
	B"01110001" when B"0101110001",  -- INDEX 369
	B"01010001" when B"0101110010",  -- INDEX 370
	B"00100101" when B"0101110011",  -- INDEX 371
	B"11110100" when B"0101110100",  -- INDEX 372
	B"11000100" when B"0101110101",  -- INDEX 373
	B"10011110" when B"0101110110",  -- INDEX 374
	B"10000110" when B"0101110111",  -- INDEX 375
	B"10000000" when B"0101111000",  -- INDEX 376
	B"10001110" when B"0101111001",  -- INDEX 377
	B"10101101" when B"0101111010",  -- INDEX 378
	B"11011000" when B"0101111011",  -- INDEX 379
	B"00001001" when B"0101111100",  -- INDEX 380
	B"00111001" when B"0101111101",  -- INDEX 381
	B"01100000" when B"0101111110",  -- INDEX 382
	B"01111001" when B"0101111111",  -- INDEX 383
	B"01111111" when B"0110000000",  -- INDEX 384
	B"01110011" when B"0110000001",  -- INDEX 385
	B"01010110" when B"0110000010",  -- INDEX 386
	B"00101011" when B"0110000011",  -- INDEX 387
	B"11111010" when B"0110000100",  -- INDEX 388
	B"11001010" when B"0110000101",  -- INDEX 389
	B"10100010" when B"0110000110",  -- INDEX 390
	B"10001000" when B"0110000111",  -- INDEX 391
	B"10000000" when B"0110001000",  -- INDEX 392
	B"10001011" when B"0110001001",  -- INDEX 393
	B"10101000" when B"0110001010",  -- INDEX 394
	B"11010001" when B"0110001011",  -- INDEX 395
	B"00000010" when B"0110001100",  -- INDEX 396
	B"00110010" when B"0110001101",  -- INDEX 397
	B"01011011" when B"0110001110",  -- INDEX 398
	B"01110110" when B"0110001111",  -- INDEX 399
	B"01111111" when B"0110010000",  -- INDEX 400
	B"01110110" when B"0110010001",  -- INDEX 401
	B"01011011" when B"0110010010",  -- INDEX 402
	B"00110010" when B"0110010011",  -- INDEX 403
	B"00000010" when B"0110010100",  -- INDEX 404
	B"11010001" when B"0110010101",  -- INDEX 405
	B"10101000" when B"0110010110",  -- INDEX 406
	B"10001011" when B"0110010111",  -- INDEX 407
	B"10000000" when B"0110011000",  -- INDEX 408
	B"10001000" when B"0110011001",  -- INDEX 409
	B"10100010" when B"0110011010",  -- INDEX 410
	B"11001010" when B"0110011011",  -- INDEX 411
	B"11111010" when B"0110011100",  -- INDEX 412
	B"00101011" when B"0110011101",  -- INDEX 413
	B"01010110" when B"0110011110",  -- INDEX 414
	B"01110011" when B"0110011111",  -- INDEX 415
	B"01111111" when B"0110100000",  -- INDEX 416
	B"01111001" when B"0110100001",  -- INDEX 417
	B"01100000" when B"0110100010",  -- INDEX 418
	B"00111001" when B"0110100011",  -- INDEX 419
	B"00001001" when B"0110100100",  -- INDEX 420
	B"11011000" when B"0110100101",  -- INDEX 421
	B"10101101" when B"0110100110",  -- INDEX 422
	B"10001110" when B"0110100111",  -- INDEX 423
	B"10000000" when B"0110101000",  -- INDEX 424
	B"10000110" when B"0110101001",  -- INDEX 425
	B"10011110" when B"0110101010",  -- INDEX 426
	B"11000100" when B"0110101011",  -- INDEX 427
	B"11110100" when B"0110101100",  -- INDEX 428
	B"00100101" when B"0110101101",  -- INDEX 429
	B"01010001" when B"0110101110",  -- INDEX 430
	B"01110001" when B"0110101111",  -- INDEX 431
	B"01111111" when B"0110110000",  -- INDEX 432
	B"01111011" when B"0110110001",  -- INDEX 433
	B"01100100" when B"0110110010",  -- INDEX 434
	B"00111110" when B"0110110011",  -- INDEX 435
	B"00001111" when B"0110110100",  -- INDEX 436
	B"11011101" when B"0110110101",  -- INDEX 437
	B"10110001" when B"0110110110",  -- INDEX 438
	B"10010001" when B"0110110111",  -- INDEX 439
	B"10000001" when B"0110111000",  -- INDEX 440
	B"10000100" when B"0110111001",  -- INDEX 441
	B"10011010" when B"0110111010",  -- INDEX 442
	B"11000000" when B"0110111011",  -- INDEX 443
	B"11101111" when B"0110111100",  -- INDEX 444
	B"00100000" when B"0110111101",  -- INDEX 445
	B"01001101" when B"0110111110",  -- INDEX 446
	B"01101110" when B"0110111111",  -- INDEX 447
	B"01111111" when B"0111000000",  -- INDEX 448
	B"01111100" when B"0111000001",  -- INDEX 449
	B"01100111" when B"0111000010",  -- INDEX 450
	B"01000010" when B"0111000011",  -- INDEX 451
	B"00010011" when B"0111000100",  -- INDEX 452
	B"11100010" when B"0111000101",  -- INDEX 453
	B"10110101" when B"0111000110",  -- INDEX 454
	B"10010011" when B"0111000111",  -- INDEX 455
	B"10000010" when B"0111001000",  -- INDEX 456
	B"10000011" when B"0111001001",  -- INDEX 457
	B"10011000" when B"0111001010",  -- INDEX 458
	B"10111100" when B"0111001011",  -- INDEX 459
	B"11101011" when B"0111001100",  -- INDEX 460
	B"00011101" when B"0111001101",  -- INDEX 461
	B"01001010" when B"0111001110",  -- INDEX 462
	B"01101100" when B"0111001111",  -- INDEX 463
	B"01111110" when B"0111010000",  -- INDEX 464
	B"01111101" when B"0111010001",  -- INDEX 465
	B"01101001" when B"0111010010",  -- INDEX 466
	B"01000101" when B"0111010011",  -- INDEX 467
	B"00010111" when B"0111010100",  -- INDEX 468
	B"11100101" when B"0111010101",  -- INDEX 469
	B"10110111" when B"0111010110",  -- INDEX 470
	B"10010101" when B"0111010111",  -- INDEX 471
	B"10000010" when B"0111011000",  -- INDEX 472
	B"10000011" when B"0111011001",  -- INDEX 473
	B"10010110" when B"0111011010",  -- INDEX 474
	B"10111010" when B"0111011011",  -- INDEX 475
	B"11101000" when B"0111011100",  -- INDEX 476
	B"00011010" when B"0111011101",  -- INDEX 477
	B"01001000" when B"0111011110",  -- INDEX 478
	B"01101011" when B"0111011111",  -- INDEX 479
	B"01111110" when B"0111100000",  -- INDEX 480
	B"01111101" when B"0111100001",  -- INDEX 481
	B"01101010" when B"0111100010",  -- INDEX 482
	B"01000111" when B"0111100011",  -- INDEX 483
	B"00011001" when B"0111100100",  -- INDEX 484
	B"11100111" when B"0111100101",  -- INDEX 485
	B"10111001" when B"0111100110",  -- INDEX 486
	B"10010101" when B"0111100111",  -- INDEX 487
	B"10000010" when B"0111101000",  -- INDEX 488
	B"10000010" when B"0111101001",  -- INDEX 489
	B"10010110" when B"0111101010",  -- INDEX 490
	B"10111001" when B"0111101011",  -- INDEX 491
	B"11100111" when B"0111101100",  -- INDEX 492
	B"00011001" when B"0111101101",  -- INDEX 493
	B"01000111" when B"0111101110",  -- INDEX 494
	B"01101010" when B"0111101111",  -- INDEX 495
	B"01111110" when B"0111110000",  -- INDEX 496
	B"01111110" when B"0111110001",  -- INDEX 497
	B"01101011" when B"0111110010",  -- INDEX 498
	B"01000111" when B"0111110011",  -- INDEX 499
	B"00011001" when B"0111110100",  -- INDEX 500
	B"11100111" when B"0111110101",  -- INDEX 501
	B"10111001" when B"0111110110",  -- INDEX 502
	B"10010110" when B"0111110111",  -- INDEX 503
	B"10000011" when B"0111111000",  -- INDEX 504
	B"10000010" when B"0111111001",  -- INDEX 505
	B"10010101" when B"0111111010",  -- INDEX 506
	B"10111001" when B"0111111011",  -- INDEX 507
	B"11100111" when B"0111111100",  -- INDEX 508
	B"00011001" when B"0111111101",  -- INDEX 509
	B"01000111" when B"0111111110",  -- INDEX 510
	B"01101010" when B"0111111111",  -- INDEX 511
	B"01111110" when B"1000000000",  -- INDEX 512
	B"01111110" when B"1000000001",  -- INDEX 513
	B"01101010" when B"1000000010",  -- INDEX 514
	B"01000111" when B"1000000011",  -- INDEX 515
	B"00011001" when B"1000000100",  -- INDEX 516
	B"11100111" when B"1000000101",  -- INDEX 517
	B"10111000" when B"1000000110",  -- INDEX 518
	B"10010101" when B"1000000111",  -- INDEX 519
	B"10000010" when B"1000001000",  -- INDEX 520
	B"10000011" when B"1000001001",  -- INDEX 521
	B"10010110" when B"1000001010",  -- INDEX 522
	B"10111010" when B"1000001011",  -- INDEX 523
	B"11101000" when B"1000001100",  -- INDEX 524
	B"00011010" when B"1000001101",  -- INDEX 525
	B"01001000" when B"1000001110",  -- INDEX 526
	B"01101011" when B"1000001111",  -- INDEX 527
	B"01111110" when B"1000010000",  -- INDEX 528
	B"01111101" when B"1000010001",  -- INDEX 529
	B"01101001" when B"1000010010",  -- INDEX 530
	B"01000101" when B"1000010011",  -- INDEX 531
	B"00010111" when B"1000010100",  -- INDEX 532
	B"11100101" when B"1000010101",  -- INDEX 533
	B"10110111" when B"1000010110",  -- INDEX 534
	B"10010100" when B"1000010111",  -- INDEX 535
	B"10000010" when B"1000011000",  -- INDEX 536
	B"10000011" when B"1000011001",  -- INDEX 537
	B"10010111" when B"1000011010",  -- INDEX 538
	B"10111100" when B"1000011011",  -- INDEX 539
	B"11101011" when B"1000011100",  -- INDEX 540
	B"00011101" when B"1000011101",  -- INDEX 541
	B"01001010" when B"1000011110",  -- INDEX 542
	B"01101101" when B"1000011111",  -- INDEX 543
	B"01111110" when B"1000100000",  -- INDEX 544
	B"01111101" when B"1000100001",  -- INDEX 545
	B"01101000" when B"1000100010",  -- INDEX 546
	B"01000011" when B"1000100011",  -- INDEX 547
	B"00010100" when B"1000100100",  -- INDEX 548
	B"11100010" when B"1000100101",  -- INDEX 549
	B"10110100" when B"1000100110",  -- INDEX 550
	B"10010010" when B"1000100111",  -- INDEX 551
	B"10000001" when B"1000101000",  -- INDEX 552
	B"10000100" when B"1000101001",  -- INDEX 553
	B"10011010" when B"1000101010",  -- INDEX 554
	B"10111111" when B"1000101011",  -- INDEX 555
	B"11101110" when B"1000101100",  -- INDEX 556
	B"00100001" when B"1000101101",  -- INDEX 557
	B"01001110" when B"1000101110",  -- INDEX 558
	B"01101111" when B"1000101111",  -- INDEX 559
	B"01111111" when B"1000110000",  -- INDEX 560
	B"01111011" when B"1000110001",  -- INDEX 561
	B"01100101" when B"1000110010",  -- INDEX 562
	B"00111111" when B"1000110011",  -- INDEX 563
	B"00001111" when B"1000110100",  -- INDEX 564
	B"11011101" when B"1000110101",  -- INDEX 565
	B"10110000" when B"1000110110",  -- INDEX 566
	B"10010000" when B"1000110111",  -- INDEX 567
	B"10000001" when B"1000111000",  -- INDEX 568
	B"10000101" when B"1000111001",  -- INDEX 569
	B"10011101" when B"1000111010",  -- INDEX 570
	B"11000011" when B"1000111011",  -- INDEX 571
	B"11110011" when B"1000111100",  -- INDEX 572
	B"00100110" when B"1000111101",  -- INDEX 573
	B"01010010" when B"1000111110",  -- INDEX 574
	B"01110001" when B"1000111111",  -- INDEX 575
	B"01111111" when B"1001000000",  -- INDEX 576
	B"01111010" when B"1001000001",  -- INDEX 577
	B"01100001" when B"1001000010",  -- INDEX 578
	B"00111010" when B"1001000011",  -- INDEX 579
	B"00001001" when B"1001000100",  -- INDEX 580
	B"11011000" when B"1001000101",  -- INDEX 581
	B"10101100" when B"1001000110",  -- INDEX 582
	B"10001101" when B"1001000111",  -- INDEX 583
	B"10000000" when B"1001001000",  -- INDEX 584
	B"10000111" when B"1001001001",  -- INDEX 585
	B"10100001" when B"1001001010",  -- INDEX 586
	B"11001001" when B"1001001011",  -- INDEX 587
	B"11111010" when B"1001001100",  -- INDEX 588
	B"00101100" when B"1001001101",  -- INDEX 589
	B"01010111" when B"1001001110",  -- INDEX 590
	B"01110100" when B"1001001111",  -- INDEX 591
	B"01111111" when B"1001010000",  -- INDEX 592
	B"01111000" when B"1001010001",  -- INDEX 593
	B"01011101" when B"1001010010",  -- INDEX 594
	B"00110100" when B"1001010011",  -- INDEX 595
	B"00000010" when B"1001010100",  -- INDEX 596
	B"11010001" when B"1001010101",  -- INDEX 597
	B"10100111" when B"1001010110",  -- INDEX 598
	B"10001010" when B"1001010111",  -- INDEX 599
	B"10000000" when B"1001011000",  -- INDEX 600
	B"10001010" when B"1001011001",  -- INDEX 601
	B"10100110" when B"1001011010",  -- INDEX 602
	B"11010000" when B"1001011011",  -- INDEX 603
	B"00000001" when B"1001011100",  -- INDEX 604
	B"00110011" when B"1001011101",  -- INDEX 605
	B"01011100" when B"1001011110",  -- INDEX 606
	B"01110111" when B"1001011111",  -- INDEX 607
	B"01111111" when B"1001100000",  -- INDEX 608
	B"01110101" when B"1001100001",  -- INDEX 609
	B"01010111" when B"1001100010",  -- INDEX 610
	B"00101101" when B"1001100011",  -- INDEX 611
	B"11111011" when B"1001100100",  -- INDEX 612
	B"11001010" when B"1001100101",  -- INDEX 613
	B"10100001" when B"1001100110",  -- INDEX 614
	B"10000111" when B"1001100111",  -- INDEX 615
	B"10000000" when B"1001101000",  -- INDEX 616
	B"10001101" when B"1001101001",  -- INDEX 617
	B"10101011" when B"1001101010",  -- INDEX 618
	B"11010111" when B"1001101011",  -- INDEX 619
	B"00001001" when B"1001101100",  -- INDEX 620
	B"00111001" when B"1001101101",  -- INDEX 621
	B"01100001" when B"1001101110",  -- INDEX 622
	B"01111010" when B"1001101111",  -- INDEX 623
	B"01111111" when B"1001110000",  -- INDEX 624
	B"01110010" when B"1001110001",  -- INDEX 625
	B"01010010" when B"1001110010",  -- INDEX 626
	B"00100110" when B"1001110011",  -- INDEX 627
	B"11110100" when B"1001110100",  -- INDEX 628
	B"11000100" when B"1001110101",  -- INDEX 629
	B"10011101" when B"1001110110",  -- INDEX 630
	B"10000101" when B"1001110111",  -- INDEX 631
	B"10000001" when B"1001111000",  -- INDEX 632
	B"10010000" when B"1001111001",  -- INDEX 633
	B"10110000" when B"1001111010",  -- INDEX 634
	B"11011100" when B"1001111011",  -- INDEX 635
	B"00001110" when B"1001111100",  -- INDEX 636
	B"00111110" when B"1001111101",  -- INDEX 637
	B"01100101" when B"1001111110",  -- INDEX 638
	B"01111011" when B"1001111111",  -- INDEX 639
	B"01111111" when B"1010000000",  -- INDEX 640
	B"01101111" when B"1010000001",  -- INDEX 641
	B"01001110" when B"1010000010",  -- INDEX 642
	B"00100001" when B"1010000011",  -- INDEX 643
	B"11101111" when B"1010000100",  -- INDEX 644
	B"11000000" when B"1010000101",  -- INDEX 645
	B"10011010" when B"1010000110",  -- INDEX 646
	B"10000100" when B"1010000111",  -- INDEX 647
	B"10000001" when B"1010001000",  -- INDEX 648
	B"10010010" when B"1010001001",  -- INDEX 649
	B"10110011" when B"1010001010",  -- INDEX 650
	B"11100001" when B"1010001011",  -- INDEX 651
	B"00010011" when B"1010001100",  -- INDEX 652
	B"01000010" when B"1010001101",  -- INDEX 653
	B"01100111" when B"1010001110",  -- INDEX 654
	B"01111100" when B"1010001111",  -- INDEX 655
	B"01111110" when B"1010010000",  -- INDEX 656
	B"01101101" when B"1010010001",  -- INDEX 657
	B"01001011" when B"1010010010",  -- INDEX 658
	B"00011101" when B"1010010011",  -- INDEX 659
	B"11101011" when B"1010010100",  -- INDEX 660
	B"10111100" when B"1010010101",  -- INDEX 661
	B"10011000" when B"1010010110",  -- INDEX 662
	B"10000011" when B"1010010111",  -- INDEX 663
	B"10000010" when B"1010011000",  -- INDEX 664
	B"10010100" when B"1010011001",  -- INDEX 665
	B"10110110" when B"1010011010",  -- INDEX 666
	B"11100100" when B"1010011011",  -- INDEX 667
	B"00010110" when B"1010011100",  -- INDEX 668
	B"01000101" when B"1010011101",  -- INDEX 669
	B"01101001" when B"1010011110",  -- INDEX 670
	B"01111101" when B"1010011111",  -- INDEX 671
	B"01111110" when B"1010100000",  -- INDEX 672
	B"01101100" when B"1010100001",  -- INDEX 673
	B"01001001" when B"1010100010",  -- INDEX 674
	B"00011011" when B"1010100011",  -- INDEX 675
	B"11101001" when B"1010100100",  -- INDEX 676
	B"10111010" when B"1010100101",  -- INDEX 677
	B"10010110" when B"1010100110",  -- INDEX 678
	B"10000011" when B"1010100111",  -- INDEX 679
	B"10000010" when B"1010101000",  -- INDEX 680
	B"10010101" when B"1010101001",  -- INDEX 681
	B"10111000" when B"1010101010",  -- INDEX 682
	B"11100110" when B"1010101011",  -- INDEX 683
	B"00011000" when B"1010101100",  -- INDEX 684
	B"01000110" when B"1010101101",  -- INDEX 685
	B"01101010" when B"1010101110",  -- INDEX 686
	B"01111101" when B"1010101111",  -- INDEX 687
	B"01111110" when B"1010110000",  -- INDEX 688
	B"01101011" when B"1010110001",  -- INDEX 689
	B"01001000" when B"1010110010",  -- INDEX 690
	B"00011001" when B"1010110011",  -- INDEX 691
	B"11100111" when B"1010110100",  -- INDEX 692
	B"10111001" when B"1010110101",  -- INDEX 693
	B"10010110" when B"1010110110",  -- INDEX 694
	B"10000011" when B"1010110111",  -- INDEX 695
	B"10000010" when B"1010111000",  -- INDEX 696
	B"10010101" when B"1010111001",  -- INDEX 697
	B"10111001" when B"1010111010",  -- INDEX 698
	B"11100111" when B"1010111011",  -- INDEX 699
	B"00011001" when B"1010111100",  -- INDEX 700
	B"01000111" when B"1010111101",  -- INDEX 701
	B"01101010" when B"1010111110",  -- INDEX 702
	B"01111101" when B"1010111111",  -- INDEX 703
	B"01111110" when B"1011000000",  -- INDEX 704
	B"01101011" when B"1011000001",  -- INDEX 705
	B"01000111" when B"1011000010",  -- INDEX 706
	B"00011001" when B"1011000011",  -- INDEX 707
	B"11100111" when B"1011000100",  -- INDEX 708
	B"10111001" when B"1011000101",  -- INDEX 709
	B"10010110" when B"1011000110",  -- INDEX 710
	B"10000011" when B"1011000111",  -- INDEX 711
	B"10000010" when B"1011001000",  -- INDEX 712
	B"10010101" when B"1011001001",  -- INDEX 713
	B"10111000" when B"1011001010",  -- INDEX 714
	B"11100110" when B"1011001011",  -- INDEX 715
	B"00011000" when B"1011001100",  -- INDEX 716
	B"01000110" when B"1011001101",  -- INDEX 717
	B"01101010" when B"1011001110",  -- INDEX 718
	B"01111101" when B"1011001111",  -- INDEX 719
	B"01111110" when B"1011010000",  -- INDEX 720
	B"01101011" when B"1011010001",  -- INDEX 721
	B"01001000" when B"1011010010",  -- INDEX 722
	B"00011010" when B"1011010011",  -- INDEX 723
	B"11101001" when B"1011010100",  -- INDEX 724
	B"10111010" when B"1011010101",  -- INDEX 725
	B"10010111" when B"1011010110",  -- INDEX 726
	B"10000011" when B"1011010111",  -- INDEX 727
	B"10000010" when B"1011011000",  -- INDEX 728
	B"10010100" when B"1011011001",  -- INDEX 729
	B"10110111" when B"1011011010",  -- INDEX 730
	B"11100100" when B"1011011011",  -- INDEX 731
	B"00010110" when B"1011011100",  -- INDEX 732
	B"01000101" when B"1011011101",  -- INDEX 733
	B"01101001" when B"1011011110",  -- INDEX 734
	B"01111101" when B"1011011111",  -- INDEX 735
	B"01111110" when B"1011100000",  -- INDEX 736
	B"01101100" when B"1011100001",  -- INDEX 737
	B"01001010" when B"1011100010",  -- INDEX 738
	B"00011101" when B"1011100011",  -- INDEX 739
	B"11101011" when B"1011100100",  -- INDEX 740
	B"10111101" when B"1011100101",  -- INDEX 741
	B"10011000" when B"1011100110",  -- INDEX 742
	B"10000011" when B"1011100111",  -- INDEX 743
	B"10000010" when B"1011101000",  -- INDEX 744
	B"10010011" when B"1011101001",  -- INDEX 745
	B"10110100" when B"1011101010",  -- INDEX 746
	B"11100001" when B"1011101011",  -- INDEX 747
	B"00010011" when B"1011101100",  -- INDEX 748
	B"01000010" when B"1011101101",  -- INDEX 749
	B"01100111" when B"1011101110",  -- INDEX 750
	B"01111100" when B"1011101111",  -- INDEX 751
	B"01111111" when B"1011110000",  -- INDEX 752
	B"01101110" when B"1011110001",  -- INDEX 753
	B"01001101" when B"1011110010",  -- INDEX 754
	B"00100000" when B"1011110011",  -- INDEX 755
	B"11101111" when B"1011110100",  -- INDEX 756
	B"11000000" when B"1011110101",  -- INDEX 757
	B"10011011" when B"1011110110",  -- INDEX 758
	B"10000100" when B"1011110111",  -- INDEX 759
	B"10000001" when B"1011111000",  -- INDEX 760
	B"10010001" when B"1011111001",  -- INDEX 761
	B"10110001" when B"1011111010",  -- INDEX 762
	B"11011101" when B"1011111011",  -- INDEX 763
	B"00001111" when B"1011111100",  -- INDEX 764
	B"00111110" when B"1011111101",  -- INDEX 765
	B"01100100" when B"1011111110",  -- INDEX 766
	B"01111011" when B"1011111111",  -- INDEX 767
	B"01111111" when B"1100000000",  -- INDEX 768
	B"01110001" when B"1100000001",  -- INDEX 769
	B"01010001" when B"1100000010",  -- INDEX 770
	B"00100101" when B"1100000011",  -- INDEX 771
	B"11110100" when B"1100000100",  -- INDEX 772
	B"11000100" when B"1100000101",  -- INDEX 773
	B"10011110" when B"1100000110",  -- INDEX 774
	B"10000110" when B"1100000111",  -- INDEX 775
	B"10000000" when B"1100001000",  -- INDEX 776
	B"10001110" when B"1100001001",  -- INDEX 777
	B"10101101" when B"1100001010",  -- INDEX 778
	B"11011000" when B"1100001011",  -- INDEX 779
	B"00001001" when B"1100001100",  -- INDEX 780
	B"00111001" when B"1100001101",  -- INDEX 781
	B"01100000" when B"1100001110",  -- INDEX 782
	B"01111001" when B"1100001111",  -- INDEX 783
	B"01111111" when B"1100010000",  -- INDEX 784
	B"01110011" when B"1100010001",  -- INDEX 785
	B"01010110" when B"1100010010",  -- INDEX 786
	B"00101011" when B"1100010011",  -- INDEX 787
	B"11111010" when B"1100010100",  -- INDEX 788
	B"11001010" when B"1100010101",  -- INDEX 789
	B"10100010" when B"1100010110",  -- INDEX 790
	B"10001000" when B"1100010111",  -- INDEX 791
	B"10000000" when B"1100011000",  -- INDEX 792
	B"10001011" when B"1100011001",  -- INDEX 793
	B"10101000" when B"1100011010",  -- INDEX 794
	B"11010001" when B"1100011011",  -- INDEX 795
	B"00000010" when B"1100011100",  -- INDEX 796
	B"00110010" when B"1100011101",  -- INDEX 797
	B"01011011" when B"1100011110",  -- INDEX 798
	B"01110110" when B"1100011111",  -- INDEX 799
	B"01111111" when B"1100100000",  -- INDEX 800
	B"01110110" when B"1100100001",  -- INDEX 801
	B"01011011" when B"1100100010",  -- INDEX 802
	B"00110010" when B"1100100011",  -- INDEX 803
	B"00000010" when B"1100100100",  -- INDEX 804
	B"11010001" when B"1100100101",  -- INDEX 805
	B"10101000" when B"1100100110",  -- INDEX 806
	B"10001011" when B"1100100111",  -- INDEX 807
	B"10000000" when B"1100101000",  -- INDEX 808
	B"10001000" when B"1100101001",  -- INDEX 809
	B"10100010" when B"1100101010",  -- INDEX 810
	B"11001010" when B"1100101011",  -- INDEX 811
	B"11111010" when B"1100101100",  -- INDEX 812
	B"00101011" when B"1100101101",  -- INDEX 813
	B"01010110" when B"1100101110",  -- INDEX 814
	B"01110011" when B"1100101111",  -- INDEX 815
	B"01111111" when B"1100110000",  -- INDEX 816
	B"01111001" when B"1100110001",  -- INDEX 817
	B"01100000" when B"1100110010",  -- INDEX 818
	B"00111001" when B"1100110011",  -- INDEX 819
	B"00001001" when B"1100110100",  -- INDEX 820
	B"11011000" when B"1100110101",  -- INDEX 821
	B"10101101" when B"1100110110",  -- INDEX 822
	B"10001110" when B"1100110111",  -- INDEX 823
	B"10000000" when B"1100111000",  -- INDEX 824
	B"10000110" when B"1100111001",  -- INDEX 825
	B"10011110" when B"1100111010",  -- INDEX 826
	B"11000100" when B"1100111011",  -- INDEX 827
	B"11110100" when B"1100111100",  -- INDEX 828
	B"00100101" when B"1100111101",  -- INDEX 829
	B"01010001" when B"1100111110",  -- INDEX 830
	B"01110001" when B"1100111111",  -- INDEX 831
	B"01111111" when B"1101000000",  -- INDEX 832
	B"01111011" when B"1101000001",  -- INDEX 833
	B"01100100" when B"1101000010",  -- INDEX 834
	B"00111110" when B"1101000011",  -- INDEX 835
	B"00001111" when B"1101000100",  -- INDEX 836
	B"11011101" when B"1101000101",  -- INDEX 837
	B"10110001" when B"1101000110",  -- INDEX 838
	B"10010001" when B"1101000111",  -- INDEX 839
	B"10000001" when B"1101001000",  -- INDEX 840
	B"10000100" when B"1101001001",  -- INDEX 841
	B"10011010" when B"1101001010",  -- INDEX 842
	B"11000000" when B"1101001011",  -- INDEX 843
	B"11101111" when B"1101001100",  -- INDEX 844
	B"00100000" when B"1101001101",  -- INDEX 845
	B"01001101" when B"1101001110",  -- INDEX 846
	B"01101110" when B"1101001111",  -- INDEX 847
	B"01111111" when B"1101010000",  -- INDEX 848
	B"01111100" when B"1101010001",  -- INDEX 849
	B"01100111" when B"1101010010",  -- INDEX 850
	B"01000010" when B"1101010011",  -- INDEX 851
	B"00010011" when B"1101010100",  -- INDEX 852
	B"11100010" when B"1101010101",  -- INDEX 853
	B"10110101" when B"1101010110",  -- INDEX 854
	B"10010011" when B"1101010111",  -- INDEX 855
	B"10000010" when B"1101011000",  -- INDEX 856
	B"10000011" when B"1101011001",  -- INDEX 857
	B"10011000" when B"1101011010",  -- INDEX 858
	B"10111100" when B"1101011011",  -- INDEX 859
	B"11101011" when B"1101011100",  -- INDEX 860
	B"00011101" when B"1101011101",  -- INDEX 861
	B"01001010" when B"1101011110",  -- INDEX 862
	B"01101100" when B"1101011111",  -- INDEX 863
	B"01111110" when B"1101100000",  -- INDEX 864
	B"01111101" when B"1101100001",  -- INDEX 865
	B"01101001" when B"1101100010",  -- INDEX 866
	B"01000101" when B"1101100011",  -- INDEX 867
	B"00010111" when B"1101100100",  -- INDEX 868
	B"11100101" when B"1101100101",  -- INDEX 869
	B"10110111" when B"1101100110",  -- INDEX 870
	B"10010101" when B"1101100111",  -- INDEX 871
	B"10000010" when B"1101101000",  -- INDEX 872
	B"10000011" when B"1101101001",  -- INDEX 873
	B"10010110" when B"1101101010",  -- INDEX 874
	B"10111010" when B"1101101011",  -- INDEX 875
	B"11101000" when B"1101101100",  -- INDEX 876
	B"00011010" when B"1101101101",  -- INDEX 877
	B"01001000" when B"1101101110",  -- INDEX 878
	B"01101011" when B"1101101111",  -- INDEX 879
	B"01111110" when B"1101110000",  -- INDEX 880
	B"01111101" when B"1101110001",  -- INDEX 881
	B"01101010" when B"1101110010",  -- INDEX 882
	B"01000111" when B"1101110011",  -- INDEX 883
	B"00011001" when B"1101110100",  -- INDEX 884
	B"11100111" when B"1101110101",  -- INDEX 885
	B"10111001" when B"1101110110",  -- INDEX 886
	B"10010101" when B"1101110111",  -- INDEX 887
	B"10000010" when B"1101111000",  -- INDEX 888
	B"10000010" when B"1101111001",  -- INDEX 889
	B"10010110" when B"1101111010",  -- INDEX 890
	B"10111001" when B"1101111011",  -- INDEX 891
	B"11100111" when B"1101111100",  -- INDEX 892
	B"00011001" when B"1101111101",  -- INDEX 893
	B"01000111" when B"1101111110",  -- INDEX 894
	B"01101010" when B"1101111111",  -- INDEX 895
	B"01111110" when B"1110000000",  -- INDEX 896
	B"01111110" when B"1110000001",  -- INDEX 897
	B"01101011" when B"1110000010",  -- INDEX 898
	B"01000111" when B"1110000011",  -- INDEX 899
	B"00011001" when B"1110000100",  -- INDEX 900
	B"11100111" when B"1110000101",  -- INDEX 901
	B"10111001" when B"1110000110",  -- INDEX 902
	B"10010110" when B"1110000111",  -- INDEX 903
	B"10000011" when B"1110001000",  -- INDEX 904
	B"10000010" when B"1110001001",  -- INDEX 905
	B"10010101" when B"1110001010",  -- INDEX 906
	B"10111001" when B"1110001011",  -- INDEX 907
	B"11100111" when B"1110001100",  -- INDEX 908
	B"00011001" when B"1110001101",  -- INDEX 909
	B"01000111" when B"1110001110",  -- INDEX 910
	B"01101010" when B"1110001111",  -- INDEX 911
	B"01111110" when B"1110010000",  -- INDEX 912
	B"01111110" when B"1110010001",  -- INDEX 913
	B"01101010" when B"1110010010",  -- INDEX 914
	B"01000111" when B"1110010011",  -- INDEX 915
	B"00011001" when B"1110010100",  -- INDEX 916
	B"11100111" when B"1110010101",  -- INDEX 917
	B"10111000" when B"1110010110",  -- INDEX 918
	B"10010101" when B"1110010111",  -- INDEX 919
	B"10000010" when B"1110011000",  -- INDEX 920
	B"10000011" when B"1110011001",  -- INDEX 921
	B"10010110" when B"1110011010",  -- INDEX 922
	B"10111010" when B"1110011011",  -- INDEX 923
	B"11101000" when B"1110011100",  -- INDEX 924
	B"00011010" when B"1110011101",  -- INDEX 925
	B"01001000" when B"1110011110",  -- INDEX 926
	B"01101011" when B"1110011111",  -- INDEX 927
	B"01111110" when B"1110100000",  -- INDEX 928
	B"01111101" when B"1110100001",  -- INDEX 929
	B"01101001" when B"1110100010",  -- INDEX 930
	B"01000101" when B"1110100011",  -- INDEX 931
	B"00010111" when B"1110100100",  -- INDEX 932
	B"11100101" when B"1110100101",  -- INDEX 933
	B"10110111" when B"1110100110",  -- INDEX 934
	B"10010100" when B"1110100111",  -- INDEX 935
	B"10000010" when B"1110101000",  -- INDEX 936
	B"10000011" when B"1110101001",  -- INDEX 937
	B"10010111" when B"1110101010",  -- INDEX 938
	B"10111100" when B"1110101011",  -- INDEX 939
	B"11101011" when B"1110101100",  -- INDEX 940
	B"00011101" when B"1110101101",  -- INDEX 941
	B"01001010" when B"1110101110",  -- INDEX 942
	B"01101101" when B"1110101111",  -- INDEX 943
	B"01111110" when B"1110110000",  -- INDEX 944
	B"01111101" when B"1110110001",  -- INDEX 945
	B"01101000" when B"1110110010",  -- INDEX 946
	B"01000011" when B"1110110011",  -- INDEX 947
	B"00010100" when B"1110110100",  -- INDEX 948
	B"11100010" when B"1110110101",  -- INDEX 949
	B"10110100" when B"1110110110",  -- INDEX 950
	B"10010010" when B"1110110111",  -- INDEX 951
	B"10000001" when B"1110111000",  -- INDEX 952
	B"10000100" when B"1110111001",  -- INDEX 953
	B"10011010" when B"1110111010",  -- INDEX 954
	B"10111111" when B"1110111011",  -- INDEX 955
	B"11101110" when B"1110111100",  -- INDEX 956
	B"00100001" when B"1110111101",  -- INDEX 957
	B"01001110" when B"1110111110",  -- INDEX 958
	B"01101111" when B"1110111111",  -- INDEX 959
	B"01111111" when B"1111000000",  -- INDEX 960
	B"01111011" when B"1111000001",  -- INDEX 961
	B"01100101" when B"1111000010",  -- INDEX 962
	B"00111111" when B"1111000011",  -- INDEX 963
	B"00001111" when B"1111000100",  -- INDEX 964
	B"11011101" when B"1111000101",  -- INDEX 965
	B"10110000" when B"1111000110",  -- INDEX 966
	B"10010000" when B"1111000111",  -- INDEX 967
	B"10000001" when B"1111001000",  -- INDEX 968
	B"10000101" when B"1111001001",  -- INDEX 969
	B"10011101" when B"1111001010",  -- INDEX 970
	B"11000011" when B"1111001011",  -- INDEX 971
	B"11110011" when B"1111001100",  -- INDEX 972
	B"00100110" when B"1111001101",  -- INDEX 973
	B"01010010" when B"1111001110",  -- INDEX 974
	B"01110001" when B"1111001111",  -- INDEX 975
	B"01111111" when B"1111010000",  -- INDEX 976
	B"01111010" when B"1111010001",  -- INDEX 977
	B"01100001" when B"1111010010",  -- INDEX 978
	B"00111010" when B"1111010011",  -- INDEX 979
	B"00001001" when B"1111010100",  -- INDEX 980
	B"11011000" when B"1111010101",  -- INDEX 981
	B"10101100" when B"1111010110",  -- INDEX 982
	B"10001101" when B"1111010111",  -- INDEX 983
	B"10000000" when B"1111011000",  -- INDEX 984
	B"10000111" when B"1111011001",  -- INDEX 985
	B"10100001" when B"1111011010",  -- INDEX 986
	B"11001001" when B"1111011011",  -- INDEX 987
	B"11111010" when B"1111011100",  -- INDEX 988
	B"00101100" when B"1111011101",  -- INDEX 989
	B"01010111" when B"1111011110",  -- INDEX 990
	B"01110100" when B"1111011111",  -- INDEX 991
	B"01111111" when B"1111100000",  -- INDEX 992
	B"01111000" when B"1111100001",  -- INDEX 993
	B"01011101" when B"1111100010",  -- INDEX 994
	B"00110100" when B"1111100011",  -- INDEX 995
	B"00000010" when B"1111100100",  -- INDEX 996
	B"11010001" when B"1111100101",  -- INDEX 997
	B"10100111" when B"1111100110",  -- INDEX 998
	B"10001010" when B"1111100111",  -- INDEX 999

-- END INPUT FM SIGNAL
	B"00000000" when others;

end input_data;
