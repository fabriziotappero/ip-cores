/*******************************************************************************
 *
 * top.v
 * Copyright 2012, Sinclair R.F., Inc.
 *
 * Top-level module for Conway's Game of Life design example.
 *
 ******************************************************************************/

module top(
);

/*******************************************************************************
 *
 * Instantiate the dual-port ping-pong memories.
 *
 ******************************************************************************/

reg [7:0] mema[8191:0];
reg [7:0] memb[8191:0];

/*******************************************************************************
 *
 * Generate the output NTSC video.
 *
 ******************************************************************************/

/*******************************************************************************
 *
 * Instantiate the SSBCC.9x8 micro controller.
 *
 ******************************************************************************/

endmodule
