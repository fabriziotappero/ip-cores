/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

module rom (clk, addr, out);
   input clk;
   input [8:0] addr;
   output reg [25:0] out;
   
   always @(posedge clk)
      case (addr)
         0: out <= 26'h30c042;
         1: out <= 26'h514045;
         2: out <= 26'h61a041;
         3: out <= 26'h71e041;
         4: out <= 26'hc046;
         5: out <= 26'h1603840;
         6: out <= 26'h1702041;
         7: out <= 26'h1717857;
         8: out <= 26'h1817847;
         9: out <= 26'h1963847;
         10: out <= 26'hf5d059;
         11: out <= 26'hf3d045;
         12: out <= 26'h1763845;
         13: out <= 26'h185f840;
         14: out <= 26'h161f856;
         15: out <= 26'h1160056;
         16: out <= 26'h1144051;
         17: out <= 26'h1214045;
         18: out <= 26'h131f840;
         19: out <= 26'h135d053;
         20: out <= 26'h1404041;
         21: out <= 26'h151c047;
         22: out <= 26'h3e041;
         23: out <= 26'h1646041;
         24: out <= 26'h174a041;
         25: out <= 26'h184e041;
         26: out <= 26'h1952041;
         27: out <= 26'h1a56041;
         28: out <= 26'hf00057;
         29: out <= 26'hf3c059;
         30: out <= 26'h1158058;
         31: out <= 26'h114405a;
         32: out <= 26'h1144051;
         33: out <= 26'h125d059;
         34: out <= 26'h1369058;
         35: out <= 26'h1464041;
         36: out <= 26'h156805a;
         37: out <= 26'h61a081;
         38: out <= 26'h619042;
         39: out <= 26'h71e081;
         40: out <= 26'h71c047;
         41: out <= 26'hc046;
         42: out <= 26'h1600040;
         43: out <= 26'h1717847;
         44: out <= 26'h5b840;
         45: out <= 26'h1800056;
         46: out <= 26'h1901056;
         47: out <= 26'h1a3c054;
         48: out <= 26'h1b68052;
         49: out <= 26'h1c69052;
         50: out <= 26'h1d3d054;
         51: out <= 26'h1e75053;
         52: out <= 26'h1d74053;
         53: out <= 26'h1f44055;
         54: out <= 26'h207c053;
         55: out <= 26'h217d053;
         56: out <= 26'h225c056;
         57: out <= 26'h165d056;
         58: out <= 26'h2345055;
         59: out <= 26'h248c052;
         60: out <= 26'h238d052;
         61: out <= 26'h2560057;
         62: out <= 26'h266c060;
         63: out <= 26'h2700062;
         64: out <= 26'h2878064;
         65: out <= 26'h2964057;
         66: out <= 26'h2a70061;
         67: out <= 26'h2b00056;
         68: out <= 26'h2c74063;
         69: out <= 26'h186385b;
         70: out <= 26'h1b97866;
         71: out <= 26'h205f860;
         72: out <= 26'h1e0385e;
         73: out <= 26'h259f868;
         74: out <= 26'h228b864;
         75: out <= 26'h196785c;
         76: out <= 26'h1ca786a;
         77: out <= 26'h175f861;
         78: out <= 26'h385d;
         79: out <= 26'h1daf86c;
         80: out <= 26'h165b863;
         81: out <= 26'h2160065;
         82: out <= 26'h238005d;
         83: out <= 26'h2481057;
         84: out <= 26'h2665058;
         85: out <= 26'h175c060;
         86: out <= 26'h1789057;
         87: out <= 26'h175c056;
         88: out <= 26'h1864058;
         89: out <= 26'h186105e;
         90: out <= 26'h1861040;
         91: out <= 26'h198d061;
         92: out <= 26'h196505e;
         93: out <= 26'h1664056;
         94: out <= 26'h1984063;
         95: out <= 26'h196505b;
         96: out <= 26'h1964062;
         97: out <= 26'h64040;
         98: out <= 26'h1990066;
         99: out <= 26'h1e91066;
         100: out <= 26'h1e7805c;
         101: out <= 26'h1e7905b;
         102: out <= 26'h205c058;
         103: out <= 26'h175d058;
         104: out <= 26'h175c05c;
         105: out <= 26'h175c05b;
         106: out <= 26'h175d065;
         107: out <= 26'h175d05d;
         108: out <= 26'hf59052;
         109: out <= 26'h1101053;
         110: out <= 26'h65052;
         111: out <= 26'h1054;
         112: out <= 26'h1679053;
         113: out <= 26'h1659055;
         114: out <= 26'h148105a;
         115: out <= 26'h155d05f;
         116: out <= 26'h1201041;
         117: out <= 26'h1359041;
         118: out <= 26'h93e041;
         119: out <= 26'h3c052;
         120: out <= 26'h54;
         121: out <= 26'h163f84f;
         122: out <= 26'h173f852;
         123: out <= 26'h184b854;
         124: out <= 26'h1953854;
         125: out <= 26'h3840;
         126: out <= 26'h175c058;
         127: out <= 26'h1859058;
         128: out <= 26'h1965057;
         129: out <= 26'h57;
         130: out <= 26'h1056;
         131: out <= 26'h1644053;
         132: out <= 26'h1658055;
         133: out <= 26'h1747851;
         134: out <= 26'h1a47853;
         135: out <= 26'h1b4f855;
         136: out <= 26'h1c57855;
         137: out <= 26'h165b856;
         138: out <= 26'h1a6805b;
         139: out <= 26'h1b5d05b;
         140: out <= 26'h1c7105a;
         141: out <= 26'h165805a;
         142: out <= 26'h1659057;
         143: out <= 26'h173c052;
         144: out <= 26'h1a3c054;
         145: out <= 26'h1d48054;
         146: out <= 26'h1e44053;
         147: out <= 26'h1f44055;
         148: out <= 26'h204c055;
         149: out <= 26'h213f851;
         150: out <= 26'h224b853;
         151: out <= 26'h2353855;
         152: out <= 26'h175f85e;
         153: out <= 26'h1a6b85f;
         154: out <= 26'h1d77860;
         155: out <= 26'h1e85062;
         156: out <= 26'h1f79063;
         157: out <= 26'h1f7c05d;
         158: out <= 26'h175d05e;
         159: out <= 26'h175c05d;
         160: out <= 26'h1a6905e;
         161: out <= 26'h1d6105b;
         162: out <= 26'h1e6505c;
         163: out <= 26'h2001056;
         164: out <= 26'h186005b;
         165: out <= 26'h196405c;
         166: out <= 26'h56;
         167: out <= 26'h1660059;
         168: out <= 26'h1b61040;
         169: out <= 26'h1c65058;
         170: out <= 26'h210105c;
         171: out <= 26'h2263858;
         172: out <= 26'h2367859;
         173: out <= 26'h2403840;
         174: out <= 26'h1963859;
         175: out <= 26'h1863840;
         176: out <= 26'h3856;
         177: out <= 26'h168b85b;
         178: out <= 26'h1b8f85c;
         179: out <= 26'h1c93861;
         180: out <= 26'h165805b;
         181: out <= 26'h165805c;
         182: out <= 26'h1b58041;
         183: out <= 26'h1c6e041;
         184: out <= 26'h1b6f85c;
         185: out <= 26'h1c6e081;
         186: out <= 26'h1b6f85c;
         187: out <= 26'h1c6e101;
         188: out <= 26'h1b6f85c;
         189: out <= 26'h1c6e201;
         190: out <= 26'h1b6f85c;
         191: out <= 26'h1c6e401;
         192: out <= 26'h1b6f85c;
         193: out <= 26'h1c6e801;
         194: out <= 26'h1c6f85c;
         195: out <= 26'h1c72801;
         196: out <= 26'h1b6f85c;
         197: out <= 26'h1b6e041;
         198: out <= 26'h166f856;
         199: out <= 26'h166f856;
         200: out <= 26'h1b8d064;
         201: out <= 26'h1c8905b;
         202: out <= 26'h71040;
         203: out <= 26'h1991059;
         204: out <= 26'h186d058;
         205: out <= 26'h5b840;
         206: out <= 26'h195b859;
         207: out <= 26'h165b858;
         208: out <= 26'h187405e;
         209: out <= 26'h1b74060;
         210: out <= 26'h1c78060;
         211: out <= 26'h2100059;
         212: out <= 26'h2200056;
         213: out <= 26'h2364056;
         214: out <= 26'h1d77840;
         215: out <= 26'h1e7b859;
         216: out <= 26'h2083856;
         217: out <= 26'h1863861;
         218: out <= 26'h1b6f862;
         219: out <= 26'h1c73863;
         220: out <= 26'h1d7505e;
         221: out <= 26'h1e75060;
         222: out <= 26'h1e7805c;
         223: out <= 26'h186105d;
         224: out <= 26'h186005c;
         225: out <= 26'h1b6d05d;
         226: out <= 26'h1c7c057;
         227: out <= 26'h1d7c05a;
         228: out <= 26'h205c05a;
         229: out <= 26'h2100059;
         230: out <= 26'h2200056;
         231: out <= 26'h2364056;
         232: out <= 26'h7f840;
         233: out <= 26'h175f859;
         234: out <= 26'h166b856;
         235: out <= 26'h1973861;
         236: out <= 26'h1a77862;
         237: out <= 26'h1c83863;
         238: out <= 26'h1057;
         239: out <= 26'h1601056;
         240: out <= 26'h165805c;
         241: out <= 26'h1765040;
         242: out <= 26'h175c05c;
         243: out <= 26'h69040;
         244: out <= 26'h1978056;
         245: out <= 26'h1a60057;
         246: out <= 26'h1c6d040;
         247: out <= 26'h1d7b85b;
         248: out <= 26'h1f5b840;
         249: out <= 26'h1b6385b;
         250: out <= 26'h5f840;
         251: out <= 26'h206785c;
         252: out <= 26'h165b858;
         253: out <= 26'h177b857;
         254: out <= 26'h186785a;
         255: out <= 26'h196b85c;
         256: out <= 26'h1a58057;
         257: out <= 26'h1869058;
         258: out <= 26'h1a6c040;
         259: out <= 26'h1a6805a;
         260: out <= 26'h105b;
         261: out <= 26'h1b7d05d;
         262: out <= 26'h1b6c060;
         263: out <= 26'h1c0805d;
         264: out <= 26'h1c7005f;
         265: out <= 26'h1c7005a;
         266: out <= 26'h1659057;
         267: out <= 26'h165805b;
         268: out <= 26'h1769058;
         269: out <= 26'h1d64040;
         270: out <= 26'h1b7505b;
         271: out <= 26'h1860058;
         272: out <= 26'h186105a;
         273: out <= 26'h64040;
         274: out <= 26'h1972041;
         275: out <= 26'h1a5a041;
         276: out <= 26'h1d5e041;
         277: out <= 26'h1e6e041;
         278: out <= 26'h1f62041;
         279: out <= 26'h2002041;
         280: out <= 26'h196405d;
         281: out <= 26'h196405f;
         282: out <= 26'h1a6805a;
         283: out <= 26'h1a6905e;
         284: out <= 26'h1a69060;
         285: out <= 26'h1d7505f;
         286: out <= 26'h1e8105e;
         287: out <= 26'h2080060;
         288: out <= 26'h1966041;
         289: out <= 26'h1a6a041;
         290: out <= 26'h1d76041;
         291: out <= 26'h1e7a041;
         292: out <= 26'h1f7e041;
         293: out <= 26'h2082041;
         294: out <= 26'h196405d;
         295: out <= 26'h196405f;
         296: out <= 26'h1a6805a;
         297: out <= 26'h1a6905e;
         298: out <= 26'h1a69060;
         299: out <= 26'h1d7505f;
         300: out <= 26'h1e8105e;
         301: out <= 26'h2080060;
         302: out <= 26'h2170056;
         303: out <= 26'h225c05b;
         304: out <= 26'h2361040;
         305: out <= 26'h2473858;
         306: out <= 26'h255b840;
         307: out <= 26'h185f858;
         308: out <= 26'h6f840;
         309: out <= 26'h2687863;
         310: out <= 26'h165b857;
         311: out <= 26'h177385b;
         312: out <= 26'h1b87862;
         313: out <= 26'h1c8b863;
         314: out <= 26'h2158057;
         315: out <= 26'h1b8505b;
         316: out <= 26'h2160040;
         317: out <= 26'h2184061;
         318: out <= 26'h1058;
         319: out <= 26'h1895064;
         320: out <= 26'h1860066;
         321: out <= 26'h2208064;
         322: out <= 26'h2288065;
         323: out <= 26'h2288061;
         324: out <= 26'h1659057;
         325: out <= 26'h1658058;
         326: out <= 26'h178505b;
         327: out <= 26'h2370040;
         328: out <= 26'h188d058;
         329: out <= 26'h1b6c05b;
         330: out <= 26'h1b6d061;
         331: out <= 26'h70040;
         332: out <= 26'h1a6805a;
         333: out <= 26'h1c7805e;
         334: out <= 26'h1e80060;
         335: out <= 26'h206405f;
         336: out <= 26'h218005d;
         337: out <= 26'h208105d;
         338: out <= 26'h238805b;
         339: out <= 26'h248c057;
         340: out <= 26'h238d057;
         341: out <= 26'h196505f;
         342: out <= 26'h256505c;
         343: out <= 26'h196405c;
         344: out <= 26'h228905b;
         345: out <= 26'h2689058;
         346: out <= 26'h2288058;
         347: out <= 26'h276805e;
         348: out <= 26'h289c05c;
         349: out <= 26'h1c9d05c;
         350: out <= 26'h2758040;
         351: out <= 26'h299c058;
         352: out <= 26'h189d058;
         353: out <= 26'h1a6905e;
         354: out <= 26'h276805d;
         355: out <= 26'h1a6905d;
         356: out <= 26'h1659040;
         357: out <= 26'h1d58057;
         358: out <= 26'h1659057;
         359: out <= 26'h1784068;
         360: out <= 26'h2a90069;
         361: out <= 26'h2b94067;
         362: out <= 26'h2c9805d;
         363: out <= 26'h2d8005c;
         364: out <= 26'h2e8c058;
         365: out <= 26'h2f6405a;
         366: out <= 26'h3088056;
         367: out <= 26'h317c05e;
         368: out <= 26'h326c040;
         369: out <= 26'h2187864;
         370: out <= 26'h175f86a;
         371: out <= 26'h24a3869;
         372: out <= 26'h2597866;
         373: out <= 26'h26af86c;
         374: out <= 26'h1d9f85d;
         375: out <= 26'h2083863;
         376: out <= 26'h23b786e;
         377: out <= 26'h1873858;
         378: out <= 26'h1967862;
         379: out <= 26'h1cbf870;
         380: out <= 26'h166b856;
         381: out <= 26'h1a7f85b;
         382: out <= 26'h1bc7872;
         383: out <= 26'h7b840;
         384: out <= 26'h1e84066;
         385: out <= 26'h1e7805a;
         386: out <= 26'h1f9005c;
         387: out <= 26'h1f7c040;
         388: out <= 26'h1a8005a;
         389: out <= 26'h60040;
         390: out <= 26'h40;
         391: out <= 26'h188c05b;
         392: out <= 26'h2000064;
         393: out <= 26'h2269061;
         394: out <= 26'h1064;
         395: out <= 26'h5d;
         396: out <= 26'h56;
         397: out <= 26'h1a68061;
         398: out <= 26'h1a69065;
         399: out <= 26'h1a69059;
         400: out <= 26'h97d05e;
         401: out <= 26'h925065;
         402: out <= 26'h924056;
         403: out <= 26'ha7805f;
         404: out <= 26'ha29057;
         405: out <= 26'ha2805d;
         406: out <= 26'ha28059;
         407: out <= 26'ha2905b;
         408: out <= 26'hb80062;
         409: out <= 26'hc81062;
         410: out <= 26'hc30058;
         411: out <= 26'hc31057;
         412: out <= 26'hd0005a;
         413: out <= 26'he0105a;
         414: out <= 26'he38058;
         415: out <= 26'he38057;
         416: out <= 26'he39066;
         417: out <= 26'he3905c;
         default: out <= 0;
      endcase
endmodule
