//File name=Module name=JTAG_SpW  2005-1-18      btltz@mail.china.com      btltz from CASIC,China 
//Description:   JTAG organization for SpaceWire node device ,  Approximate area:
//Origin:        SpaceWire Std - Draft-1 of ESTEC,ESA
//--     TODO:
////////////////////////////////////////////////////////////////////////////////////

/*synthesis translate_off*/
`include "timescale.v"
/*synthesis translate_on */
module JTAG_SpW #()
               ( output TDO,
                 input TDI,
		   input TCK
                );


endmodule

