import RegFile::*;

