-- AHB2HPI enable 
  constant CFG_AHB2HPI  : integer := CONFIG_AHB2HPI_ENABLE;

