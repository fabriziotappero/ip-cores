----==============================================================----
----                                                              ----
---- Filename: hw_loops5_top_tb.vhd                               ----
---- Module description: Simple testbench for the "hw_loops5_top" ----
----                     top-level module                         ----
----                                                              ----
---- Author: Nikolaos Kavvadias                                   ----
----         nkavv@skiathos.physics.auth.gr                       ----
----                                                              ---- 
----                                                              ----
---- Downloaded from: http://wwww.opencores.org/cores/hwlu        ----
----                                                              ----
---- To Do:                                                       ----
----         1. Should be improved. A more thorough testbench is  ----
----            needed.                                           ----
----         2. The testbench file for the top-level module will  ----
----            be generated by corresponding C tool.             ----
----                                                              ----
---- Author: Nikolaos Kavvadias                                   ----
----         nkavv@skiathos.physics.auth.gr                       ----
----                                                              ----
----==============================================================----
----                                                              ----
---- Copyright (C) 2004 Nikolaos Kavvadias                        ----
----                    nick-kavi.8m.com                          ----
----                    nkavv@skiathos.physics.auth.gr            ----
----                    nick_ka_vi@hotmail.com                    ----
----                                                              ----
---- This source file may be used and distributed without         ----
---- restriction provided that this copyright statement is not    ----
---- removed from the file and that any derivative work contains  ----
---- the original copyright notice and the associated disclaimer. ----
----                                                              ----
---- This source file is free software; you can redistribute it   ----
---- and/or modify it under the terms of the GNU Lesser General   ----
---- Public License as published by the Free Software Foundation; ----
---- either version 2.1 of the License, or (at your option) any   ----
---- later version.                                               ----
----                                                              ----
---- This source is distributed in the hope that it will be       ----
---- useful, but WITHOUT ANY WARRANTY; without even the implied   ----
---- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ----
---- PURPOSE. See the GNU Lesser General Public License for more  ----
---- details.                                                     ----
----                                                              ----
---- You should have received a copy of the GNU Lesser General    ----
---- Public License along with this source; if not, download it   ----
---- from <http://www.opencores.org/lgpl.shtml>                   ----
----                                                              ----
----==============================================================----
--
-- CVS Revision History
--    

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_textio.all;
use STD.textio.all;


entity hwloop_top_tb is
  generic (	
    DW  : integer := 8;
    NLP : integer := 5    
  );
end hwloop_top_tb;
                              
                              
architecture tb_architecture of hwloop_top_tb is
--
-- Component declaration of the DUT
component hw_looping is
  generic (
    DW : integer := 8;
    NLP : integer := 5
  );
  port (                 
    clk            : in std_logic;
    reset          : in std_logic;
	task_loop5_end : in std_logic;
    loop1_count    : in std_logic_vector(DW-1 downto 0);
    loop2_count    : in std_logic_vector(DW-1 downto 0);
    loop3_count    : in std_logic_vector(DW-1 downto 0);
    loop4_count    : in std_logic_vector(DW-1 downto 0);
    loop5_count    : in std_logic_vector(DW-1 downto 0);
    index1         : out std_logic_vector(DW-1 downto 0);
    index2         : out std_logic_vector(DW-1 downto 0);
    index3         : out std_logic_vector(DW-1 downto 0);
    index4         : out std_logic_vector(DW-1 downto 0);
    index5         : out std_logic_vector(DW-1 downto 0);   
    loops_end      : out std_logic
  );
end component;
-- 
-- Signal declarations
-- Stimulus signals - signals mapped to the I/IO ports of tested entity
signal clk            : std_logic;
signal reset          : std_logic;
signal task_loop5_end : std_logic;
signal loop1_count    : std_logic_vector(DW-1 downto 0);    
signal loop2_count    : std_logic_vector(DW-1 downto 0);    
signal loop3_count    : std_logic_vector(DW-1 downto 0);    
signal loop4_count    : std_logic_vector(DW-1 downto 0);    
signal loop5_count    : std_logic_vector(DW-1 downto 0);    
-- Signals mapped to the output ports of tested entity
signal index1         : std_logic_vector(DW-1 downto 0);    
signal index2         : std_logic_vector(DW-1 downto 0);    
signal index3         : std_logic_vector(DW-1 downto 0);    
signal index4         : std_logic_vector(DW-1 downto 0);    
signal index5         : std_logic_vector(DW-1 downto 0);    
signal loops_end      : std_logic;                     
--
-- Constant declarations
constant CLK_PERIOD : time := 10 ns;

begin

  -- Unit Under Test port map
  UUT : hw_looping
    generic map (    
      DW => DW,
      NLP => NLP
    )
    port map (
      clk => clk,
      reset => reset,
	  task_loop5_end => task_loop5_end,
      loop1_count => loop1_count,
      loop2_count => loop2_count,
      loop3_count => loop3_count,
      loop4_count => loop4_count,
      loop5_count => loop5_count,
      index1 => index1,
      index2 => index2,
      index3 => index3,
      index4 => index4,
      index5 => index5,
	  loops_end => loops_end
    );
    
CLK_GEN_PROC: process(clk)
begin
  if (clk = 'U') then 
    clk <= '1'; 
  else 
    clk <= not clk after CLK_PERIOD/2; 
  end if;
end process CLK_GEN_PROC;	

DATA_STIM: process
begin
  reset <= '0';
  task_loop5_end <= '0';
  loop1_count <= X"00";
  loop2_count <= X"00";
  loop3_count <= X"00";
  loop4_count <= X"00";
  loop5_count <= X"00";
  wait for CLK_PERIOD;
  --
  reset <= '1';
  task_loop5_end <= '0';
  loop1_count <= X"00";
  loop2_count <= X"00";
  loop3_count <= X"00";
  loop4_count <= X"00";
  loop5_count <= X"00";
  wait for CLK_PERIOD;
  --
  reset <= '0';		   
  task_loop5_end <= '1';
  loop1_count <= X"04";
  loop2_count <= X"06";
  loop3_count <= X"02";
  loop4_count <= X"04";
  loop5_count <= X"03";
  wait for CLK_PERIOD;
  --
  -- Apply same inputs (written in some kind of 
  -- configuration memory) for large amount of time, 
  -- e.g. 1000 clock periods
  wait for 1000*CLK_PERIOD;
  --            
end process DATA_STIM;

end tb_architecture;


configuration TESTBENCH_FOR_hw_looping of hwloop_top_tb is
	for tb_architecture
		for UUT : hw_looping
			use entity work.hw_looping(structural);
		end for;
	end for;
end TESTBENCH_FOR_hw_looping;
