-------------------------------------------------------------------------------
--
-- The skip unit.
-- Skip conditions are checked here and communicated to the decoder unit.
--
-- $Id: t400_skip-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_skip_rtl_c0 of t400_skip is

  for rtl
  end for;

end t400_skip_rtl_c0;
