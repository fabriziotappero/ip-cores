library verilog;
use verilog.vl_types.all;
entity mobile_sdr is
    generic(
        tCK             : integer := 6000;
        tCK3_min        : integer := 6000;
        tCK2_min        : integer := 9600;
        tCK1_min        : integer := 0;
        tAC3            : integer := 5000;
        tAC2            : integer := 8000;
        tAC1            : integer := 0;
        tHZ3            : integer := 5000;
        tHZ2            : integer := 8000;
        tHZ1            : integer := 0;
        tOH             : integer := 2500;
        tMRD            : integer := 2;
        tRAS            : integer := 42000;
        tRC             : integer := 60000;
        tRFC            : integer := 97500;
        tRCD            : integer := 18000;
        tRP             : integer := 18000;
        tRRD            : integer := 2;
        tWRa            : integer := 7500;
        tWRm            : integer := 15000;
        tCH             : integer := 2600;
        tCL             : integer := 2600;
        tXSR            : integer := 120000;
        ADDR_BITS       : integer := 13;
        ROW_BITS        : integer := 13;
        DQ_BITS         : integer := 16;
        DM_BITS         : integer := 2;
        COL_BITS        : integer := 10;
        BA_BITS         : integer := 2;
        part_mem_bits   : integer := 10;
        part_size       : integer := 256;
        NOP             : integer := 39;
        ACTIVATE        : integer := 35;
        READ            : integer := 37;
        READ_AP         : integer := 53;
        READ_SUSPEND    : integer := 5;
        READ_AP_SUSPEND : integer := 21;
        WRITE           : integer := 36;
        WRITE_AP        : integer := 52;
        WRITE_SUSPEND   : integer := 4;
        WRITE_AP_SUSPEND: integer := 20;
        BURST_TERMINATE : integer := 38;
        POWER_DOWN_CI   : integer := 15;
        POWER_DOWN_NOP  : integer := 7;
        DEEP_POWER_DOWN : integer := 6;
        PRECHARGE       : integer := 34;
        PRECHARGE_ALL   : integer := 50;
        AUTO_REFRESH    : integer := 33;
        SELF_REFRESH    : integer := 1;
        LOAD_MODE       : integer := 32;
        CKE_DISABLE     : integer := 31;
        DEBUG           : integer := 1;
        ERR_MAX_REPORTED: integer := -1;
        ERR_MAX         : integer := -1;
        MSGLENGTH       : integer := 256;
        ERR_CODES       : integer := 16;
        ERR_MISC        : integer := 1;
        ERR_CMD         : integer := 2;
        ERR_STATUS      : integer := 3;
        ERR_tMRD        : integer := 4;
        ERR_tRAS        : integer := 5;
        ERR_tRC         : integer := 6;
        ERR_tRFC        : integer := 7;
        ERR_tRCD        : integer := 8;
        ERR_tRP         : integer := 9;
        ERR_tRRD        : integer := 11;
        ERR_tWR         : integer := 12;
        ERR_tCH         : integer := 13;
        ERR_tCL         : integer := 14;
        ERR_tXSR        : integer := 15;
        ERR_tCK_MIN     : integer := 16
    );
    port(
        clk             : in     vl_logic;
        cke             : in     vl_logic;
        addr            : in     vl_logic_vector;
        ba              : in     vl_logic_vector;
        cs_n            : in     vl_logic;
        ras_n           : in     vl_logic;
        cas_n           : in     vl_logic;
        we_n            : in     vl_logic;
        dq              : inout  vl_logic_vector;
        dqm             : in     vl_logic_vector
    );
end mobile_sdr;
