-- PS/2 interface
  constant CFG_PS2_ENABLE  : integer := CONFIG_PS2_ENABLE;

