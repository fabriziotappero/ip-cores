-- ------------------------------------------------------------------------
-- Copyright (C) 2005 Arif Endro Nugroho
-- All rights reserved.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY ARIF ENDRO NUGROHO "AS IS" AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL ARIF ENDRO NUGROHO BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
-- ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
-- 
-- End Of License.
-- ------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity input is
   port (
      clock   : in  bit;
      clear   : in  bit;
      start   : out bit;
      rom_pos : out integer;
      rxin    : out bit_vector (07 downto 00)
      );
end input;

architecture test_bench of input is

type rom_bank is array ( 00000 to 19999 ) of bit_vector (7 downto 0);

constant input_bank : rom_bank :=
(

 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000"

);

signal input_counter : integer range 0 to 19999 := 0;
signal start_fifo    : bit_vector (7 downto 0) := ( B"0100_0000" );
signal clk : bit;

begin

process (clk, clear)
begin
if (clear = '1') then
    rxin <= (others => '0');
elsif (clk = '1' and clk'event) then
    rxin <= input_bank(input_counter);
end if;
end process;

process (clk, clear)
begin
if (clear = '1') then
    input_counter <= 0;
elsif (clk = '1' and clk'event) then
    if (input_counter < 19999) then
    input_counter <= input_counter + 1;
    else
    input_counter <= 0;
    end if;
end if;
end process;

rom_pos <= input_counter;

process (clk, clear)
begin
if (clear = '1') then
    start_fifo <= B"0100_0000";
elsif ( clk = '1' and clk'event) then
    start_fifo <= start_fifo (6 downto 0) & start_fifo (7);
end if;
end process;

clk   <= clock;
start <= start_fifo (7);

end test_bench;
