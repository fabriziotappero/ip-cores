-- -------------------------------------------------------------------------
-- -------------------------------------------------------------------------
--
-- Revision Control Information
--
-- $RCSfile: timing_adapter_32.vhd,v $
-- $Source: /ipbu/cvs/sio/projects/TriSpeedEthernet/src/testbench/models/vhdl/ethernet_model/gen/timing_adapter_32.vhd,v $
--
-- $Revision: #1 $
-- $Date: 2008/08/09 $
-- Check in by : $Author: sc-build $
-- Author      : SKNg/TTChong
--
-- Project     : Triple Speed Ethernet - 10/100/1000 MAC
--
-- Description : (Simulation only)
--
-- Timing adapater  (from 3 to zero ready latency) Client Interface Ethernet Traffic Generator
-- Instantiating a FIFO unit 
-- 
-- ALTERA Confidential and Proprietary
-- Copyright 2006 (c) Altera Corporation
-- All rights reserved
--
-- -------------------------------------------------------------------------
-- -------------------------------------------------------------------------

-- --------------------------------------------------------------------------------
--| Avalon Streaming Timing Adapter
-- --------------------------------------------------------------------------------

--IP Functional Simulation Model
--VERSION_BEGIN 7.1SP1 cbx_mgl 2007:06:11:16:05:04:SJ cbx_simgen 2007:03:19:18:39:32:SJ  VERSION_END


-- Legal Notice: � 2003 Altera Corporation. All rights reserved.
-- You may only use these  simulation  model  output files for simulation
-- purposes and expressly not for synthesis or any other purposes (in which
-- event  Altera disclaims all warranties of any kind). Your use of  Altera
-- Corporation's design tools, logic functions and other software and tools,
-- and its AMPP partner logic functions, and any output files any of the
-- foregoing (including device programming or simulation files), and any
-- associated documentation or information  are expressly subject to the
-- terms and conditions of the  Altera Program License Subscription Agreement
-- or other applicable license agreement, including, without limitation, that
-- your use is for the sole purpose of programming logic devices manufactured
-- by Altera and sold by Altera or its authorized distributors.  Please refer
-- to the applicable agreement for further details.


--synopsys translate_off

 LIBRARY altera_mf;
 USE altera_mf.altera_mf_components.all;

 LIBRARY sgate;
 USE sgate.sgate_pack.all;

--synthesis_resources = altsyncram 1 lut 9 mux21 15 oper_add 3 oper_less_than 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;


 
 ENTITY  timing_adapter_32 IS 
     PORT 
     ( 
         -- Interface: clk
         clk                :   IN      STD_LOGIC;
         reset              :   IN      STD_LOGIC;

         -- Interface: in
         in_ready           :   OUT     STD_LOGIC;
         in_valid           :   IN      STD_LOGIC;
         in_data            :   IN      STD_LOGIC_VECTOR (31 DOWNTO 0);
         in_startofpacket   :   IN      STD_LOGIC;
         in_endofpacket     :   IN      STD_LOGIC;
         in_empty           :   IN      STD_LOGIC_VECTOR (1 DOWNTO 0);
         in_error           :   IN      STD_LOGIC;
         -- Interface: out
         out_ready          :   IN      STD_LOGIC;
         out_valid          :   OUT     STD_LOGIC;
         out_data           :   OUT     STD_LOGIC_VECTOR (31 DOWNTO 0);
         out_startofpacket  :   OUT     STD_LOGIC;
         out_endofpacket    :   OUT     STD_LOGIC;
         out_empty          :   OUT     STD_LOGIC_VECTOR (1 DOWNTO 0);
         out_error          :   OUT     STD_LOGIC
     ); 
 END timing_adapter_32;

 ARCHITECTURE RTL OF timing_adapter_32 IS


	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_204q	:	STD_LOGIC := '0';
	 SIGNAL  wire_ni_w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_100_580q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_101_582q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_102_584q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_103_586q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_104_588q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_105_590q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_106_592q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_107_594q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_108_596q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_109_598q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_10_400q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_110_600q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_111_602q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_112_604q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_113_606q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_114_608q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_115_610q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_116_612q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_117_614q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_118_616q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_119_618q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_11_402q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_120_620q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_121_622q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_122_624q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_123_626q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_124_628q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_125_630q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_126_632q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_127_634q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_128_636q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_129_638q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_12_404q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_130_640q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_131_642q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_132_644q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_133_646q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_134_648q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_135_650q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_136_652q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_137_654q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_138_656q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_139_658q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_13_406q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_140_660q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_141_662q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_142_664q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_143_666q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_144_668q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_145_670q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_146_672q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_147_674q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_148_676q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_149_678q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_14_408q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_150_680q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_151_682q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_152_684q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_153_686q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_154_688q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_155_690q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_156_692q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_157_694q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_158_696q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_159_698q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_15_410q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_160_700q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_161_702q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_162_704q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_163_706q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_164_708q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_165_710q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_166_712q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_167_714q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_168_716q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_169_718q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_16_412q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_170_720q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_171_722q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_172_724q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_173_726q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_174_728q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_175_730q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_176_732q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_177_734q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_178_736q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_179_738q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_17_414q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_180_740q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_181_742q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_182_744q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_183_746q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_184_748q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_185_750q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_186_752q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_187_754q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_188_756q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_189_758q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_18_416q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_190_760q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_191_762q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_192_764q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_193_766q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_194_768q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_195_770q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_196_772q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_197_774q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_198_776q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_199_778q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_19_418q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_1_382q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_200_780q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_201_782q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_202_784q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_203_786q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_204_788q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_205_790q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_206_792q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_207_794q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_208_796q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_209_798q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_20_420q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_210_800q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_211_802q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_212_804q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_213_806q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_214_808q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_215_810q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_216_812q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_217_814q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_218_816q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_219_818q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_21_422q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_220_820q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_221_822q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_222_824q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_223_826q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_224_828q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_225_830q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_226_832q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_227_834q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_228_836q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_229_838q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_22_424q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_230_840q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_231_842q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_232_844q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_233_846q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_234_848q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_235_850q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_236_852q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_237_854q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_238_856q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_239_858q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_23_426q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_240_860q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_241_862q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_242_864q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_243_866q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_244_868q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_245_870q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_246_872q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_247_874q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_248_876q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_249_878q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_24_428q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_250_880q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_251_882q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_252_884q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_253_886q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_254_888q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_255_890q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_256_892q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_257_894q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_258_896q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_259_898q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_25_430q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_260_900q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_261_902q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_262_904q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_263_906q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_264_908q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_265_910q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_266_912q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_267_914q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_268_916q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_269_918q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_26_432q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_270_920q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_271_922q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_272_924q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_273_926q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_274_928q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_275_930q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_276_932q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_277_934q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_278_936q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_279_938q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_27_434q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_280_940q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_281_942q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_282_944q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_283_946q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_284_948q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_285_950q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_286_952q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_287_954q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_288_956q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_289_958q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_28_436q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_290_960q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_291_962q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_292_964q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_293_966q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_294_968q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_295_970q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_296_972q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_29_438q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_2_384q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_30_440q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_31_442q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_32_444q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_33_446q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_34_448q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_35_450q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_36_452q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_37_454q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_38_456q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_39_458q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_3_386q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_40_460q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_41_462q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_42_464q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_43_466q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_44_468q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_45_470q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_46_472q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_47_474q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_48_476q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_49_478q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_4_388q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_50_480q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_51_482q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_52_484q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_53_486q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_54_488q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_55_490q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_56_492q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_57_494q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_58_496q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_59_498q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_5_390q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_60_500q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_61_502q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_62_504q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_63_506q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_64_508q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_65_510q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_66_512q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_67_514q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_68_516q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_69_518q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_6_392q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_70_520q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_71_522q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_72_524q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_73_526q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_74_528q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_75_530q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_76_532q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_77_534q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_78_536q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_79_538q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_7_394q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_80_540q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_81_542q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_82_544q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_83_546q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_84_548q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_85_550q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_86_552q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_87_554q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_88_556q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_89_558q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_8_396q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_90_560q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_91_562q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_92_564q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_93_566q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_94_568q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_95_570q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_96_572q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_97_574q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_98_576q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_99_578q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_9_398q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_187q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q	:	STD_LOGIC := '0';
	 SIGNAL	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q	:	STD_LOGIC := '0';
	 SIGNAL  wire_nO_w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_nO_w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_nO_w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_nO_w84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_100_567m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_101_569m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_102_571m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_103_573m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_104_575m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_105_577m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_106_579m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_107_581m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_108_583m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_109_585m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_10_387m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_110_587m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_111_589m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_112_591m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_113_593m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_114_595m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_115_597m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_116_599m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_117_601m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_118_603m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_119_605m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_11_389m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_120_607m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_121_609m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_122_611m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_123_613m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_124_615m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_125_617m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_126_619m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_127_621m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_128_623m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_129_625m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_12_391m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_130_627m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_131_629m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_132_631m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_133_633m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_134_635m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_135_637m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_136_639m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_137_641m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_138_643m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_139_645m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_13_393m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_140_647m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_141_649m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_142_651m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_143_653m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_144_655m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_145_657m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_146_659m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_147_661m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_148_663m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_149_665m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_14_395m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_150_667m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_151_669m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_152_671m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_153_673m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_154_675m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_155_677m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_156_679m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_157_681m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_158_683m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_159_685m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_15_397m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_160_687m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_161_689m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_162_691m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_163_693m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_164_695m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_165_697m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_166_699m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_167_701m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_168_703m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_169_705m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_16_399m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_170_707m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_171_709m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_172_711m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_173_713m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_174_715m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_175_717m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_176_719m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_177_721m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_178_723m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_179_725m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_17_401m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_180_727m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_181_729m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_182_731m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_183_733m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_184_735m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_185_737m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_186_739m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_187_741m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_188_743m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_189_745m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_18_403m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_190_747m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_191_749m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_192_751m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_193_753m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_194_755m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_195_757m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_196_759m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_197_761m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_198_763m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_199_765m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_19_405m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_200_767m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_201_769m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_202_771m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_203_773m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_204_775m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_205_777m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_206_779m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_207_781m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_208_783m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_209_785m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_20_407m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_210_787m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_211_789m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_212_791m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_213_793m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_214_795m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_215_797m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_216_799m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_217_801m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_218_803m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_219_805m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_21_409m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_220_807m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_221_809m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_222_811m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_223_813m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_224_815m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_225_817m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_226_819m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_227_821m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_228_823m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_229_825m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_22_411m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_230_827m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_231_829m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_232_831m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_233_833m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_234_835m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_235_837m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_236_839m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_237_841m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_238_843m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_239_845m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_23_413m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_240_847m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_241_849m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_242_851m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_243_853m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_244_855m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_245_857m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_246_859m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_247_861m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_248_863m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_249_865m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_24_415m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_250_867m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_251_869m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_252_871m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_253_873m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_254_875m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_255_877m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_256_879m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_257_881m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_258_883m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_259_885m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_25_417m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_260_887m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_261_889m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_262_891m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_263_893m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_264_895m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_265_897m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_266_899m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_267_901m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_268_903m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_269_905m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_26_419m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_270_907m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_271_909m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_272_911m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_273_913m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_274_915m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_275_917m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_276_919m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_277_921m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_278_923m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_279_925m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_27_421m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_280_927m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_281_929m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_282_931m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_283_933m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_284_935m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_285_937m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_286_939m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_287_941m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_288_943m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_289_945m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_28_423m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_290_947m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_291_949m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_292_951m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_293_953m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_294_955m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_295_957m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_296_959m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_297_961m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_298_963m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_299_965m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_29_425m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_300_967m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_301_969m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_302_971m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_303_973m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_30_427m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_31_429m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_32_431m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_33_433m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_34_435m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_35_437m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_36_439m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_37_441m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_38_443m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_39_445m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_40_447m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_41_449m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_42_451m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_43_453m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_44_455m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_45_457m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_46_459m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_47_461m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_48_463m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_49_465m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_50_467m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_51_469m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_52_471m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_53_473m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_54_475m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_55_477m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_56_479m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_57_481m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_58_483m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_59_485m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_60_487m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_61_489m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_62_491m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_63_493m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_64_495m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_65_497m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_66_499m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_67_501m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_68_503m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_69_505m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_70_507m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_71_509m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_72_511m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_73_513m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_74_515m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_75_517m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_76_519m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_77_521m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_78_523m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_79_525m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_80_527m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_81_529m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_82_531m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_83_533m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_84_535m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_85_537m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_86_539m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_87_541m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_88_543m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_89_545m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_8_383m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_90_547m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_91_549m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_92_551m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_93_553m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_94_555m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_95_557m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_96_559m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_97_561m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_98_563m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_99_565m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_9_385m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_0_184m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_1_189m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_2_192m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_0_176m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_1_175m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_2_174m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_0_180m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_1_185m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_2_191m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_4_334m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_0_190m_dataout	:	STD_LOGIC;
	 SIGNAL	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_1_193m_dataout	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_a	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_b	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_a	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_b	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_a	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_b	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_o	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_i	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_lessthan0_2_a	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_lessthan0_2_b	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_lessthan0_2_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_o	:	STD_LOGIC;
	 SIGNAL  wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_sel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_3_195_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_3_981_dataout :	STD_LOGIC;
	 SIGNAL  s_wire_vcc :	STD_LOGIC;
 BEGIN

	wire_gnd <= '0';
	wire_w_lg_reset102w(0) <= NOT reset;
	wire_w106w(0) <= NOT s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_3_195_dataout;
	in_ready <= wire_timing_adapter_32_lessthan0_2_o;
	out_data <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_o
 & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_o);
	out_empty <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_o & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_o);
	out_endofpacket <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_o;
	out_error <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_o;
	out_startofpacket <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_o;
	out_valid <= timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_187q;
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(0));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(1));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(2));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(3));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(4));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(5));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(6));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout <= (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout AND wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o(7));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout <= (wire_nO_w88w(0) AND in_valid);
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout <= (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_187q AND out_ready);
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_3_195_dataout <= (in_valid AND (wire_nO_w88w(0) AND s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout));
	s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_3_981_dataout <= (((NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(0))) AND (NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(1)))) AND (NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(2))));
	s_wire_vcc <= '1';
	PROCESS (clk, reset)
	BEGIN
		IF (reset = '1') THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_204q <= '1';
		ELSIF (clk = '1' AND clk'event) THEN
			IF (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_3_195_dataout = '0') THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_204q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_2_192m_dataout;
			END IF;
		END IF;
	END PROCESS;
	wire_ni_w103w(0) <= NOT timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_204q;
	PROCESS (clk, reset)
	BEGIN
		IF (reset = '1') THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q <= '0';
		ELSIF (clk = '1' AND clk'event) THEN
			IF (s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout = '1') THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(0);
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(1);
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clk, reset)
	BEGIN
		IF (reset = '1') THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_100_580q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_101_582q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_102_584q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_103_586q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_104_588q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_105_590q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_106_592q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_107_594q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_108_596q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_109_598q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_10_400q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_110_600q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_111_602q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_112_604q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_113_606q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_114_608q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_115_610q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_116_612q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_117_614q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_118_616q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_119_618q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_11_402q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_120_620q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_121_622q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_122_624q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_123_626q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_124_628q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_125_630q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_126_632q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_127_634q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_128_636q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_129_638q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_12_404q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_130_640q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_131_642q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_132_644q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_133_646q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_134_648q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_135_650q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_136_652q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_137_654q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_138_656q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_139_658q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_13_406q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_140_660q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_141_662q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_142_664q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_143_666q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_144_668q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_145_670q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_146_672q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_147_674q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_148_676q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_149_678q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_14_408q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_150_680q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_151_682q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_152_684q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_153_686q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_154_688q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_155_690q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_156_692q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_157_694q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_158_696q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_159_698q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_15_410q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_160_700q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_161_702q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_162_704q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_163_706q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_164_708q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_165_710q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_166_712q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_167_714q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_168_716q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_169_718q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_16_412q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_170_720q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_171_722q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_172_724q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_173_726q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_174_728q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_175_730q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_176_732q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_177_734q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_178_736q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_179_738q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_17_414q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_180_740q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_181_742q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_182_744q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_183_746q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_184_748q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_185_750q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_186_752q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_187_754q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_188_756q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_189_758q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_18_416q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_190_760q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_191_762q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_192_764q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_193_766q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_194_768q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_195_770q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_196_772q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_197_774q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_198_776q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_199_778q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_19_418q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_1_382q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_200_780q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_201_782q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_202_784q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_203_786q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_204_788q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_205_790q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_206_792q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_207_794q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_208_796q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_209_798q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_20_420q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_210_800q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_211_802q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_212_804q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_213_806q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_214_808q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_215_810q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_216_812q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_217_814q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_218_816q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_219_818q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_21_422q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_220_820q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_221_822q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_222_824q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_223_826q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_224_828q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_225_830q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_226_832q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_227_834q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_228_836q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_229_838q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_22_424q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_230_840q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_231_842q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_232_844q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_233_846q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_234_848q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_235_850q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_236_852q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_237_854q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_238_856q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_239_858q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_23_426q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_240_860q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_241_862q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_242_864q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_243_866q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_244_868q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_245_870q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_246_872q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_247_874q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_248_876q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_249_878q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_24_428q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_250_880q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_251_882q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_252_884q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_253_886q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_254_888q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_255_890q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_256_892q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_257_894q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_258_896q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_259_898q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_25_430q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_260_900q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_261_902q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_262_904q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_263_906q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_264_908q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_265_910q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_266_912q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_267_914q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_268_916q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_269_918q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_26_432q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_270_920q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_271_922q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_272_924q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_273_926q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_274_928q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_275_930q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_276_932q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_277_934q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_278_936q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_279_938q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_27_434q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_280_940q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_281_942q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_282_944q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_283_946q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_284_948q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_285_950q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_286_952q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_287_954q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_288_956q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_289_958q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_28_436q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_290_960q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_291_962q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_292_964q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_293_966q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_294_968q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_295_970q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_296_972q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_29_438q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_2_384q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_30_440q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_31_442q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_32_444q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_33_446q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_34_448q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_35_450q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_36_452q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_37_454q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_38_456q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_39_458q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_3_386q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_40_460q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_41_462q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_42_464q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_43_466q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_44_468q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_45_470q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_46_472q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_47_474q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_48_476q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_49_478q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_4_388q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_50_480q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_51_482q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_52_484q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_53_486q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_54_488q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_55_490q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_56_492q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_57_494q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_58_496q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_59_498q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_5_390q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_60_500q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_61_502q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_62_504q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_63_506q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_64_508q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_65_510q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_66_512q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_67_514q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_68_516q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_69_518q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_6_392q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_70_520q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_71_522q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_72_524q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_73_526q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_74_528q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_75_530q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_76_532q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_77_534q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_78_536q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_79_538q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_7_394q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_80_540q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_81_542q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_82_544q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_83_546q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_84_548q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_85_550q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_86_552q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_87_554q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_88_556q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_89_558q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_8_396q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_90_560q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_91_562q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_92_564q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_93_566q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_94_568q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_95_570q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_96_572q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_97_574q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_98_576q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_99_578q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_9_398q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_187q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q <= '0';
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q <= '0';
		ELSIF (clk = '1' AND clk'event) THEN
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_4_334m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_100_580q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_107_581m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_101_582q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_108_583m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_102_584q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_109_585m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_103_586q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_110_587m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_104_588q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_111_589m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_105_590q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_112_591m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_106_592q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_113_593m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_107_594q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_114_595m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_108_596q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_115_597m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_109_598q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_116_599m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_10_400q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_17_401m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_110_600q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_117_601m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_111_602q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_118_603m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_112_604q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_119_605m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_113_606q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_120_607m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_114_608q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_121_609m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_115_610q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_122_611m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_116_612q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_123_613m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_117_614q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_124_615m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_118_616q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_125_617m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_119_618q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_126_619m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_11_402q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_18_403m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_120_620q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_127_621m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_121_622q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_128_623m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_122_624q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_129_625m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_123_626q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_130_627m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_124_628q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_131_629m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_125_630q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_132_631m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_126_632q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_133_633m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_127_634q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_134_635m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_128_636q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_135_637m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_129_638q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_136_639m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_12_404q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_19_405m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_130_640q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_137_641m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_131_642q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_138_643m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_132_644q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_139_645m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_133_646q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_140_647m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_134_648q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_141_649m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_135_650q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_142_651m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_136_652q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_143_653m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_137_654q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_144_655m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_138_656q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_145_657m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_139_658q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_146_659m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_13_406q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_20_407m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_140_660q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_147_661m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_141_662q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_148_663m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_142_664q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_149_665m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_143_666q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_150_667m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_144_668q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_151_669m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_145_670q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_152_671m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_146_672q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_153_673m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_147_674q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_154_675m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_148_676q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_155_677m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_149_678q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_156_679m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_14_408q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_21_409m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_150_680q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_157_681m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_151_682q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_158_683m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_152_684q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_159_685m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_153_686q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_160_687m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_154_688q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_161_689m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_155_690q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_162_691m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_156_692q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_163_693m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_157_694q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_164_695m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_158_696q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_165_697m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_159_698q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_166_699m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_15_410q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_22_411m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_160_700q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_167_701m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_161_702q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_168_703m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_162_704q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_169_705m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_163_706q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_170_707m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_164_708q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_171_709m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_165_710q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_172_711m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_166_712q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_173_713m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_167_714q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_174_715m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_168_716q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_175_717m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_169_718q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_176_719m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_16_412q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_23_413m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_170_720q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_177_721m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_171_722q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_178_723m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_172_724q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_179_725m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_173_726q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_180_727m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_174_728q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_181_729m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_175_730q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_182_731m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_176_732q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_183_733m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_177_734q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_184_735m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_178_736q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_185_737m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_179_738q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_186_739m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_17_414q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_24_415m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_180_740q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_187_741m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_181_742q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_188_743m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_182_744q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_189_745m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_183_746q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_190_747m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_184_748q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_191_749m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_185_750q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_192_751m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_186_752q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_193_753m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_187_754q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_194_755m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_188_756q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_195_757m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_189_758q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_196_759m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_18_416q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_25_417m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_190_760q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_197_761m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_191_762q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_198_763m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_192_764q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_199_765m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_193_766q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_200_767m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_194_768q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_201_769m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_195_770q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_202_771m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_196_772q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_203_773m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_197_774q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_204_775m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_198_776q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_205_777m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_199_778q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_206_779m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_19_418q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_26_419m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_1_382q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_8_383m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_200_780q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_207_781m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_201_782q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_208_783m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_202_784q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_209_785m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_203_786q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_210_787m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_204_788q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_211_789m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_205_790q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_212_791m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_206_792q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_213_793m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_207_794q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_214_795m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_208_796q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_215_797m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_209_798q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_216_799m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_20_420q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_27_421m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_210_800q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_217_801m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_211_802q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_218_803m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_212_804q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_219_805m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_213_806q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_220_807m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_214_808q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_221_809m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_215_810q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_222_811m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_216_812q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_223_813m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_217_814q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_224_815m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_218_816q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_225_817m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_219_818q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_226_819m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_21_422q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_28_423m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_220_820q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_227_821m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_221_822q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_228_823m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_222_824q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_229_825m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_223_826q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_230_827m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_224_828q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_231_829m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_225_830q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_232_831m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_226_832q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_233_833m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_227_834q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_234_835m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_228_836q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_235_837m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_229_838q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_236_839m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_22_424q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_29_425m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_230_840q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_237_841m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_231_842q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_238_843m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_232_844q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_239_845m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_233_846q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_240_847m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_234_848q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_241_849m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_235_850q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_242_851m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_236_852q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_243_853m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_237_854q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_244_855m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_238_856q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_245_857m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_239_858q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_246_859m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_23_426q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_30_427m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_240_860q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_247_861m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_241_862q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_248_863m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_242_864q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_249_865m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_243_866q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_250_867m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_244_868q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_251_869m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_245_870q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_252_871m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_246_872q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_253_873m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_247_874q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_254_875m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_248_876q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_255_877m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_249_878q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_256_879m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_24_428q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_31_429m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_250_880q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_257_881m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_251_882q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_258_883m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_252_884q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_259_885m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_253_886q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_260_887m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_254_888q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_261_889m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_255_890q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_262_891m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_256_892q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_263_893m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_257_894q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_264_895m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_258_896q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_265_897m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_259_898q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_266_899m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_25_430q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_32_431m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_260_900q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_267_901m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_261_902q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_268_903m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_262_904q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_269_905m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_263_906q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_270_907m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_264_908q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_271_909m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_265_910q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_272_911m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_266_912q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_273_913m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_267_914q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_274_915m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_268_916q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_275_917m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_269_918q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_276_919m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_26_432q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_33_433m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_270_920q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_277_921m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_271_922q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_278_923m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_272_924q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_279_925m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_273_926q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_280_927m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_274_928q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_281_929m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_275_930q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_282_931m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_276_932q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_283_933m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_277_934q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_284_935m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_278_936q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_285_937m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_279_938q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_286_939m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_27_434q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_34_435m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_280_940q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_287_941m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_281_942q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_288_943m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_282_944q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_289_945m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_283_946q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_290_947m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_284_948q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_291_949m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_285_950q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_292_951m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_286_952q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_293_953m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_287_954q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_294_955m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_288_956q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_295_957m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_289_958q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_296_959m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_28_436q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_35_437m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_290_960q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_297_961m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_291_962q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_298_963m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_292_964q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_299_965m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_293_966q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_300_967m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_294_968q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_301_969m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_295_970q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_302_971m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_296_972q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_303_973m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_29_438q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_36_439m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_2_384q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_9_385m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_30_440q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_37_441m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_31_442q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_38_443m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_32_444q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_39_445m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_33_446q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_40_447m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_34_448q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_41_449m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_35_450q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_42_451m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_36_452q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_43_453m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_37_454q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_44_455m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_38_456q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_45_457m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_39_458q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_46_459m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_3_386q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_10_387m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_40_460q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_47_461m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_41_462q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_48_463m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_42_464q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_49_465m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_43_466q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_50_467m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_44_468q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_51_469m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_45_470q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_52_471m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_46_472q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_53_473m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_47_474q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_54_475m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_48_476q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_55_477m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_49_478q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_56_479m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_4_388q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_11_389m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_50_480q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_57_481m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_51_482q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_58_483m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_52_484q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_59_485m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_53_486q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_60_487m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_54_488q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_61_489m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_55_490q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_62_491m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_56_492q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_63_493m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_57_494q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_64_495m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_58_496q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_65_497m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_59_498q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_66_499m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_5_390q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_12_391m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_60_500q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_67_501m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_61_502q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_68_503m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_62_504q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_69_505m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_63_506q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_70_507m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_64_508q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_71_509m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_65_510q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_72_511m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_66_512q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_73_513m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_67_514q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_74_515m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_68_516q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_75_517m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_69_518q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_76_519m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_6_392q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_13_393m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_70_520q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_77_521m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_71_522q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_78_523m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_72_524q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_79_525m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_73_526q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_80_527m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_74_528q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_81_529m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_75_530q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_82_531m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_76_532q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_83_533m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_77_534q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_84_535m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_78_536q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_85_537m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_79_538q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_86_539m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_7_394q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_14_395m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_80_540q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_87_541m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_81_542q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_88_543m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_82_544q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_89_545m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_83_546q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_90_547m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_84_548q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_91_549m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_85_550q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_92_551m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_86_552q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_93_553m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_87_554q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_94_555m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_88_556q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_95_557m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_89_558q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_96_559m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_8_396q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_15_397m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_90_560q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_97_561m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_91_562q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_98_563m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_92_564q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_99_565m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_93_566q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_100_567m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_94_568q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_101_569m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_95_570q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_102_571m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_96_572q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_103_573m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_97_574q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_104_575m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_98_576q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_105_577m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_99_578q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_106_579m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_9_398q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_16_399m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_187q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_1_193m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout;
				timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout;
		END IF;
	END PROCESS;
	wire_nO_w88w(0) <= NOT timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q;
	wire_nO_w80w(0) <= NOT timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q;
	wire_nO_w82w(0) <= NOT timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q;
	wire_nO_w84w(0) <= NOT timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_100_567m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_93_566q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_101_569m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_94_568q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_102_571m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_95_570q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_103_573m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_96_572q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_104_575m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_97_574q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_105_577m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_98_576q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_106_579m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_99_578q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_107_581m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_100_580q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_108_583m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_101_582q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_109_585m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_102_584q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_10_387m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_3_386q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_110_587m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_103_586q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_111_589m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_104_588q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_112_591m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_105_590q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_113_593m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_106_592q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_114_595m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_107_594q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_115_597m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_108_596q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_116_599m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_109_598q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_117_601m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_110_600q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_118_603m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_111_602q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_119_605m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_112_604q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_11_389m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_4_388q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_120_607m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_113_606q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_121_609m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_114_608q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_122_611m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_115_610q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_123_613m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_116_612q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_124_615m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_117_614q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_125_617m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_118_616q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_126_619m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_119_618q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_127_621m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_120_620q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_128_623m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_121_622q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_129_625m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_122_624q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_12_391m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_5_390q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_130_627m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_123_626q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_131_629m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_124_628q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_132_631m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_125_630q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_133_633m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_126_632q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_134_635m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_127_634q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_135_637m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_128_636q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_136_639m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_129_638q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_137_641m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_130_640q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_138_643m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_131_642q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_139_645m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_132_644q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_13_393m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_6_392q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_140_647m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_133_646q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_141_649m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_134_648q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_142_651m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_135_650q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_143_653m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_136_652q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_144_655m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_137_654q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_145_657m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_138_656q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_146_659m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_139_658q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_147_661m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_140_660q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_148_663m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_141_662q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_149_665m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_142_664q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_14_395m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_7_394q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_150_667m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_143_666q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_151_669m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_144_668q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_152_671m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_145_670q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_153_673m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_146_672q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_154_675m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_147_674q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_155_677m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_3_340_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_148_676q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_156_679m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_149_678q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_157_681m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_150_680q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_158_683m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_151_682q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_159_685m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_152_684q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_15_397m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_8_396q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_160_687m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_153_686q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_161_689m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_154_688q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_162_691m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_155_690q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_163_693m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_156_692q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_164_695m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_157_694q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_165_697m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_158_696q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_166_699m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_159_698q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_167_701m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_160_700q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_168_703m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_161_702q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_169_705m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_162_704q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_16_399m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_9_398q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_170_707m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_163_706q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_171_709m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_164_708q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_172_711m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_165_710q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_173_713m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_166_712q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_174_715m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_167_714q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_175_717m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_168_716q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_176_719m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_169_718q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_177_721m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_170_720q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_178_723m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_171_722q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_179_725m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_172_724q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_17_401m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_10_400q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_180_727m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_173_726q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_181_729m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_174_728q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_182_731m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_175_730q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_183_733m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_176_732q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_184_735m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_177_734q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_185_737m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_178_736q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_186_739m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_179_738q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_187_741m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_180_740q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_188_743m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_181_742q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_189_745m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_182_744q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_18_403m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_11_402q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_190_747m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_183_746q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_191_749m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_184_748q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_192_751m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_4_341_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_185_750q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_193_753m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_186_752q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_194_755m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_187_754q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_195_757m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_188_756q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_196_759m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_189_758q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_197_761m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_190_760q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_198_763m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_191_762q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_199_765m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_192_764q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_19_405m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_12_404q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_200_767m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_193_766q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_201_769m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_194_768q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_202_771m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_195_770q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_203_773m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_196_772q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_204_775m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_197_774q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_205_777m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_198_776q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_206_779m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_199_778q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_207_781m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_200_780q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_208_783m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_201_782q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_209_785m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_202_784q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_20_407m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_13_406q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_210_787m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_203_786q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_211_789m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_204_788q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_212_791m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_205_790q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_213_793m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_206_792q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_214_795m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_207_794q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_215_797m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_208_796q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_216_799m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_209_798q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_217_801m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_210_800q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_218_803m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_211_802q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_219_805m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_212_804q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_21_409m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_14_408q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_220_807m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_213_806q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_221_809m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_214_808q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_222_811m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_215_810q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_223_813m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_216_812q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_224_815m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_217_814q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_225_817m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_218_816q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_226_819m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_219_818q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_227_821m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_220_820q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_228_823m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_221_822q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_229_825m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_5_342_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_222_824q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_22_411m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_15_410q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_230_827m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_223_826q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_231_829m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_224_828q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_232_831m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_225_830q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_233_833m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_226_832q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_234_835m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_227_834q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_235_837m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_228_836q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_236_839m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_229_838q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_237_841m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_230_840q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_238_843m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_231_842q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_239_845m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_232_844q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_23_413m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_16_412q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_240_847m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_233_846q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_241_849m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_234_848q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_242_851m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_235_850q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_243_853m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_236_852q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_244_855m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_237_854q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_245_857m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_238_856q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_246_859m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_239_858q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_247_861m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_240_860q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_248_863m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_241_862q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_249_865m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_242_864q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_24_415m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_17_414q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_250_867m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_243_866q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_251_869m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_244_868q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_252_871m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_245_870q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_253_873m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_246_872q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_254_875m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_247_874q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_255_877m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_248_876q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_256_879m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_249_878q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_257_881m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_250_880q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_258_883m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_251_882q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_259_885m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_252_884q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_25_417m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_18_416q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_260_887m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_253_886q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_261_889m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_254_888q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_262_891m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_255_890q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_263_893m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_256_892q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_264_895m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_257_894q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_265_897m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_258_896q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_266_899m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_6_343_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_259_898q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_267_901m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_260_900q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_268_903m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_261_902q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_269_905m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_262_904q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_26_419m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_19_418q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_270_907m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_263_906q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_271_909m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_264_908q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_272_911m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_265_910q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_273_913m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_266_912q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_274_915m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_267_914q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_275_917m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_268_916q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_276_919m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_269_918q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_277_921m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_270_920q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_278_923m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_271_922q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_279_925m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_272_924q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_27_421m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_20_420q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_280_927m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_273_926q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_281_929m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_274_928q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_282_931m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_275_930q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_283_933m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_276_932q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_284_935m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_277_934q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_285_937m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_278_936q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_286_939m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_279_938q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_287_941m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_280_940q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_288_943m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_281_942q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_289_945m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_282_944q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_28_423m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_21_422q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_290_947m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_283_946q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_291_949m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_284_948q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_292_951m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_285_950q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_293_953m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_286_952q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_294_955m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_287_954q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_295_957m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_288_956q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_296_959m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_289_958q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_297_961m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_290_960q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_298_963m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_291_962q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_299_965m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_292_964q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_29_425m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_22_424q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_300_967m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_293_966q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_301_969m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_294_968q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_302_971m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_295_970q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_303_973m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_7_344_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_296_972q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_30_427m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_23_426q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_31_429m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_24_428q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_32_431m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_25_430q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_33_433m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_26_432q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_34_435m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_27_434q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_35_437m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_28_436q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_36_439m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_29_438q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_37_441m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_30_440q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_38_443m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_31_442q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_39_445m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_32_444q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_40_447m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_33_446q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_41_449m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_34_448q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_42_451m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_35_450q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_43_453m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_36_452q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_44_455m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_37_454q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_45_457m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_38_456q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_46_459m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_39_458q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_47_461m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_40_460q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_48_463m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_41_462q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_49_465m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_42_464q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_50_467m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_43_466q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_51_469m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_44_468q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_52_471m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_45_470q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_53_473m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_46_472q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_54_475m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_47_474q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_55_477m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_48_476q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_56_479m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_49_478q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_57_481m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_50_480q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_58_483m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_51_482q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_59_485m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_52_484q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_60_487m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_53_486q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_61_489m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_54_488q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_62_491m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_55_490q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_63_493m_dataout <= in_data(13) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_56_492q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_64_495m_dataout <= in_data(14) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_57_494q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_65_497m_dataout <= in_data(15) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_58_496q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_66_499m_dataout <= in_data(16) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_59_498q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_67_501m_dataout <= in_data(17) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_60_500q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_68_503m_dataout <= in_data(18) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_61_502q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_69_505m_dataout <= in_data(19) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_62_504q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_70_507m_dataout <= in_data(20) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_63_506q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_71_509m_dataout <= in_data(21) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_64_508q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_72_511m_dataout <= in_data(22) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_65_510q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_73_513m_dataout <= in_data(23) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_66_512q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_74_515m_dataout <= in_data(24) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_67_514q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_75_517m_dataout <= in_data(25) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_68_516q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_76_519m_dataout <= in_data(26) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_69_518q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_77_521m_dataout <= in_data(27) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_70_520q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_78_523m_dataout <= in_data(28) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_71_522q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_79_525m_dataout <= in_data(29) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_72_524q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_80_527m_dataout <= in_data(30) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_73_526q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_81_529m_dataout <= in_data(31) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_1_338_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_74_528q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_82_531m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_75_530q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_83_533m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_76_532q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_84_535m_dataout <= in_empty(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_77_534q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_85_537m_dataout <= in_endofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_78_536q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_86_539m_dataout <= in_startofpacket WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_79_538q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_87_541m_dataout <= in_data(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_80_540q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_88_543m_dataout <= in_data(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_81_542q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_89_545m_dataout <= in_data(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_82_544q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_8_383m_dataout <= in_error WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_1_382q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_90_547m_dataout <= in_data(3) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_83_546q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_91_549m_dataout <= in_data(4) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_84_548q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_92_551m_dataout <= in_data(5) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_85_550q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_93_553m_dataout <= in_data(6) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_86_552q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_94_555m_dataout <= in_data(7) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_87_554q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_95_557m_dataout <= in_data(8) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_88_556q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_96_559m_dataout <= in_data(9) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_89_558q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_97_561m_dataout <= in_data(10) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_90_560q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_98_563m_dataout <= in_data(11) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_91_562q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_99_565m_dataout <= in_data(12) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_2_339_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_92_564q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_9_385m_dataout <= in_empty(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_0_337_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_2_384q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_0_184m_dataout <= timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_204q AND NOT(s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_1_189m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_0_184m_dataout OR s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_3_981_dataout;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_2_192m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_1_189m_dataout WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout = '1'  ELSE wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_empty_0_184m_dataout;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_0_176m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_o(1) AND NOT(timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_1_175m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_o(2) AND NOT(timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_2_174m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_o(3) AND NOT(timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_0_180m_dataout <= timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q OR (((NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(0))) AND (NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(1)))) AND (NOT (timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q XOR wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o(2))));
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_1_185m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_0_180m_dataout WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_0_178_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_2_191m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_1_185m_dataout AND NOT(s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_4_334m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_2_191m_dataout WHEN wire_w106w(0) = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_full_205q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(0) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(1) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o(2) WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout = '1'  ELSE timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q;
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_0_190m_dataout <= wire_ni_w103w(0) AND NOT(s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_3_981_dataout);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_1_193m_dataout <= wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_out_valid_0_190m_dataout WHEN s_wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_always1_1_186_dataout = '1'  ELSE wire_ni_w103w(0);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_a <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_b <= ( "0" & "0" & "1");
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167 :  oper_add
	  GENERIC MAP (
		sgate_representation => 0,
		width_a => 3,
		width_b => 3,
		width_o => 3
	  )
	  PORT MAP ( 
		a => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_a,
		b => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_b,
		cin => wire_gnd,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add0_167_o
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_a <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_2_201q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_1_202q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_rd_addr_0_203q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_b <= ( "0" & "0" & "1");
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168 :  oper_add
	  GENERIC MAP (
		sgate_representation => 0,
		width_a => 3,
		width_b => 3,
		width_o => 3
	  )
	  PORT MAP ( 
		a => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_a,
		b => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_b,
		cin => wire_gnd,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add1_168_o
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_a <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q & "1");
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_b <= ( wire_nO_w84w & wire_nO_w82w & wire_nO_w80w & "1");
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172 :  oper_add
	  GENERIC MAP (
		sgate_representation => 0,
		width_a => 4,
		width_b => 4,
		width_o => 4
	  )
	  PORT MAP ( 
		a => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_a,
		b => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_b,
		cin => wire_gnd,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_add2_172_o
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_i <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_2_198q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_1_199q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_wr_addr_0_200q);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336 :  oper_decoder
	  GENERIC MAP (
		width_i => 3,
		width_o => 8
	  )
	  PORT MAP ( 
		i => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_i,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_336_o
	  );
	wire_timing_adapter_32_lessthan0_2_a <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_2_174m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_1_175m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_fill_level_0_176m_dataout);
	wire_timing_adapter_32_lessthan0_2_b <= ( "0" & "1" & "1");
	timing_adapter_32_lessthan0_2 :  oper_less_than
	  GENERIC MAP (
		sgate_representation => 0,
		width_a => 3,
		width_b => 3
	  )
	  PORT MAP ( 
		a => wire_timing_adapter_32_lessthan0_2_a,
		b => wire_timing_adapter_32_lessthan0_2_b,
		cin => wire_gnd,
		o => wire_timing_adapter_32_lessthan0_2_o
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_260_900q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_223_826q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_186_752q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_149_678q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_112_604q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_75_530q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_38_456q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_1_382q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_345_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_261_902q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_224_828q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_187_754q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_150_680q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_113_606q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_76_532q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_39_458q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_2_384q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_346_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_262_904q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_225_830q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_188_756q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_151_682q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_114_608q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_77_534q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_40_460q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_3_386q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_347_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_263_906q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_226_832q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_189_758q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_152_684q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_115_610q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_78_536q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_41_462q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_4_388q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_348_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_264_908q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_227_834q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_190_760q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_153_686q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_116_612q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_79_538q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_42_464q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_5_390q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_349_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_265_910q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_228_836q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_191_762q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_154_688q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_117_614q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_80_540q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_43_466q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_6_392q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_350_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_266_912q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_229_838q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_192_764q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_155_690q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_118_616q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_81_542q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_44_468q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_7_394q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_351_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_267_914q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_230_840q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_193_766q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_156_692q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_119_618q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_82_544q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_45_470q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_8_396q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_352_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_268_916q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_231_842q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_194_768q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_157_694q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_120_620q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_83_546q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_46_472q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_9_398q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_353_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_269_918q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_232_844q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_195_770q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_158_696q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_121_622q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_84_548q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_47_474q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_10_400q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_354_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_270_920q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_233_846q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_196_772q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_159_698q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_122_624q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_85_550q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_48_476q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_11_402q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_355_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_271_922q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_234_848q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_197_774q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_160_700q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_123_626q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_86_552q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_49_478q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_12_404q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_356_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_272_924q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_235_850q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_198_776q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_161_702q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_124_628q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_87_554q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_50_480q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_13_406q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_357_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_273_926q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_236_852q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_199_778q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_162_704q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_125_630q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_88_556q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_51_482q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_14_408q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_358_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_274_928q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_237_854q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_200_780q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_163_706q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_126_632q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_89_558q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_52_484q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_15_410q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_359_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_275_930q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_238_856q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_201_782q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_164_708q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_127_634q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_90_560q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_53_486q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_16_412q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_360_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_276_932q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_239_858q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_202_784q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_165_710q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_128_636q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_91_562q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_54_488q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_17_414q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_361_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_277_934q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_240_860q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_203_786q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_166_712q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_129_638q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_92_564q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_55_490q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_18_416q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_362_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_278_936q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_241_862q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_204_788q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_167_714q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_130_640q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_93_566q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_56_492q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_19_418q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_363_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_279_938q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_242_864q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_205_790q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_168_716q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_131_642q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_94_568q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_57_494q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_20_420q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_364_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_280_940q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_243_866q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_206_792q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_169_718q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_132_644q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_95_570q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_58_496q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_21_422q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_365_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_281_942q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_244_868q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_207_794q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_170_720q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_133_646q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_96_572q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_59_498q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_22_424q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_366_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_282_944q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_245_870q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_208_796q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_171_722q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_134_648q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_97_574q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_60_500q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_23_426q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_367_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_283_946q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_246_872q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_209_798q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_172_724q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_135_650q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_98_576q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_61_502q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_24_428q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_368_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_284_948q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_247_874q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_210_800q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_173_726q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_136_652q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_99_578q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_62_504q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_25_430q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_369_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_285_950q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_248_876q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_211_802q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_174_728q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_137_654q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_100_580q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_63_506q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_26_432q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_370_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_286_952q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_249_878q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_212_804q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_175_730q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_138_656q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_101_582q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_64_508q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_27_434q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_371_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_287_954q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_250_880q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_213_806q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_176_732q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_139_658q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_102_584q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_65_510q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_28_436q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_372_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_288_956q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_251_882q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_214_808q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_177_734q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_140_660q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_103_586q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_66_512q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_29_438q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_373_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_289_958q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_252_884q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_215_810q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_178_736q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_141_662q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_104_588q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_67_514q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_30_440q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_374_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_290_960q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_253_886q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_216_812q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_179_738q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_142_664q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_105_590q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_68_516q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_31_442q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_375_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_291_962q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_254_888q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_217_814q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_180_740q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_143_666q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_106_592q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_69_518q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_32_444q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_376_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_292_964q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_255_890q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_218_816q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_181_742q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_144_668q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_107_594q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_70_520q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_33_446q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_377_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_293_966q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_256_892q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_219_818q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_182_744q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_145_670q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_108_596q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_71_522q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_34_448q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_378_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_294_968q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_257_894q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_220_820q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_183_746q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_146_672q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_109_598q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_72_524q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_35_450q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_379_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_295_970q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_258_896q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_221_822q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_184_748q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_147_674q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_110_600q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_73_526q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_36_452q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_380_sel
	  );
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_data <= ( timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_296_972q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_259_898q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_222_824q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_185_750q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_148_676q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_111_602q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_74_528q & timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_37_454q);
	wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_sel <= ( wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_2_206m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_1_207m_dataout & wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_rd_addr_0_208m_dataout);
	timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381 :  oper_mux
	  GENERIC MAP (
		width_data => 8,
		width_sel => 3
	  )
	  PORT MAP ( 
		data => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_data,
		o => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_o,
		sel => wire_timing_adapter_32_timing_adapter_fifo_32_timing_adapter_fifo_mem_381_sel
	  );

 END RTL; --timing_adapter_32
 --synopsys translate_on
--VALID FILE
