2800
0a00
0003
