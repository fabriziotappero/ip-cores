library verilog;
use verilog.vl_types.all;
entity pc_gen_ctl_reg_clr is
    port(
        pc_gen_ctl_i    : in     vl_logic_vector(2 downto 0);
        pc_gen_ctl_o    : out    vl_logic_vector(2 downto 0);
        clk             : in     vl_logic;
        clr             : in     vl_logic;
        hold            : in     vl_logic
    );
end pc_gen_ctl_reg_clr;
