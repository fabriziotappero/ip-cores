----------------------------------------------------------------------
----                                                              ----
----  cod3_synth.vhd                                              ----
----                                                              ----
----  This file is part of the turbo decoder IP core project      ----
----  http://www.opencores.org/projects/turbocodes/               ----
----                                                              ----
----  Author(s):                                                  ----
----      - David Brochart(dbrochart@opencores.org)               ----
----                                                              ----
----  All additional information is available in the README.txt   ----
----  file.                                                       ----
----                                                              ----
----------------------------------------------------------------------
----                                                              ----
---- Copyright (C) 2005 Authors                                   ----
----                                                              ----
---- This source file may be used and distributed without         ----
---- restriction provided that this copyright statement is not    ----
---- removed from the file and that any derivative work contains  ----
---- the original copyright notice and the associated disclaimer. ----
----                                                              ----
---- This source file is free software; you can redistribute it   ----
---- and/or modify it under the terms of the GNU Lesser General   ----
---- Public License as published by the Free Software Foundation; ----
---- either version 2.1 of the License, or (at your option) any   ----
---- later version.                                               ----
----                                                              ----
---- This source is distributed in the hope that it will be       ----
---- useful, but WITHOUT ANY WARRANTY; without even the implied   ----
---- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ----
---- PURPOSE. See the GNU Lesser General Public License for more  ----
---- details.                                                     ----
----                                                              ----
---- You should have received a copy of the GNU Lesser General    ----
---- Public License along with this source; if not, download it   ----
---- from http://www.opencores.org/lgpl.shtml                     ----
----                                                              ----
----------------------------------------------------------------------



architecture synth of cod3 is
begin
    process (inSig)
        variable tmp : std_logic_vector(2 downto 0);
    begin
        tmp(0) := ((not inSig(6)) and (not inSig(5)) and (not inSig(3))) or ((not inSig(6)) and inSig(5) and (not inSig(2))) or (inSig(6) and (not inSig(4)) and (not inSig(1))) or ((inSig(6)) and (inSig(4)) and (not inSig(0)));
        tmp(1) := ((not inSig(6)) and (not inSig(5))) or (inSig(6) and (not inSig(4)));
        tmp(2) := not inSig(6);
        outCod <= tmp;
    end process;
end;
