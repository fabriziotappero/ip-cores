-------------------------------------------------------------------------------
-- $Id: ram_loader-c.vhd 77 2009-04-01 19:53:14Z arniml $
-------------------------------------------------------------------------------

configuration ram_loader_rtl_c0 of ram_loader is

  for rtl
  end for;

end ram_loader_rtl_c0;
