// ===========================================================================
// File    : crc32d16N.v
// Author  : cwinward
// Date    : Sat Dec 8 14:00:37 MST 2007
// Project : TI PHY design
//
// Copyright (c) notice
// This code adheres to the GNU public license
//
// ===========================================================================
//
// $Id: crc32d16.v,v 1.1.1.1 2007-12-08 22:27:00 cmagleby Exp $
//
// ===========================================================================
//
// $Log: not supported by cvs2svn $
//
// ===========================================================================
// Function :  CRC for TLP packet
//             This was generated by a c program owned by gutzlogic.
// ===========================================================================
// ===========================================================================


module crc32d16(/*AUTOARG*/
   // Outputs
   crc, 
   // Inputs
   clk, resetN, load, d, init,en
   );


   input clk;
   input resetN;
   input load;
   input [15:0] d;
   input [31:0] init;
   input        en;
   output [31:0] crc;
   reg [31:0]    crc;
   

   always @(posedge clk or negedge resetN)
     begin
        if(~resetN)
          crc <= #1 32'hFFFF_FFFF;
        else if(load)
          crc <= #1 init;
        else
          if(en)
            begin
               crc[0] <= #1 d[3] ^ d[5] ^ d[6] ^ d[9] ^ d[15] ^ crc[16] ^ crc[22] ^ crc[25] ^ crc[26] 
              ^ crc[28];
               crc[1] <= #1 d[2] ^ d[3] ^ d[4] ^ d[6] ^ d[8] ^ d[9] ^ d[14] ^ d[15] ^ crc[16] ^ 
                         crc[17] ^ crc[22] ^ crc[23] ^ crc[25] ^ crc[27] ^ crc[28] ^ crc[29];
               crc[2] <= #1 d[1] ^ d[2] ^ d[6] ^ d[7] ^ d[8] ^ d[9] ^ d[13] ^ d[14] ^ d[15] ^ 
                         crc[16] ^ crc[17] ^ crc[18] ^ crc[22] ^ crc[23] ^ crc[24] ^ crc[25] ^ crc[29] ^ crc[30];
               crc[3] <= #1 d[0] ^ d[1] ^ d[5] ^ d[6] ^ d[7] ^ d[8] ^ d[12] ^ d[13] ^ d[14] ^ 
                         crc[17] ^ crc[18] ^ crc[19] ^ crc[23] ^ crc[24] ^ crc[25] ^ crc[26] ^ crc[30] ^ crc[31];
               crc[4] <= #1 d[0] ^ d[3] ^ d[4] ^ d[7] ^ d[9] ^ d[11] ^ d[12] ^ d[13] ^ d[15] ^ 
                         crc[16] ^ crc[18] ^ crc[19] ^ crc[20] ^ crc[22] ^ crc[24] ^ crc[27] ^ crc[28] ^ crc[31];
               crc[5] <= #1 d[2] ^ d[5] ^ d[8] ^ d[9] ^ d[10] ^ d[11] ^ d[12] ^ d[14] ^ d[15] 
                 ^ crc[16] ^ crc[17] ^ crc[19] ^ crc[20] ^ crc[21] ^ crc[22] ^ crc[23] ^ crc[26] ^ 
                         crc[29];
               crc[6] <= #1 d[1] ^ d[4] ^ d[7] ^ d[8] ^ d[9] ^ d[10] ^ d[11] ^ d[13] ^ d[14] ^ 
                         crc[17] ^ crc[18] ^ crc[20] ^ crc[21] ^ crc[22] ^ crc[23] ^ crc[24] ^ crc[27] ^ crc[30];
               crc[7] <= #1 d[0] ^ d[5] ^ d[7] ^ d[8] ^ d[10] ^ d[12] ^ d[13] ^ d[15] ^ crc[16] 
                 ^ crc[18] ^ crc[19] ^ crc[21] ^ crc[23] ^ crc[24] ^ crc[26] ^ crc[31];
               crc[8] <= #1 d[3] ^ d[4] ^ d[5] ^ d[7] ^ d[11] ^ d[12] ^ d[14] ^ d[15] ^ crc[16] 
                 ^ crc[17] ^ crc[19] ^ crc[20] ^ crc[24] ^ crc[26] ^ crc[27] ^ crc[28];
               crc[9] <= #1 d[2] ^ d[3] ^ d[4] ^ d[6] ^ d[10] ^ d[11] ^ d[13] ^ d[14] ^ crc[17] 
                 ^ crc[18] ^ crc[20] ^ crc[21] ^ crc[25] ^ crc[27] ^ crc[28] ^ crc[29];
               crc[10] <= #1 d[1] ^ d[2] ^ d[6] ^ d[10] ^ d[12] ^ d[13] ^ d[15] ^ crc[16] ^ crc[18] 
                 ^ crc[19] ^ crc[21] ^ crc[25] ^ crc[29] ^ crc[30];
               crc[11] <= #1 d[0] ^ d[1] ^ d[3] ^ d[6] ^ d[11] ^ d[12] ^ d[14] ^ d[15] ^ crc[16] 
                 ^ crc[17] ^ crc[19] ^ crc[20] ^ crc[25] ^ crc[28] ^ crc[30] ^ crc[31];
               crc[12] <= #1 d[0] ^ d[2] ^ d[3] ^ d[6] ^ d[9] ^ d[10] ^ d[11] ^ d[13] ^ d[14] ^ 
                          d[15] ^ crc[16] ^ crc[17] ^ crc[18] ^ crc[20] ^ crc[21] ^ crc[22] ^ crc[25] ^ crc[28] 
                 ^ crc[29] ^ crc[31];
               crc[13] <= #1 d[1] ^ d[2] ^ d[5] ^ d[8] ^ d[9] ^ d[10] ^ d[12] ^ d[13] ^ d[14] ^ 
                          crc[17] ^ crc[18] ^ crc[19] ^ crc[21] ^ crc[22] ^ crc[23] ^ crc[26] ^ crc[29] ^ crc[30];
               crc[14] <= #1 d[0] ^ d[1] ^ d[4] ^ d[7] ^ d[8] ^ d[9] ^ d[11] ^ d[12] ^ d[13] ^ 
                          crc[18] ^ crc[19] ^ crc[20] ^ crc[22] ^ crc[23] ^ crc[24] ^ crc[27] ^ crc[30] ^ crc[31];
               crc[15] <= #1 d[0] ^ d[3] ^ d[6] ^ d[7] ^ d[8] ^ d[10] ^ d[11] ^ d[12] ^ crc[19] ^ 
                          crc[20] ^ crc[21] ^ crc[23] ^ crc[24] ^ crc[25] ^ crc[28] ^ crc[31];
               crc[16] <= #1 d[2] ^ d[3] ^ d[7] ^ d[10] ^ d[11] ^ d[15] ^ crc[0] ^ crc[16] ^ crc[20] 
                 ^ crc[21] ^ crc[24] ^ crc[28] ^ crc[29];
               crc[17] <= #1 d[1] ^ d[2] ^ d[6] ^ d[9] ^ d[10] ^ d[14] ^ crc[1] ^ crc[17] ^ crc[21] ^ 
                          crc[22] ^ crc[25] ^ crc[29] ^ crc[30];
               crc[18] <= #1 d[0] ^ d[1] ^ d[5] ^ d[8] ^ d[9] ^ d[13] ^ crc[2] ^ crc[18] ^ crc[22] ^ 
                          crc[23] ^ crc[26] ^ crc[30] ^ crc[31];
               crc[19] <= #1 d[0] ^ d[4] ^ d[7] ^ d[8] ^ d[12] ^ crc[3] ^ crc[19] ^ crc[23] ^ crc[24] ^ 
                          crc[27] ^ crc[31];
               crc[20] <= #1 d[3] ^ d[6] ^ d[7] ^ d[11] ^ crc[4] ^ crc[20] ^ crc[24] ^ crc[25] ^ crc[28];
               crc[21] <= #1 d[2] ^ d[5] ^ d[6] ^ d[10] ^ crc[5] ^ crc[21] ^ crc[25] ^ crc[26] ^ crc[29];
               crc[22] <= #1 d[1] ^ d[3] ^ d[4] ^ d[6] ^ d[15] ^ crc[6] ^ crc[16] ^ crc[25] ^ crc[27] ^ 
                          crc[28] ^ crc[30];
               crc[23] <= #1 d[0] ^ d[2] ^ d[6] ^ d[9] ^ d[14] ^ d[15] ^ crc[7] ^ crc[16] ^ crc[17] ^ 
                          crc[22] ^ crc[25] ^ crc[29] ^ crc[31];
               crc[24] <= #1 d[1] ^ d[5] ^ d[8] ^ d[13] ^ d[14] ^ crc[8] ^ crc[17] ^ crc[18] ^ crc[23] 
                 ^ crc[26] ^ crc[30];
               crc[25] <= #1 d[0] ^ d[4] ^ d[7] ^ d[12] ^ d[13] ^ crc[9] ^ crc[18] ^ crc[19] ^ crc[24] 
                 ^ crc[27] ^ crc[31];
               crc[26] <= #1 d[5] ^ d[9] ^ d[11] ^ d[12] ^ d[15] ^ crc[10] ^ crc[16] ^ crc[19] ^ crc[20] 
                 ^ crc[22] ^ crc[26];
               crc[27] <= #1 d[4] ^ d[8] ^ d[10] ^ d[11] ^ d[14] ^ crc[11] ^ crc[17] ^ crc[20] ^ crc[21] 
                 ^ crc[23] ^ crc[27];
               crc[28] <= #1 d[3] ^ d[7] ^ d[9] ^ d[10] ^ d[13] ^ crc[12] ^ crc[18] ^ crc[21] ^ crc[22] 
                 ^ crc[24] ^ crc[28];
               crc[29] <= #1 d[2] ^ d[6] ^ d[8] ^ d[9] ^ d[12] ^ crc[13] ^ crc[19] ^ crc[22] ^ crc[23] 
                 ^ crc[25] ^ crc[29];
               crc[30] <= #1 d[1] ^ d[5] ^ d[7] ^ d[8] ^ d[11] ^ crc[14] ^ crc[20] ^ crc[23] ^ crc[24] 
                 ^ crc[26] ^ crc[30];
               crc[31] <= #1 d[0] ^ d[4] ^ d[6] ^ d[7] ^ d[10] ^ crc[15] ^ crc[21] ^ crc[24] ^ crc[25] 
                 ^ crc[27] ^ crc[31];
            end // if (en)
          else
            crc <= #1 crc;
     end
        
endmodule


