-- SVGA controller
  constant CFG_SVGA_ENABLE : integer := CONFIG_SVGA_ENABLE;

