////////////////////////////////////////////////////////////////////////////
//
// Copyright 2014  Ken Campbell
//
//   Licensed under the Apache License, Version 2.0 (the "License");
//   you may not use this file except in compliance with the License.
//   You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in writing, software
//   distributed under the License is distributed on an "AS IS" BASIS,
//   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//   See the License for the specific language governing permissions and
//   limitations under the License.
//
/////////////////////////////////////

/////////////////////////////////////////////////////////
//  the test bench package.
//
package tb_pkg;

  `include "tb_types.sv"
  `include "gfuncts.sv"
  `include "lst_item.sv"
  `include "tb_cmd.sv"
  `include "cmd_lst.sv"
  
endpackage:  tb_pkg // tb
  
