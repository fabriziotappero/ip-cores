Paste timesim model here