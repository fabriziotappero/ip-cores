-- DDRMP controller
  constant CFG_DDRMP_EN  	: integer := CONFIG_DDRMP;
  constant CFG_DDRMP_EN2P    	: integer := CONFIG_DDRMP_EN2P;
  constant CFG_DDRMP_NCS    	: integer := CONFIG_DDRMP_NCS;
  constant CFG_DDRMP_NDEV    	: integer := CONFIG_DDRMP_NDEV;
  constant CFG_DDRMP_NBITS    	: integer := CONFIG_DDRMP_NBITS;
  constant CFG_DDRMP_MBITS    	: integer := CONFIG_DDRMP_MBITS;
  constant CFG_DDRMP_PERIOD    	: integer := 1000/CONFIG_DDRMP_FREQ;

