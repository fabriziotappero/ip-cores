    vector_stim_in : process ( clock_tb )
                    variable i  : integer := 0;
type out_vector is record
      A           : std_logic_vector(8 downto 1)    ;
      B           : std_logic_vector(8 downto 1)    ;
      S           : std_logic_vector(4 downto 1)    ;
      Y           : std_logic_vector(8 downto 1)    ;
      CLR         : std_logic                       ;
      CLK         : std_logic                       ;
      C           : std_logic                       ;
      V           : std_logic                       ;
      Z           : std_logic                       ;
 end record;
type out_vectors is array (natural range <>) of out_vector;
constant vectors  : out_vectors :=  (
("UUUUUUUU", "UUUUUUUU", "UUUU", "UUUUUUUU", '1', '1', 'U', 'U', 'U'),
("01010101", "00000001", "0000", "00000000", '1', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "00000000", '1', '1', '0', '0', '0'),
("01010101", "00000010", "0000", "00000000", '1', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "00000000", '1', '1', '0', '0', '0'),
("01010101", "00000100", "0000", "00000000", '0', '1', '0', '0', '0'),
("01010101", "00000100", "0000", "00000000", '0', '1', '0', '0', '0'),
("01010101", "00000100", "0000", "00000000", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "01011001", '0', '1', '0', '0', '0'),
("01010101", "00001000", "0000", "01011001", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00010000", "0000", "01011101", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00100000", "0000", "01100101", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "01010101", '0', '1', '0', '0', '0'),
("01010101", "01000000", "0000", "01110101", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0000", "01010101", '0', '1', '0', '0', '0'),
("01010101", "10000000", "0000", "10010101", '0', '1', '0', '0', '0'),
("01010101", "00000001", "0010", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0010", "11010101", '0', '1', '0', '0', '0'),
("01010101", "00000010", "0010", "01010100", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0010", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00000100", "0010", "01010011", '0', '1', '0', '0', '0'),
("01010101", "00010000", "0010", "01010101", '0', '1', '0', '0', '0'),
("01010101", "01000000", "0010", "01010001", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0010", "01000101", '0', '1', '0', '0', '0'),
("01010101", "10000000", "0010", "00010101", '0', '1', '0', '0', '0'),
("01010101", "00000001", "0100", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0100", "11010101", '0', '1', '0', '0', '0'),
("01010101", "00000010", "0101", "10101010", '0', '1', '0', '0', '0'),
("01010101", "00000000", "0101", "01010101", '0', '1', '0', '0', '0'),
("01010101", "00000100", "0100", "00010101", '0', '1', '0', '0', '0'),
("01010101", "00010000", "0101", "01010101", '0', '1', '0', '0', '0'),
("01010101", "01000000", "0010", "01010000", '0', '1', '1', '0', '0'),
("01010101", "00000000", "0010", "01010101", '0', '1', '0', '0', '0'),
("01010101", "10000000", "0010", "00010101", '0', '1', '0', '0', '0'),
("01010101", "10000000", "0010", "01010101", '0', '1', '0', '0', '0'));
                 begin
                    if (clock_tb'event and clock_tb = '1') then
                        if ( i <= vectors'high) then
                            A <= vectors(i).A;
                            B <= vectors(i).B;
                            S <= vectors(i).S;
                            --Y <= vectors(i).Y;
                            CLR <= vectors(i).CLR;
                            CLK <= vectors(i).CLK;
                            --C <= vectors(i).C;
                            --V <= vectors(i).V;
                            --Z <= vectors(i).Z;
                            
                            i := i + 1;
                        else
                            finished <= '1';
                        end if;
                    else
                        CLK <= clock_tb;
                    end if;

                end process vector_stim_in;

