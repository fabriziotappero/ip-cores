/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

/* v0(a)+v1(a)+v2(a) == a^3 in GF(3^m) */

/* c == v0(a) */
module v0(a, c);
    input [193:0] a;
    output [193:0] c;
    assign c[1:0] = a[1:0];
    assign c[3:2] = a[131:130];
    assign c[5:4] = a[67:66];
    assign c[7:6] = a[3:2];
    assign c[9:8] = a[133:132];
    assign c[11:10] = a[69:68];
    assign c[13:12] = a[5:4];
    assign c[15:14] = a[135:134];
    assign c[17:16] = a[71:70];
    assign c[19:18] = a[193:192];
    assign c[21:20] = {a[128], a[129]};
    assign c[23:22] = a[73:72];
    assign c[25:24] = {a[178], a[179]};
    assign c[27:26] = a[131:130];
    assign c[29:28] = {a[66], a[67]};
    assign c[31:30] = {a[180], a[181]};
    assign c[33:32] = a[133:132];
    assign c[35:34] = {a[68], a[69]};
    assign c[37:36] = {a[182], a[183]};
    assign c[39:38] = a[127:126];
    assign c[41:40] = {a[70], a[71]};
    assign c[43:42] = {a[184], a[185]};
    assign c[45:44] = a[145:144];
    assign c[47:46] = a[81:80];
    assign c[49:48] = a[17:16];
    assign c[51:50] = a[147:146];
    assign c[53:52] = a[83:82];
    assign c[55:54] = a[19:18];
    assign c[57:56] = a[149:148];
    assign c[59:58] = a[85:84];
    assign c[61:60] = a[21:20];
    assign c[63:62] = a[135:134];
    assign c[65:64] = a[87:86];
    assign c[67:66] = {a[192], a[193]};
    assign c[69:68] = a[145:144];
    assign c[71:70] = {a[80], a[81]};
    assign c[73:72] = a[25:24];
    assign c[75:74] = a[147:146];
    assign c[77:76] = {a[82], a[83]};
    assign c[79:78] = a[27:26];
    assign c[81:80] = a[149:148];
    assign c[83:82] = {a[84], a[85]};
    assign c[85:84] = a[29:28];
    assign c[87:86] = a[143:142];
    assign c[89:88] = {a[86], a[87]};
    assign c[91:90] = a[31:30];
    assign c[93:92] = a[161:160];
    assign c[95:94] = a[97:96];
    assign c[97:96] = a[33:32];
    assign c[99:98] = a[163:162];
    assign c[101:100] = a[99:98];
    assign c[103:102] = a[35:34];
    assign c[105:104] = a[165:164];
    assign c[107:106] = a[101:100];
    assign c[109:108] = a[37:36];
    assign c[111:110] = a[151:150];
    assign c[113:112] = a[103:102];
    assign c[115:114] = a[39:38];
    assign c[117:116] = a[161:160];
    assign c[119:118] = {a[96], a[97]};
    assign c[121:120] = a[41:40];
    assign c[123:122] = a[163:162];
    assign c[125:124] = {a[98], a[99]};
    assign c[127:126] = a[43:42];
    assign c[129:128] = a[165:164];
    assign c[131:130] = {a[100], a[101]};
    assign c[133:132] = a[45:44];
    assign c[135:134] = a[159:158];
    assign c[137:136] = {a[102], a[103]};
    assign c[139:138] = a[47:46];
    assign c[141:140] = a[177:176];
    assign c[143:142] = a[113:112];
    assign c[145:144] = a[49:48];
    assign c[147:146] = a[179:178];
    assign c[149:148] = a[115:114];
    assign c[151:150] = a[51:50];
    assign c[153:152] = a[181:180];
    assign c[155:154] = a[117:116];
    assign c[157:156] = a[53:52];
    assign c[159:158] = a[167:166];
    assign c[161:160] = a[119:118];
    assign c[163:162] = a[55:54];
    assign c[165:164] = a[177:176];
    assign c[167:166] = {a[112], a[113]};
    assign c[169:168] = a[57:56];
    assign c[171:170] = a[179:178];
    assign c[173:172] = {a[114], a[115]};
    assign c[175:174] = a[59:58];
    assign c[177:176] = a[181:180];
    assign c[179:178] = {a[116], a[117]};
    assign c[181:180] = a[61:60];
    assign c[183:182] = a[175:174];
    assign c[185:184] = {a[118], a[119]};
    assign c[187:186] = a[63:62];
    assign c[189:188] = a[193:192];
    assign c[191:190] = a[129:128];
    assign c[193:192] = a[65:64];
endmodule
/* c == v1(a) */
module v1(a, c);
    input [193:0] a;
    output [193:0] c;
    assign c[1:0] = a[179:178];
    assign c[3:2] = {a[122], a[123]};
    assign c[5:4] = 0;
    assign c[7:6] = a[181:180];
    assign c[9:8] = {a[124], a[125]};
    assign c[11:10] = 0;
    assign c[13:12] = a[183:182];
    assign c[15:14] = {a[126], a[127]};
    assign c[17:16] = 0;
    assign c[19:18] = a[7:6];
    assign c[21:20] = a[137:136];
    assign c[23:22] = 0;
    assign c[25:24] = a[9:8];
    assign c[27:26] = a[139:138];
    assign c[29:28] = a[75:74];
    assign c[31:30] = a[11:10];
    assign c[33:32] = a[125:124];
    assign c[35:34] = a[77:76];
    assign c[37:36] = a[13:12];
    assign c[39:38] = a[135:134];
    assign c[41:40] = a[79:78];
    assign c[43:42] = a[15:14];
    assign c[45:44] = a[129:128];
    assign c[47:46] = {a[72], a[73]};
    assign c[49:48] = {a[186], a[187]};
    assign c[51:50] = a[139:138];
    assign c[53:52] = {a[74], a[75]};
    assign c[55:54] = {a[188], a[189]};
    assign c[57:56] = a[133:132];
    assign c[59:58] = {a[76], a[77]};
    assign c[61:60] = {a[190], a[191]};
    assign c[63:62] = a[151:150];
    assign c[65:64] = {a[78], a[79]};
    assign c[67:66] = a[23:22];
    assign c[69:68] = a[137:136];
    assign c[71:70] = a[89:88];
    assign c[73:72] = 0;
    assign c[75:74] = a[155:154];
    assign c[77:76] = a[91:90];
    assign c[79:78] = 0;
    assign c[81:80] = a[141:140];
    assign c[83:82] = a[93:92];
    assign c[85:84] = 0;
    assign c[87:86] = a[151:150];
    assign c[89:88] = a[95:94];
    assign c[91:90] = 0;
    assign c[93:92] = a[145:144];
    assign c[95:94] = {a[88], a[89]};
    assign c[97:96] = 0;
    assign c[99:98] = a[155:154];
    assign c[101:100] = {a[90], a[91]};
    assign c[103:102] = 0;
    assign c[105:104] = a[149:148];
    assign c[107:106] = {a[92], a[93]};
    assign c[109:108] = 0;
    assign c[111:110] = a[167:166];
    assign c[113:112] = {a[94], a[95]};
    assign c[115:114] = 0;
    assign c[117:116] = a[153:152];
    assign c[119:118] = a[105:104];
    assign c[121:120] = 0;
    assign c[123:122] = a[171:170];
    assign c[125:124] = a[107:106];
    assign c[127:126] = 0;
    assign c[129:128] = a[157:156];
    assign c[131:130] = a[109:108];
    assign c[133:132] = 0;
    assign c[135:134] = a[167:166];
    assign c[137:136] = a[111:110];
    assign c[139:138] = 0;
    assign c[141:140] = a[161:160];
    assign c[143:142] = {a[104], a[105]};
    assign c[145:144] = 0;
    assign c[147:146] = a[171:170];
    assign c[149:148] = {a[106], a[107]};
    assign c[151:150] = 0;
    assign c[153:152] = a[165:164];
    assign c[155:154] = {a[108], a[109]};
    assign c[157:156] = 0;
    assign c[159:158] = a[183:182];
    assign c[161:160] = {a[110], a[111]};
    assign c[163:162] = 0;
    assign c[165:164] = a[169:168];
    assign c[167:166] = a[121:120];
    assign c[169:168] = 0;
    assign c[171:170] = a[187:186];
    assign c[173:172] = a[123:122];
    assign c[175:174] = 0;
    assign c[177:176] = a[173:172];
    assign c[179:178] = a[125:124];
    assign c[181:180] = 0;
    assign c[183:182] = a[183:182];
    assign c[185:184] = a[127:126];
    assign c[187:186] = 0;
    assign c[189:188] = a[177:176];
    assign c[191:190] = {a[120], a[121]};
    assign c[193:192] = 0;
endmodule
/* c == v2(a) */
module v2(a, c);
    input [193:0] a;
    output [193:0] c;
    assign c[1:0] = a[187:186];
    assign c[3:2] = 0;
    assign c[5:4] = 0;
    assign c[7:6] = a[189:188];
    assign c[9:8] = 0;
    assign c[11:10] = 0;
    assign c[13:12] = a[191:190];
    assign c[15:14] = 0;
    assign c[17:16] = 0;
    assign c[19:18] = a[185:184];
    assign c[21:20] = 0;
    assign c[23:22] = 0;
    assign c[25:24] = 0;
    assign c[27:26] = a[123:122];
    assign c[29:28] = 0;
    assign c[31:30] = 0;
    assign c[33:32] = a[141:140];
    assign c[35:34] = 0;
    assign c[37:36] = 0;
    assign c[39:38] = a[143:142];
    assign c[41:40] = 0;
    assign c[43:42] = 0;
    assign c[45:44] = a[137:136];
    assign c[47:46] = 0;
    assign c[49:48] = 0;
    assign c[51:50] = a[131:130];
    assign c[53:52] = 0;
    assign c[55:54] = 0;
    assign c[57:56] = a[141:140];
    assign c[59:58] = 0;
    assign c[61:60] = 0;
    assign c[63:62] = a[143:142];
    assign c[65:64] = 0;
    assign c[67:66] = 0;
    assign c[69:68] = a[153:152];
    assign c[71:70] = 0;
    assign c[73:72] = 0;
    assign c[75:74] = a[139:138];
    assign c[77:76] = 0;
    assign c[79:78] = 0;
    assign c[81:80] = a[157:156];
    assign c[83:82] = 0;
    assign c[85:84] = 0;
    assign c[87:86] = a[159:158];
    assign c[89:88] = 0;
    assign c[91:90] = 0;
    assign c[93:92] = a[153:152];
    assign c[95:94] = 0;
    assign c[97:96] = 0;
    assign c[99:98] = a[147:146];
    assign c[101:100] = 0;
    assign c[103:102] = 0;
    assign c[105:104] = a[157:156];
    assign c[107:106] = 0;
    assign c[109:108] = 0;
    assign c[111:110] = a[159:158];
    assign c[113:112] = 0;
    assign c[115:114] = 0;
    assign c[117:116] = a[169:168];
    assign c[119:118] = 0;
    assign c[121:120] = 0;
    assign c[123:122] = a[155:154];
    assign c[125:124] = 0;
    assign c[127:126] = 0;
    assign c[129:128] = a[173:172];
    assign c[131:130] = 0;
    assign c[133:132] = 0;
    assign c[135:134] = a[175:174];
    assign c[137:136] = 0;
    assign c[139:138] = 0;
    assign c[141:140] = a[169:168];
    assign c[143:142] = 0;
    assign c[145:144] = 0;
    assign c[147:146] = a[163:162];
    assign c[149:148] = 0;
    assign c[151:150] = 0;
    assign c[153:152] = a[173:172];
    assign c[155:154] = 0;
    assign c[157:156] = 0;
    assign c[159:158] = a[175:174];
    assign c[161:160] = 0;
    assign c[163:162] = 0;
    assign c[165:164] = a[185:184];
    assign c[167:166] = 0;
    assign c[169:168] = 0;
    assign c[171:170] = a[171:170];
    assign c[173:172] = 0;
    assign c[175:174] = 0;
    assign c[177:176] = a[189:188];
    assign c[179:178] = 0;
    assign c[181:180] = 0;
    assign c[183:182] = a[191:190];
    assign c[185:184] = 0;
    assign c[187:186] = 0;
    assign c[189:188] = a[185:184];
    assign c[191:190] = 0;
    assign c[193:192] = 0;
endmodule
