// sdram.v

// Generated using ACDS version 13.0 156 at 2013.08.15.18:11:30

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,                //        clk.clk
		input  wire        reset_reset_n,          //      reset.reset_n
		input  wire [24:0] sdram_s1_address,       //   sdram_s1.address
		input  wire [3:0]  sdram_s1_byteenable_n,  //           .byteenable_n
		input  wire        sdram_s1_chipselect,    //           .chipselect
		input  wire [31:0] sdram_s1_writedata,     //           .writedata
		input  wire        sdram_s1_read_n,        //           .read_n
		input  wire        sdram_s1_write_n,       //           .write_n
		output wire [31:0] sdram_s1_readdata,      //           .readdata
		output wire        sdram_s1_readdatavalid, //           .readdatavalid
		output wire        sdram_s1_waitrequest,   //           .waitrequest
		output wire [12:0] sdram_wire_addr,        // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //           .ba
		output wire        sdram_wire_cas_n,       //           .cas_n
		output wire        sdram_wire_cke,         //           .cke
		output wire        sdram_wire_cs_n,        //           .cs_n
		inout  wire [31:0] sdram_wire_dq,          //           .dq
		output wire [3:0]  sdram_wire_dqm,         //           .dqm
		output wire        sdram_wire_ras_n,       //           .ras_n
		output wire        sdram_wire_we_n,        //           .we_n
		output wire        sdram_clk_clk           //  sdram_clk.clk
	);

	wire    up_clocks_0_sys_clk_clk;            // up_clocks_0:sys_clk -> [rst_controller:clk, sdram_controller:clk]
	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> sdram_controller:reset_n
	wire    rst_controller_001_reset_out_reset; // rst_controller_001:reset_out -> up_clocks_0:reset

	sdram_sdram_controller sdram_controller (
		.clk            (up_clocks_0_sys_clk_clk),         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset), // reset.reset_n
		.az_addr        (sdram_s1_address),                //    s1.address
		.az_be_n        (sdram_s1_byteenable_n),           //      .byteenable_n
		.az_cs          (sdram_s1_chipselect),             //      .chipselect
		.az_data        (sdram_s1_writedata),              //      .writedata
		.az_rd_n        (sdram_s1_read_n),                 //      .read_n
		.az_wr_n        (sdram_s1_write_n),                //      .write_n
		.za_data        (sdram_s1_readdata),               //      .readdata
		.za_valid       (sdram_s1_readdatavalid),          //      .readdatavalid
		.za_waitrequest (sdram_s1_waitrequest),            //      .waitrequest
		.zs_addr        (sdram_wire_addr),                 //  wire.export
		.zs_ba          (sdram_wire_ba),                   //      .export
		.zs_cas_n       (sdram_wire_cas_n),                //      .export
		.zs_cke         (sdram_wire_cke),                  //      .export
		.zs_cs_n        (sdram_wire_cs_n),                 //      .export
		.zs_dq          (sdram_wire_dq),                   //      .export
		.zs_dqm         (sdram_wire_dqm),                  //      .export
		.zs_ras_n       (sdram_wire_ras_n),                //      .export
		.zs_we_n        (sdram_wire_we_n)                  //      .export
	);

	sdram_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (up_clocks_0_sys_clk_clk),            //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk)                       //            sdram_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (up_clocks_0_sys_clk_clk),        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

endmodule
