//Jul.5.2004 reduce critical path cell

`include "define.h"
module 
shifter(a,c,shift_func,shift_amount);
	input [31:0] a;
	output [31:0] c;
	input [1:0] shift_func;
	input [4:0] shift_amount;

	 reg [31:0] c=0;




endmodule