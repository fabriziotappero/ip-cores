-- Testbench for Filters H_a1-4(z)
-- Uses a sine sweep as stimuli
-- 
-- This program is free software; you can redistribute it and/or modify it under the terms of the GNU General Public License
-- as published by the Free Software Foundation; either version 3 of the License, or (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License along with this program; 
-- if not, see <http://www.gnu.org/licenses/>.


library ieee;
library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;
use ieee.math_real.all;

use work.analytic_filter_h_a1_pkg.all;
use work.analytic_filter_h_a2_pkg.all;
use work.analytic_filter_h_a3_pkg.all;
use work.analytic_filter_h_a4_pkg.all;

entity analytic_filter_tb is
	generic(
		clk_period : time := 10 ns;
		input_data_width : integer := 16;
		output_data_width : integer := 16;
		filter_delay_in_clks : integer  := 7; --delay of hilbert filter
    data_width : integer := 16
	);
end analytic_filter_tb; 

architecture analytic_filter_tb_arch of analytic_filter_tb is
  signal x : std_logic_vector(input_data_width-1 downto 0) := (others => '0'); --input
  signal i,q : std_logic_vector(output_data_width-1 downto 0); --output
  signal i_real,q_real : real;
  signal x_real : real;
  signal anal_data_i : std_logic_vector(input_data_width-1 downto 0);
  signal clk : std_logic := '0';
  signal rst : std_logic;

  type filter_in_table is array (0 to 1034) of std_logic_vector(15 downto 0);

  -- sine sweep
  constant filter_in_force : filter_in_table :=
    (
     to_stdlogicvector(bit_vector'(X"7FFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FF7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FE9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FD0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FA7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F68"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F0D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E8E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7DE2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D02"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7BE2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A79"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"78BC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"769F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7416"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7116"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6D93"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6981"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"64D6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5F87"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"598B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"52DB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4B71"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"434B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3A68"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"30CA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2679"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1B7F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0FEC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"03D4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F751"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EA82"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DD8B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D098"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C3D9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B781"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ABCC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A0F5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"973D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8EE4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"882C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8353"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8092"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"801E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8220"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"86B8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8DF5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"97D9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A450"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B334"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C445"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D731"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EB8D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"00D7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"167D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2BDA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"403C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"52ED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6336"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7067"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"79DF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F16"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FA5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7B4F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7205"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"63F1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5174"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3B2D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"21F3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"06D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EAFC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CFCB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B6A3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A0E5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FDB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"84A1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8012"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"82B3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8CA2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9D8D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B4AC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D0C5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F038"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1110"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3124"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4E36"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6620"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"76FA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F4A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E28"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7359"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5F67"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"43A0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"220B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FD49"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D863"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B68F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9AE7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"881B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"802D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"842D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9413"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AEA8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D193"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F985"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"227F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4837"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6687"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"79ED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FF5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7793"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"615E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3F93"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"15ED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E947"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BF10"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9CA4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8699"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"801A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8A66"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A483"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CB45"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F99D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2936"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"534A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"719F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F76"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A5D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"62AB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3B9C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0AF3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D835"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AB83"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8C4E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8010"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8940"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A6C3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D3EA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"091C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3D09"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"664B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D1B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7CDD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6523"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"39FC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"035B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CBBA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9E1D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"83E4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"82C7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9B7C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C958"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"030C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3C71"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"690F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EDA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"788B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"570B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"217E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E3E8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AC88"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8896"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8107"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"982E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C8E8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0791"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"44AB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"70AC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E20"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3F3F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FF51"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BF3C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"906C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8006"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9319"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C4DB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"07A9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"489A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"74CD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EF5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6387"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2A25"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E3B9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A59D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8327"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8789"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B1F6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F579"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3CB1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"707C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F8A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"644F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2751"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DCBA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9DDF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80A3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FB4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C665"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"11D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5729"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D35"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7596"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"427D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F660"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AD91"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"83C7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8977"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BD0F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0B04"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"54F3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D62"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"73A5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3B06"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EA0E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A1D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"807A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9488"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D62B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"29ED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6BF0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F4B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5AED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0E39"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BAE5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8655"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"88C0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C1B6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"179A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"62D5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"60C0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1349"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BC47"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85C6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8AC6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C981"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"237F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6C0A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E59"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5081"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F944"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A536"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"801F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9DF7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EFB7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4A67"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D75"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6CD6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"20DC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C29A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8602"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8D36"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D4E4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"352D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7775"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"755D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2F64"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CD99"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8916"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8AA8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D217"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3543"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7890"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"72BA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2699"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C26F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"843C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"934A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E6E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4AA2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F00"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"61D2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0536"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A4F2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8033"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AFD4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"14EF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6C4A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7AD7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3607"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CC1A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"859C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"93B2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ED52"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5449"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"50D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E7B4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FD3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8906"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D8FC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"45C8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F4C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5A53"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F1B3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9396"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"875D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D710"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4658"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F9B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"55EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E908"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8DEF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8CD3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E756"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"55CB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F6C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"41EF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CE96"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"837D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9EE4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0AE5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E0B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"750F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1948"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A7D8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8172"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C7A9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3EB0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F80"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"510B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DB47"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85BA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9CAA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0C6D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"713E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6FEB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"08E1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9987"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"881F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E571"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5B9D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C6F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2872"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AE1B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"814B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CD58"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4A26"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FA4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"396C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BB15"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8014"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C308"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4281"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FF9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3D6F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BCF6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8014"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C529"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"467D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FA1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3515"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B354"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8155"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D40C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5535"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C58"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1F36"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A08C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8849"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F14F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6A71"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6FA4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FA75"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8B33"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9D15"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1D08"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7CB8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5075"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C953"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C86D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5095"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C3B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"185B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"980F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"90DB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0BEE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"791F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5727"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CD8B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8001"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CBEB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"56B3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"78B1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"07F0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8D58"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9F50"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2883"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FB5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3825"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AA56"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"87E1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FCD2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"75EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"592F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CA78"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8047"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DA9B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6570"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6C8E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E5F2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"815A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C370"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"55B2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7649"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F920"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"850B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B641"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4B25"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A3E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"02DA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8770"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B187"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"47E9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7AD4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"02F3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"86D6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B487"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4C8A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7879"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F96B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"83A2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BFBB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"583C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7193"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E66D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"805A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D490"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6885"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"62C8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CB18"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"81C2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F458"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7872"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"47E5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AAFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8E89"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1E51"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1DEF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8DD4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ADA0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4CEA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"74D8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E69F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8006"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E264"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7383"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4DE9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AC86"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9022"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"26BF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F38"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0AA8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"84C9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C6ED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6620"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5E5E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BBB1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8978"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1B35"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FE0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0FA4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8536"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C8A7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6948"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"582A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B19A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9051"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2DA6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7CDD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F580"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8031"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E808"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"798A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"374F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9458"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AE34"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5814"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"666D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BF3C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8B2B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"278F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D2C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F1F6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8002"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F579"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E12"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2138"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"87AE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CA8F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6FB2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"46E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9AE9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AA8E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5952"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6140"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B2EA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"957C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"40F7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"718C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CA99"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8951"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2ABE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A48"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DEC7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8351"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1905"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E31"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EDC5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0CED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F8A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F6DD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"803D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"06E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FD8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F9D9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8029"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"06F8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FC1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F6AD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"807B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0D35"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F08"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ED65"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"81E1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"197B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C91"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DE3B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85E6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2B5D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"766B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C9EA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8ED4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"41B2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6A04"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B229"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9F65"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5A10"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"54A3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9A38"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BA1C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"704A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3448"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"873C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E01A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E4E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0912"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8009"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0F96"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7CD4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D6E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8BDF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4244"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6557"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A699"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AFAA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6CB1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3584"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85D7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EA13"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FE8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F357"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"83A5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2FC1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E8A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AFC0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A999"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6AA8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3515"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8484"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F2F0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FBB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E22C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8A87"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"46A6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5C6E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"982B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C98F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7BFD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"07A5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8128"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"29B4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E4D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AA1E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B4B2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"74E5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1A57"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8001"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1CBE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7360"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B049"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B067"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"73C5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1A58"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"800E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"21F8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6FA5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A825"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BB61"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"79BA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"07A8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"827E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"389D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6017"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"951D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D895"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FE5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E231"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9084"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5B64"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3C5B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"82A4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0B25"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"76D5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AFC5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B863"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A9D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FE23"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"86A1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4BEA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4A80"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85DA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0232"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"78A3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B0C1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BA8E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C4F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F3DB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8BDB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"599D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"37BB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80AD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1F6F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6981"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"973D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E00E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F38"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C54C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AB12"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7814"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FD49"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8A0F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5A05"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"32A8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8007"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2E47"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5C87"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8AB6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FE54"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7671"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A4BA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D1D7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FE3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C7A1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ADC3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7B18"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ED78"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9454"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6BBC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"11A8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8598"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"55D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3140"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8028"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3CF1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4AD6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"81E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"23F7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5E2F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"886B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0CD6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6BDC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"91A0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F8BB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"74DB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9BB0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E834"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A50"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A536"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DB63"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D51"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AD34"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D22E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EC8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B2FF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CC64"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F62"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B630"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C9D8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F88"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B696"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CA75"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F5D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B429"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CE3E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EBA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AF10"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D555"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D33"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A7A1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DFEC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A16"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9E73"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EE2C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7478"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"946A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"001F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6B3F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8ACE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"157E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5D49"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8350"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2D85"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"499B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8004"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"46BC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2FAE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8339"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5ED9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0FC9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8F2F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"72B0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EB6B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A58F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E6D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C59B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C6CA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7E15"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A306"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F14F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E65"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"89AE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"20F4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4E0A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4EC6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1EF0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8B44"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"71A3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E742"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AD7F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FF8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B180"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E35A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7293"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8B02"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"22E5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"480A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80AB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5C45"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"07A8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9A08"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D32"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C20E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D464"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"772F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8E15"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2019"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"46EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"815B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"62CB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F99C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A616"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AC27"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F287"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6601"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"81BE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"47BF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1B05"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"931B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7C13"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BFF8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DDA4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6FF0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"851A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3D78"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"23B5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9022"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7B5C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BFB9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E0E4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6CAC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"82C8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4837"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1468"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9A6C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F5E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AB83"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FC99"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5935"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8038"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6382"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EC3B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BA22"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7B91"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8D72"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3010"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2A25"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"90C9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D89"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B13A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FA2E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5754"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80E2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6AF2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DB11"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CE14"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"718C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"82BF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5063"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"004A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AF76"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D0E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8D27"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3703"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1C2F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9CEB"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FF5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"98B7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"23F4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2DDE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"934A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F7E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A0B9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"197B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3607"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FCA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EF3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A2CF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1858"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3555"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"911C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F75"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9E73"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"209A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2BB7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"97C4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"94C8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"31B9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"186F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A5FA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D4D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"88F4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"49EA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FAED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BEED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7243"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80A2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"64DC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D485"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E527"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"58C2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8411"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7A6D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AAC2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"17A9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2C5D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9C79"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EA2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"895A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4E51"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EEF4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CF8D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"64D2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8166"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7795"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ADE6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1820"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"278D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A2DD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7BC1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8390"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5F8A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D3A2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EF30"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"49C9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8E46"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FFF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8E15"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4B11"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EBBA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D97E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"58D8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"878B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F38"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"93C3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"43CA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F1BF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D64A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5955"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"883E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FA7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FFE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4C25"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E51D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E536"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4B71"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"912D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F38"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"85B6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"614C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C747"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0762"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2AC5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AA10"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"73AE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"802E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"78F4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9F7E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3A65"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F3AE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DCE2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4D63"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9319"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7DBF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"81F1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6E35"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AF6B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2933"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"02E3"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D1BD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"53D2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"90A4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7DFE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8197"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"70F0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A899"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"34D4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F2EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E456"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4142"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9FE9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"755D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80AC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7D61"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FF6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"58D4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C5EE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"16A5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0E55"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"CE3E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"50D0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"96D4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7928"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"802F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7CF5"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8EE9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5D5A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BCA0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2524"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FB36"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"E481"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"39AD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AC0C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"68E0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8899"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7EED"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"80B8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"78B7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9429"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"5992"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BCF6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2987"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F19F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F2F0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"278A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C016"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"553A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"9949"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"73D4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"83C2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7FD8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8148"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"791F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"908B"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"6240"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ADE6"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3FAC"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D45A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"16B4"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"FE83"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"EC9E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"275F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C5FF"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4AE2"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A64C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"663C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8FAD"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"77E8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"8307"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7F94"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"802D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7DDE"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"861D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"7417"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"934E"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"63F1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"A5F0"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4F48"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"BC2C"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"37E8"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"D448"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1F6F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"ECCA"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0732"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0481"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"F038"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"1A8F"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"DB3A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"2E61"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"C8A7"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"3FA9"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"B8B1"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"4E4D"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"AB5A"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0),
     to_stdlogicvector(bit_vector'(X"0000"))(15 DOWNTO 0));

begin
    analytic_filter_inst : analytic_filter_h_a4 --change this to analytic_filter_h_ax to test other filters
    generic map(
--      input_data_width  => input_data_width,  --uncomment this for analytic_filter_h_a1
--      output_data_width => output_data_width, --uncomment this for analytic_filter_h_a1
--			filter_delay_in_clks => filter_delay_in_clks --uncomment this for analytic_filter_h_a1
      data_width => data_width --uncomment this for analytic_filter_h_a3-4
    )
    port map(
      rst_i           => rst,
      clk_i           => clk,
	    data_str_i 	=> '1',
	    data_i 			=> anal_data_i,
	    data_i_o 		=> i,
	    data_q_o 		=> q,
	    data_str_o 	=> open
    );
    
    clk <= not clk after clk_period/2;
    rst <= '1', '0' after 20 ns;

    --choose scaling, not all filters have the full dynamic range
    anal_data_i <= x;
--    anal_data_i <= std_logic_vector(shift_right(signed(x),1));
--    anal_data_i <= std_logic_vector(shift_right(signed(x),2));

    x_real <= real(to_integer(signed(x)))/ 2.0**(input_data_width-1);
    i_real <= real(to_integer(signed(i)))/ 2.0**(output_data_width-1);
    q_real <= real(to_integer(signed(q)))/ 2.0**(output_data_width-1);
    
  --choose imput stimuli:
--    x <= x"7FFF", x"0000" after 40 ns; --impulse response
--    x <= x"7FFF"; --step response

  filter_in_gen: process
  begin
    x <= filter_in_force(0);
    wait for clk_period*3;
    x <= filter_in_force(1);
    wait for clk_period;
    for n in 0 to 1034 loop
      if n + 2 <= 1034 then
        x <= filter_in_force(n + 2);
      end if;
      wait for clk_period;
    end loop;
    assert false report "**** test complete. ****" severity note;
  end process filter_in_gen;

end analytic_filter_tb_arch;