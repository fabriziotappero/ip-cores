-------------------------------------------------------------------------------
--
-- T8243 Core
--
-- $Id: t8243_core-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-------------------------------------------------------------------------------

configuration t8243_core_rtl_c0 of t8243_core is

  for rtl
  end for;

end t8243_core_rtl_c0;
