--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:            15:34, 2001.04.22. *
--* Tested entity name:                         wb_bus_dnsize *
--* File name contains tested entity: $DSN\src\wb_bus_dnsize.vhd *
--*************************************************************

library ieee,wb_tk,synopsys;
use ieee.std_logic_1164.all;
use wb_tk.technology.all;
use synopsys.std_logic_arith.all;
use wb_tk.wb_test.all;

entity wb_bus_dnsize_tb is
	generic(
		m_bus_width : POSITIVE := 64;
		m_addr_width : POSITIVE := 6;
		s_bus_width : POSITIVE := 16;
		s_addr_width : POSITIVE := 8;
		little_endien : BOOLEAN := true );
end wb_bus_dnsize_tb;

architecture TB of wb_bus_dnsize_tb is
	component wb_bus_dnsize
	generic(
		m_bus_width : POSITIVE := m_bus_width;
		m_addr_width : POSITIVE := m_addr_width;
		s_bus_width : POSITIVE := s_bus_width;
		s_addr_width : POSITIVE := s_addr_width;
		little_endien : BOOLEAN := little_endien
	);
	port(
		m_adr_i : in std_logic_vector((m_addr_width-1) downto 0);
		m_sel_i : in std_logic_vector(((m_bus_width/8)-1) downto 0);
		m_dat_i : in std_logic_vector((m_bus_width-1) downto 0);
		m_dat_oi : in std_logic_vector((m_bus_width-1) downto 0);
		m_dat_o : out std_logic_vector((m_bus_width-1) downto 0);
		m_cyc_i : in std_logic;
		m_ack_o : out std_logic;
		m_ack_oi : in std_logic;
		m_err_o : out std_logic;
		m_err_oi : in std_logic;
		m_rty_o : out std_logic;
		m_rty_oi : in std_logic;
		m_we_i : in std_logic;
		m_stb_i : in std_logic;
		s_adr_o : out std_logic_vector((s_addr_width-1) downto 0);
		s_sel_o : out std_logic_vector(((s_bus_width/8)-1) downto 0);
		s_dat_i : in std_logic_vector((s_bus_width-1) downto 0);
		s_dat_o : out std_logic_vector((s_bus_width-1) downto 0);
		s_cyc_o : out std_logic;
		s_ack_i : in std_logic;
		s_err_i : in std_logic;
		s_rty_i : in std_logic;
		s_we_o : out std_logic;
		s_stb_o : out std_logic
	);
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal m_adr_i : std_logic_vector((m_addr_width-1) downto 0);
	signal m_sel_i : std_logic_vector(((m_bus_width/8)-1) downto 0) := (others => '0');
	signal m_dat_i : std_logic_vector((m_bus_width-1) downto 0);
	signal m_dat_oi : std_logic_vector((m_bus_width-1) downto 0) := (others => 'U');
	signal m_cyc_i : std_logic;
	signal m_ack_oi : std_logic := 'U';
	signal m_err_oi : std_logic := 'U';
	signal m_rty_oi : std_logic := 'U';
	signal m_we_i : std_logic;
	signal m_stb_i : std_logic;
	signal s_dat_i : std_logic_vector((s_bus_width-1) downto 0);
	signal s_ack_i : std_logic;
	signal s_err_i : std_logic;
	signal s_rty_i : std_logic;
	-- Observed signals - signals mapped to the output ports of tested entity
	signal m_dat_o : std_logic_vector((m_bus_width-1) downto 0);
	signal m_ack_o : std_logic;
	signal m_err_o : std_logic;
	signal m_rty_o : std_logic;
	signal s_adr_o : std_logic_vector((s_addr_width-1) downto 0);
	signal s_sel_o : std_logic_vector(((s_bus_width/8)-1) downto 0);
	signal s_dat_o : std_logic_vector((s_bus_width-1) downto 0);
	signal s_cyc_o : std_logic;
	signal s_we_o : std_logic;
	signal s_stb_o : std_logic;

	signal clk_i: std_logic;
	signal rst_i: std_logic;
begin

	-- Unit Under Test port map
	UUT : wb_bus_dnsize
		port map
			(m_adr_i => m_adr_i,
			m_sel_i => m_sel_i,
			m_dat_i => m_dat_i,
			m_dat_oi => m_dat_oi,
			m_dat_o => m_dat_o,
			m_cyc_i => m_cyc_i,
			m_ack_o => m_ack_o,
			m_ack_oi => m_ack_oi,
			m_err_o => m_err_o,
			m_err_oi => m_err_oi,
			m_rty_o => m_rty_o,
			m_rty_oi => m_rty_oi,
			m_we_i => m_we_i,
			m_stb_i => m_stb_i,
			s_adr_o => s_adr_o,
			s_sel_o => s_sel_o,
			s_dat_i => s_dat_i,
			s_dat_o => s_dat_o,
			s_cyc_o => s_cyc_o,
			s_ack_i => s_ack_i,
			s_err_i => s_err_i,
			s_rty_i => s_rty_i,
			s_we_o => s_we_o,
			s_stb_o => s_stb_o );

	clk: process is
	begin
		clk_i <= '0';
		wait for 25ns;
		clk_i <= '1';
		wait for 25ns;
	end process;
	
	reset: process is
	begin
		rst_i <= '1';
		wait for 150ns;
		rst_i <= '0';
		wait;
	end process;
	
	master: process is
	begin
		m_we_i <= '0';
		m_cyc_i <= '0';
		m_stb_i <= '0';
		m_adr_i <= (others => '0');
		m_dat_i <= (others => '0');
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';
		wait until clk_i'EVENT and clk_i = '1';

		wr_val(clk_i, m_adr_i,m_dat_o,m_dat_i,m_we_i,m_cyc_i,m_stb_i,m_ack_o,"000101","1111111011011100101110101001100001110110010101000011001000010000");
		rd_val(clk_i, m_adr_i,m_dat_o,m_dat_i,m_we_i,m_cyc_i,m_stb_i,m_ack_o,"000101","1111111011011100101110101001100001110110010101000011001000010000");
--		wr_val(clk_i, m_adr_i,m_dat_o,m_dat_i,m_we_i,m_cyc_i,m_stb_i,m_ack_o,"000101","01110110010101000011001000010000");
--		rd_val(clk_i, m_adr_i,m_dat_o,m_dat_i,m_we_i,m_cyc_i,m_stb_i,m_ack_o,"000101","01110110010101000011001000010000");

		m_sel_i <= add_one(m_sel_i);
--		if (sel_i = "1111") then wait; end if;
	end process;

	s_ack_i <= s_stb_o;
	s_dat_i <= (others => '1');
	s_err_i <= '0';
	s_rty_i <= '0';
end TB;

configuration TB_wb_bus_dnsize of wb_bus_dnsize_tb is
	for TB
		for UUT : wb_bus_dnsize
			use entity work.wb_bus_dnsize(wb_bus_dnsize);
		end for;
	end for;
end TB_wb_bus_dnsize;

