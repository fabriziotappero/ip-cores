-------------------------------------------------------------------------------------------------100
--| Modular Oscilloscope
--| UNSL - Argentine
--|
--| File: eppwbn_16bit_test_tbench_text.vhd
--| Version: 0.01
--| Tested in: Actel APA300
--|-------------------------------------------------------------------------------------------------
--| Description:
--|   EPP - Wishbone bridge. 
--|   This file is only for test purposes. Testing eppwbn 16 bit. Test bench.
--|   It may not work for other than Actel Libero software.
--|-------------------------------------------------------------------------------------------------
--| File history:
--|   0.01  | mar-2009 | First release
----------------------------------------------------------------------------------------------------
--| Copyright � 2009, Facundo Aguilera.
--|
--| This VHDL design file is an open design; you can redistribute it and/or
--| modify it and/or implement it after contacting the author.
----------------------------------------------------------------------------------------------------


-- NOTE:  It may not work for other than Actel Libero software.
--        You can download Libero for free from Actel website.





-- Generated by WaveFormer Lite Version 12.30a at 12:26:42 on 3/13/2009
-- Stimulator for stimulus

-- Generation Settings:
--   Export type: Stimulus only (reactive export not enabled)
--                Delays, Samples, Markers, etc will not generate code.

-- Clock Domains:

--   Unclocked
--   ---------
--     Signals:
--       rst
--       nSelectIn
--       Data
--       nAutoFd
--       nStrobe
--       nInit

library ieee, std;
use ieee.std_logic_1164.all;
library syncad_vhdl_lib;
use syncad_vhdl_lib.TBDefinitions.all;
-- Additional libraries used by Model Under Test.
library IEEE;
use work.eppwbn_pgk.all;
-- End Additional libraries used by Model Under Test.

entity stimulus is
  port (
    clk : inout std_logic := '0';
    rst : inout std_logic := '0';
    nSelectIn : inout std_logic := '0';
    Data : inout std_logic_vector(7 downto 0) := "00000000";
    nAutoFd : inout std_logic := '1';
    nStrobe : inout std_logic := '0';
    nInit : inout std_logic := '1');

end stimulus;

architecture STIMULATOR of stimulus is

  -- Control Signal Declarations
  signal tb_status : TStatus;
  signal tb_ParameterInitFlag : boolean := false;

  -- Parm Declarations
  signal clk_MinHL : time := 0 ns;
  signal clk_MaxHL : time := 0 ns;
  signal clk_MinLH : time := 0 ns;
  signal clk_MaxLH : time := 0 ns;
  signal clk_JFall : time := 0 ns;
  signal clk_JRise : time := 0 ns;
  signal clk_Duty : real := 0.0;
  signal clk_Period : time := 0 ns;
  signal clk_Offset : time := 0 ns;

  -- Status Control block.

begin

  process
    variable good : boolean;
  begin
    wait until tb_ParameterInitFlag;
    tb_status <= TB_ONCE;
    wait for 360000 ns;
    tb_status <= TB_DONE;
    wait;
  end process;

  -- Parm Assignment Block
  AssignParms : process
    variable clk_MinHL_real : real;
    variable clk_MaxHL_real : real;
    variable clk_MinLH_real : real;
    variable clk_MaxLH_real : real;
    variable clk_JFall_real : real;
    variable clk_JRise_real : real;
    variable clk_Duty_real : real;
    variable clk_Period_real : real;
    variable clk_Offset_real : real;
  begin
    clk_MinHL_real := 0.0;
    clk_MinHL <= clk_MinHL_real * 1 ns;
    clk_MaxHL_real := 0.0;
    clk_MaxHL <= clk_MaxHL_real * 1 ns;
    clk_MinLH_real := 0.0;
    clk_MinLH <= clk_MinLH_real * 1 ns;
    clk_MaxLH_real := 0.0;
    clk_MaxLH <= clk_MaxLH_real * 1 ns;
    clk_JFall_real := 0.0;
    clk_JFall <= clk_JFall_real * 1 ns;
    clk_JRise_real := 0.0;
    clk_JRise <= clk_JRise_real * 1 ns;
    clk_Duty_real := 50.0;
    clk_Duty <= clk_Duty_real;
    clk_Period_real := 100.0;
    clk_Period <= clk_Period_real * 1 ns;
    clk_Offset_real := 0.0;
    clk_Offset <= clk_Offset_real * 1 ns;
    tb_ParameterInitFlag <= true;
    wait;
  end process;

  -- Clocks

  -- Clock Instantiation
  tb_clk : entity syncad_vhdl_lib.tb_clock_minmax
    generic map (name => "tb_clk",
                initialize => true,
                state1 => '1',
                state2 => '0')
    port map (tb_status,
              clk,
              clk_MinLH,
              clk_MaxLH,
              clk_MinHL,
              clk_MaxHL,
              clk_Offset,
              clk_Period,
              clk_Duty,
              clk_JRise,
              clk_JFall);

  -- Clocked Sequences

  -- Sequence: Unclocked
  Unclocked : process
  begin
    -- Initial Reset
    wait for 700 ns;
    rst <= '1';
    wait for 800 ns;
    rst <= '0';
    
    
    -------------------- Test Negotiation
    -- Negotiation
    --  st0
    wait for 800 ns;
    Data <= x"40";
    nStrobe <= '1';
    --  st1
    wait for 800 ns;
    nSelectIn <= '1';
    nAutoFd <= '0';
    --  st3
    wait for 800 ns;
    nStrobe <= '0';
    --  st4
    wait for 800 ns;
    nAutoFd <= '1';
    nStrobe <= '1';
    
    -------------------- Test write add 0x10 data 0x1234
    -- Add WR
    wait for 800 ns;
    Data <= x"10";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 800 ns;
    Data <= x"12";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 800 ns;
    Data <= x"34";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -------------------- Test write add 0x55 data 0x4321
    -- Add WR
    wait for 800 ns;
    Data <= x"55";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';

    -- Data WR
    wait for 800 ns;
    Data <= x"43";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 400 ns;
    Data <= x"21";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -------------------- Test write add changed (fist 56 then 57) data 0x1122
    -- Add WR
    wait for 800 ns;
    Data <= x"56";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';

    -- Data WR
    wait for 800 ns;
    Data <= x"33";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Add WR
    wait for 800 ns;
    Data <= x"57";
    nSelectIn <= '0';
    nStrobe <= '0';
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 800 ns;
    Data <= x"11";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 800 ns;
    Data <= x"22";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -------------------- Test write add 0x58 data 0x99 with timeout
    wait for 800 ns;
    Data <= x"58";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
   
    -- Data WR
    wait for 800 ns;
    Data <= x"99";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
   
    wait for 120000 ns;
    
   -------------------- Test write add 0x59 data 0x5678
    -- Add WR
    wait for 800 ns;
    Data <= x"59";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';

    -- Data WR
    wait for 800 ns;
    Data <= x"56";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data WR
    wait for 800 ns;
    Data <= x"78";    -- DATA
    nAutoFd <= '0';   -- DataSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nAutoFd <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -------------------- Test add read (it must be 0x59)
    -- Adr RE
    wait for 800 ns;
    Data <= "ZZZZZZZZ";   -- DATA ('Z...')
    wait for 800 ns;      
    nSelectIn <= '0';       -- DataSTB
    wait for 800 ns;
    nSelectIn <= '1';
    
    
    -------------------- Test data read add 0x10 (it must be 0x1234)
    -- Add WR
    wait for 800 ns;
    Data <= x"10";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    nAutoFd <= '0';    -- DataSTB
    wait for 200 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 200 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    nAutoFd <= '0';    -- DataSTB
    wait for 400 ns;
    nAutoFd <= '1';
    
    -------------------- Test data read add 0x55 (it must be 0x4321)
    -- Add WR
    wait for 800 ns;
    Data <= x"55";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    

    -------------------- Test data read add 0x56 (it must be 0x0000)
    -- Add WR
    wait for 800 ns;
    Data <= x"56";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -------------------- Test data read add 0x57 (it must be 0x1122)
    -- Add WR
    wait for 800 ns;
    Data <= x"57";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -------------------- Test data read add 0x57 (it must be 0x1122)
    -- Add WR
    wait for 800 ns;
    Data <= x"57";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';    
    
    -------------------- Test data read add 0x58 (it must be 0x0000)
    -- Add WR
    wait for 800 ns;
    Data <= x"58";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';    
    
    -------------------- Test data read add 0x59 (it must be 0x5678)
    -- Add WR
    wait for 800 ns;
    Data <= x"59";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';    
    
    -------------------- Test data read add 0x55 then 0x10 (it must be 0x1234)
    -- Add WR
    wait for 800 ns;
    Data <= x"55";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Add WR
    wait for 800 ns;
    Data <= x"10";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 1600 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';   
    
    -------------------- Test data read add 0x55 with timeout then 0x59 (it must be 0x5678)
    -- Add WR
    wait for 800 ns;
    Data <= x"55";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    wait for 120000 ns;
    
    -- Add WR
    wait for 800 ns;
    Data <= x"59";    -- DATA
    nSelectIn <= '0'; -- AddSTB
    nStrobe <= '0';   -- WR
    wait for 800 ns;
    nSelectIn <= '1';
    wait for 800 ns;
    nStrobe <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';
    
    -- Data RE
    wait for 400 ns;
    Data <= "ZZZZZZZZ";-- DATA ('Z...')
    wait for 800 ns;      
    nAutoFd <= '0';    -- DataSTB
    wait for 800 ns;
    nAutoFd <= '1';   
   
    
    wait;
  end process;
end STIMULATOR;

-- Test Bench wrapper for stimulus and Model Under Test
library ieee, std;
use ieee.std_logic_1164.all;
library syncad_vhdl_lib;
use syncad_vhdl_lib.TBDefinitions.all;
-- Additional libraries used by Model Under Test.
library IEEE;
use work.eppwbn_pgk.all;
-- End Additional libraries used by Model Under Test.

entity testbench is
end testbench;
architecture tbGeneratedCode of testbench is
  signal clk : std_logic;
  signal rst : std_logic;
  signal nSelectIn : std_logic;
  signal Data : std_logic_vector(7 downto 0);
  signal nAutoFd : std_logic;
  signal nStrobe : std_logic;
  signal nInit : std_logic;
  signal nAck : std_logic;
  signal busy : std_logic;
  signal PError : std_logic;
  signal Sel : std_logic;
  signal PeriphLogicH : std_logic;
  signal nFault : std_logic;

  -- Stimulator instance

begin

  stimulus_0 : entity work.stimulus
    port map (clk => clk,
              rst => rst,
              nSelectIn => nSelectIn,
              Data => Data,
              nAutoFd => nAutoFd,
              nStrobe => nStrobe,
              nInit => nInit);

  -- Instantiation of Model Under Test.
  eppwbn_16bit_test_0 : entity work.eppwbn_16bit_test
    port map (nStrobe => nStrobe,
              Data => Data,
              nAck => nAck,
              busy => busy,
              PError => PError,
              Sel => Sel,
              nAutoFd => nAutoFd,
              PeriphLogicH => PeriphLogicH,
              nInit => nInit,
              nFault => nFault,
              nSelectIn => nSelectIn,
              rst => rst,
              clk => clk);
end tbGeneratedCode;
