-------------------------------------------------------------------------------
--
-- The decoder unit.
-- Implements the instruction opcodes and controls all units of the T400 core.
--
-- $Id: t400_decoder-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_decoder_rtl_c0 of t400_decoder is

  for rtl
  end for;

end t400_decoder_rtl_c0;
