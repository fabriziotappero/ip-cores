--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Built for project 'SD Bootloader'.
--------------------------------------------------------------------------------
-- This file contains object code in the form of a VHDL byte table constant.
-- This constant can be used to initialize FPGA memories for synthesis or
-- simulation.
-- Note that the object code is stored as a plain byte table in byte address
-- order. This table knows nothing of data endianess and can be used to
-- initialize 32-, 16- or 8-bit-wide memory -- memory initialization functions
-- can be found in package mips_pkg.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.mips_pkg.all;

package obj_code_pkg is

-- Hardcoded simulation parameters ---------------------------------------------

-- Simulation clock rate
constant CLOCK_RATE : integer   := 50e6;
-- Simulation clock period
constant T : time               := (1.0e9/real(CLOCK_RATE)) * 1 ns;

-- Other simulation parameters -------------------------------------------------

constant BRAM_SIZE : integer := 4096;


-- Memory initialization data --------------------------------------------------

constant obj_code : t_obj_code(0 to 14892) := (
  X"10", X"00", X"00", X"7c", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d0", X"82", 
  X"33", X"5a", X"00", X"1f", X"34", X"1b", X"00", X"08", 
  X"13", X"5b", X"00", X"09", X"23", X"7b", X"00", X"01", 
  X"13", X"5b", X"00", X"05", X"23", X"7b", X"00", X"01", 
  X"17", X"5b", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"a3", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"72", X"00", X"00", X"00", X"00", 
  X"40", X"1b", X"70", X"00", X"40", X"1a", X"68", X"00", 
  X"00", X"1a", X"d7", X"c2", X"33", X"5a", X"00", X"01", 
  X"17", X"40", X"00", X"03", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"42", X"00", X"00", X"10", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"fe", X"40", X"84", X"60", X"00", 
  X"0f", X"f0", X"00", X"86", X"00", X"00", X"00", X"00", 
  X"3c", X"04", X"bf", X"c0", X"24", X"84", X"06", X"b8", 
  X"00", X"80", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"05", X"00", X"01", X"40", X"04", X"60", X"00", 
  X"30", X"84", X"ff", X"ff", X"00", X"85", X"28", X"25", 
  X"40", X"85", X"60", X"00", X"3c", X"04", X"00", X"07", 
  X"34", X"84", X"bf", X"fc", X"24", X"06", X"00", X"00", 
  X"24", X"05", X"00", X"ff", X"ac", X"86", X"00", X"00", 
  X"00", X"c5", X"08", X"2a", X"14", X"20", X"ff", X"fd", 
  X"20", X"c6", X"00", X"01", X"24", X"04", X"00", X"00", 
  X"24", X"06", X"00", X"00", X"24", X"05", X"00", X"ff", 
  X"8c", X"80", X"00", X"00", X"20", X"84", X"00", X"10", 
  X"00", X"c5", X"08", X"2a", X"14", X"20", X"ff", X"fc", 
  X"20", X"c6", X"00", X"01", X"3c", X"05", X"00", X"02", 
  X"40", X"04", X"60", X"00", X"30", X"84", X"ff", X"ff", 
  X"00", X"85", X"28", X"25", X"03", X"e0", X"00", X"08", 
  X"40", X"85", X"60", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"3c", X"1b", X"00", X"08", 
  X"27", X"7b", X"c0", X"4c", X"af", X"7d", X"ff", X"f0", 
  X"af", X"7f", X"ff", X"ec", X"af", X"68", X"ff", X"e8", 
  X"af", X"69", X"ff", X"e4", X"af", X"6a", X"ff", X"e0", 
  X"03", X"60", X"e8", X"21", X"40", X"08", X"70", X"00", 
  X"8d", X"1a", X"00", X"00", X"40", X"1b", X"68", X"00", 
  X"07", X"70", X"00", X"2d", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"4e", X"82", X"39", X"28", X"00", X"1f", 
  X"11", X"00", X"00", X"1f", X"39", X"28", X"00", X"1c", 
  X"11", X"00", X"00", X"13", X"00", X"00", X"00", X"00", 
  X"3c", X"08", X"20", X"01", X"ad", X"1a", X"04", X"00", 
  X"8f", X"aa", X"ff", X"e0", X"8f", X"a9", X"ff", X"e4", 
  X"8f", X"a8", X"ff", X"e8", X"8f", X"bf", X"ff", X"ec", 
  X"8f", X"bd", X"ff", X"f0", X"40", X"1b", X"70", X"00", 
  X"40", X"1a", X"68", X"00", X"00", X"1a", X"d7", X"c2", 
  X"33", X"5a", X"00", X"01", X"17", X"40", X"00", X"03", 
  X"23", X"7b", X"00", X"04", X"03", X"60", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"23", X"7b", X"00", X"04", 
  X"03", X"60", X"00", X"08", X"42", X"00", X"00", X"10", 
  X"33", X"5b", X"00", X"3f", X"3b", X"68", X"00", X"20", 
  X"11", X"00", X"00", X"14", X"3b", X"68", X"00", X"21", 
  X"11", X"00", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"3c", X"08", X"20", X"01", X"ad", X"1a", X"04", X"00", 
  X"0b", X"f0", X"00", X"b8", X"00", X"00", X"00", X"00", 
  X"33", X"5b", X"00", X"3f", X"3b", X"68", X"00", X"00", 
  X"11", X"00", X"00", X"1e", X"3b", X"68", X"00", X"04", 
  X"11", X"00", X"00", X"29", X"00", X"00", X"00", X"00", 
  X"3c", X"08", X"20", X"01", X"ad", X"1a", X"04", X"00", 
  X"0b", X"f0", X"00", X"b8", X"00", X"00", X"00", X"00", 
  X"8d", X"1a", X"00", X"04", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"01", X"62", 
  X"3c", X"0a", X"80", X"00", X"00", X"00", X"40", X"21", 
  X"03", X"6a", X"48", X"24", X"15", X"20", X"00", X"03", 
  X"00", X"0a", X"50", X"42", X"15", X"40", X"ff", X"fc", 
  X"25", X"08", X"00", X"01", X"0b", X"f0", X"01", X"18", 
  X"01", X"00", X"d8", X"21", X"0f", X"f0", X"01", X"62", 
  X"3c", X"0a", X"80", X"00", X"00", X"00", X"40", X"21", 
  X"03", X"6a", X"48", X"24", X"11", X"20", X"00", X"03", 
  X"00", X"0a", X"50", X"42", X"15", X"40", X"ff", X"fc", 
  X"25", X"08", X"00", X"01", X"0b", X"f0", X"01", X"18", 
  X"01", X"00", X"d8", X"21", X"0f", X"f0", X"01", X"62", 
  X"00", X"00", X"00", X"00", X"00", X"1a", X"41", X"82", 
  X"31", X"08", X"00", X"1f", X"00", X"1a", X"4a", X"c2", 
  X"31", X"29", X"00", X"1f", X"01", X"09", X"50", X"21", 
  X"00", X"0a", X"50", X"23", X"25", X"4a", X"00", X"1f", 
  X"01", X"5b", X"d8", X"04", X"01", X"5b", X"d8", X"06", 
  X"0b", X"f0", X"01", X"18", X"01", X"1b", X"d8", X"06", 
  X"0f", X"f0", X"01", X"62", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"41", X"82", X"31", X"08", X"00", X"1f", 
  X"00", X"1a", X"4a", X"c2", X"31", X"29", X"00", X"1f", 
  X"01", X"28", X"48", X"23", X"00", X"09", X"58", X"23", 
  X"25", X"6b", X"00", X"1f", X"01", X"1b", X"48", X"04", 
  X"3c", X"0a", X"ff", X"ff", X"35", X"4a", X"ff", X"ff", 
  X"01", X"6a", X"50", X"04", X"01", X"6a", X"50", X"06", 
  X"01", X"0a", X"50", X"04", X"01", X"2a", X"48", X"24", 
  X"01", X"40", X"50", X"27", X"0f", X"f0", X"01", X"62", 
  X"00", X"1a", X"d1", X"40", X"00", X"1a", X"d1", X"42", 
  X"03", X"6a", X"d8", X"24", X"03", X"69", X"d8", X"25", 
  X"0b", X"f0", X"01", X"18", X"00", X"00", X"00", X"00", 
  X"00", X"1a", X"4c", X"02", X"31", X"29", X"00", X"1f", 
  X"3c", X"08", X"bf", X"c0", X"25", X"08", X"04", X"88", 
  X"00", X"09", X"48", X"c0", X"01", X"09", X"40", X"20", 
  X"01", X"00", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"00", X"b8", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"60", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"61", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"62", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"63", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"64", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"65", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"66", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"67", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"af", X"bb", X"ff", X"e8", 
  X"0b", X"f0", X"01", X"20", X"af", X"bb", X"ff", X"e4", 
  X"0b", X"f0", X"01", X"20", X"af", X"bb", X"ff", X"e0", 
  X"0b", X"f0", X"01", X"20", X"37", X"6b", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"6c", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"6d", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"6e", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"6f", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"70", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"71", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"72", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"73", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"74", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"75", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"76", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"77", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"78", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"79", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"7a", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"7b", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"37", X"7c", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"af", X"bb", X"ff", X"ec", 
  X"0b", X"f0", X"01", X"20", X"37", X"7e", X"00", X"00", 
  X"0b", X"f0", X"01", X"20", X"af", X"bb", X"ff", X"f0", 
  X"af", X"bf", X"00", X"00", X"00", X"1a", X"dd", X"42", 
  X"33", X"7b", X"00", X"1f", X"3c", X"08", X"bf", X"c0", 
  X"25", X"08", X"05", X"b8", X"00", X"1b", X"d8", X"c0", 
  X"01", X"1b", X"40", X"20", X"01", X"00", X"f8", X"09", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"1b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"3b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"5b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"7b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"9b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"bb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"db", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"34", X"fb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"8f", X"bb", X"ff", X"e8", 
  X"03", X"e0", X"00", X"08", X"8f", X"bb", X"ff", X"e4", 
  X"03", X"e0", X"00", X"08", X"8f", X"bb", X"ff", X"e0", 
  X"03", X"e0", X"00", X"08", X"35", X"7b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"35", X"9b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"35", X"bb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"35", X"db", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"35", X"fb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"1b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"3b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"5b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"7b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"9b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"bb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"db", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"36", X"fb", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"37", X"1b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"37", X"3b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"37", X"5b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"37", X"7b", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"37", X"9a", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"8f", X"bb", X"ff", X"f0", 
  X"03", X"e0", X"00", X"08", X"37", X"db", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"8f", X"bb", X"ff", X"ec", 
  X"3c", X"1c", X"00", X"08", X"27", X"9c", X"3f", X"ec", 
  X"3c", X"05", X"00", X"08", X"24", X"a5", X"c0", X"00", 
  X"3c", X"04", X"00", X"08", X"24", X"84", X"c0", X"10", 
  X"3c", X"1d", X"00", X"08", X"27", X"bd", X"c4", X"38", 
  X"ac", X"a0", X"00", X"00", X"00", X"a4", X"18", X"2a", 
  X"14", X"60", X"ff", X"fd", X"24", X"a5", X"00", X"04", 
  X"3c", X"04", X"00", X"08", X"24", X"84", X"bf", X"fc", 
  X"3c", X"05", X"bf", X"c0", X"24", X"a5", X"3a", X"2c", 
  X"10", X"a4", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"3c", X"10", X"00", X"00", X"26", X"10", X"00", X"01", 
  X"12", X"00", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"8c", X"a8", X"00", X"00", X"24", X"a5", X"00", X"04", 
  X"ac", X"88", X"00", X"00", X"24", X"84", X"00", X"04", 
  X"1e", X"00", X"ff", X"fb", X"26", X"10", X"ff", X"fc", 
  X"0f", X"f0", X"01", X"f9", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"01", X"cc", X"00", X"00", X"00", X"00", 
  X"27", X"bd", X"ff", X"e8", X"24", X"02", X"00", X"03", 
  X"af", X"bf", X"00", X"14", X"10", X"82", X"00", X"1d", 
  X"00", X"80", X"28", X"21", X"2c", X"82", X"00", X"04", 
  X"10", X"40", X"00", X"0c", X"24", X"02", X"00", X"04", 
  X"24", X"02", X"00", X"01", X"10", X"82", X"00", X"12", 
  X"00", X"00", X"00", X"00", X"3c", X"04", X"bf", X"c0", 
  X"0f", X"f0", X"0d", X"fc", X"24", X"84", X"39", X"50", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"0d", X"fc", 
  X"24", X"84", X"39", X"e0", X"0b", X"f0", X"01", X"df", 
  X"00", X"00", X"00", X"00", X"10", X"82", X"00", X"12", 
  X"24", X"02", X"00", X"0d", X"14", X"82", X"ff", X"f5", 
  X"00", X"00", X"00", X"00", X"3c", X"04", X"bf", X"c0", 
  X"0f", X"f0", X"0d", X"fc", X"24", X"84", X"39", X"20", 
  X"0b", X"f0", X"01", X"dd", X"3c", X"04", X"bf", X"c0", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"0d", X"fc", 
  X"24", X"84", X"39", X"04", X"0b", X"f0", X"01", X"dd", 
  X"3c", X"04", X"bf", X"c0", X"3c", X"04", X"bf", X"c0", 
  X"0f", X"f0", X"0d", X"fc", X"24", X"84", X"38", X"f4", 
  X"0b", X"f0", X"01", X"dd", X"3c", X"04", X"bf", X"c0", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"0d", X"fc", 
  X"24", X"84", X"39", X"40", X"0b", X"f0", X"01", X"dd", 
  X"3c", X"04", X"bf", X"c0", X"3c", X"04", X"bf", X"c0", 
  X"27", X"bd", X"ff", X"c8", X"24", X"84", X"39", X"64", 
  X"af", X"bf", X"00", X"34", X"af", X"b2", X"00", X"24", 
  X"af", X"b5", X"00", X"30", X"af", X"b4", X"00", X"2c", 
  X"af", X"b3", X"00", X"28", X"af", X"b1", X"00", X"20", 
  X"0f", X"f0", X"0d", X"fc", X"af", X"b0", X"00", X"1c", 
  X"3c", X"05", X"00", X"08", X"00", X"00", X"20", X"21", 
  X"0f", X"f0", X"09", X"ff", X"24", X"a5", X"c4", X"50", 
  X"3c", X"12", X"00", X"08", X"3c", X"05", X"bf", X"c0", 
  X"26", X"44", X"c6", X"f4", X"24", X"a5", X"39", X"84", 
  X"0f", X"f0", X"0a", X"10", X"24", X"06", X"00", X"01", 
  X"14", X"40", X"00", X"3a", X"00", X"00", X"00", X"00", 
  X"3c", X"04", X"bf", X"c0", X"3c", X"11", X"00", X"08", 
  X"24", X"84", X"39", X"90", X"26", X"31", X"c6", X"74", 
  X"0f", X"f0", X"0d", X"fc", X"3c", X"13", X"00", X"04", 
  X"00", X"00", X"80", X"21", X"26", X"55", X"c6", X"f4", 
  X"02", X"20", X"a0", X"21", X"26", X"73", X"00", X"01", 
  X"02", X"a0", X"20", X"21", X"02", X"80", X"28", X"21", 
  X"24", X"06", X"00", X"80", X"0f", X"f0", X"0a", X"5e", 
  X"27", X"a7", X"00", X"10", X"14", X"40", X"00", X"25", 
  X"00", X"00", X"00", X"00", X"8f", X"a2", X"00", X"10", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"0d", 
  X"00", X"00", X"10", X"21", X"02", X"22", X"18", X"21", 
  X"90", X"63", X"00", X"00", X"24", X"42", X"00", X"01", 
  X"a2", X"03", X"00", X"00", X"8f", X"a3", X"00", X"10", 
  X"00", X"00", X"00", X"00", X"00", X"43", X"18", X"2b", 
  X"14", X"60", X"ff", X"f8", X"26", X"10", X"00", X"01", 
  X"02", X"13", X"10", X"2b", X"14", X"40", X"ff", X"eb", 
  X"02", X"a0", X"20", X"21", X"0f", X"f0", X"0b", X"18", 
  X"26", X"44", X"c6", X"f4", X"14", X"40", X"00", X"0d", 
  X"00", X"00", X"00", X"00", X"3c", X"04", X"bf", X"c0", 
  X"24", X"84", X"39", X"cc", X"0f", X"f0", X"0d", X"fc", 
  X"02", X"00", X"28", X"21", X"3c", X"04", X"bf", X"c0", 
  X"0f", X"f0", X"0d", X"fc", X"24", X"84", X"39", X"e4", 
  X"00", X"00", X"10", X"21", X"00", X"40", X"f8", X"09", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"02", X"3f", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"01", X"ce", 
  X"00", X"40", X"20", X"21", X"0b", X"f0", X"02", X"36", 
  X"3c", X"04", X"bf", X"c0", X"0f", X"f0", X"01", X"ce", 
  X"00", X"40", X"20", X"21", X"0b", X"f0", X"02", X"31", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"01", X"ce", 
  X"00", X"40", X"20", X"21", X"0b", X"f0", X"02", X"11", 
  X"3c", X"04", X"bf", X"c0", X"03", X"e0", X"00", X"08", 
  X"3c", X"02", X"40", X"21", X"00", X"85", X"28", X"21", 
  X"3c", X"02", X"20", X"00", X"24", X"07", X"ff", X"fb", 
  X"0b", X"f0", X"02", X"b6", X"24", X"06", X"ff", X"fd", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"20", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"11", X"00", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"10", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"11", X"00", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"08", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"11", X"00", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"04", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"11", X"00", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"02", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"11", X"00", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"30", X"63", X"00", X"01", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"02", X"ac", X"48", X"10", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"06", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"10", X"60", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"34", X"63", X"00", X"04", X"ac", X"43", X"10", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"34", X"63", X"00", X"02", X"ac", X"43", X"10", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"66", X"18", X"24", X"ac", X"43", X"10", X"00", 
  X"10", X"85", X"00", X"77", X"00", X"00", X"00", X"00", 
  X"90", X"83", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"03", X"46", X"00", X"00", X"08", X"46", X"03", 
  X"05", X"00", X"00", X"73", X"24", X"84", X"00", X"01", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"40", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"20", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"10", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"08", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"04", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"30", X"68", X"00", X"02", 
  X"35", X"29", X"00", X"02", X"ac", X"49", X"10", X"00", 
  X"8c", X"49", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"26", X"48", X"24", X"ac", X"49", X"10", X"00", 
  X"15", X"00", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"30", X"63", X"00", X"01", 
  X"01", X"07", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"02", X"ac", X"48", X"10", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"01", X"06", X"40", X"24", X"ac", X"48", X"10", X"00", 
  X"14", X"60", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"67", X"18", X"24", X"ac", X"43", X"10", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"34", X"63", X"00", X"02", X"ac", X"43", X"10", X"00", 
  X"8c", X"43", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"66", X"18", X"24", X"ac", X"43", X"10", X"00", 
  X"14", X"85", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"8c", X"48", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"35", X"08", X"00", X"04", X"ac", X"48", X"10", X"00", 
  X"0b", X"f0", X"02", X"c0", X"00", X"00", X"00", X"00", 
  X"3c", X"02", X"20", X"00", X"8c", X"43", X"10", X"00", 
  X"00", X"85", X"28", X"21", X"34", X"63", X"00", X"04", 
  X"ac", X"43", X"10", X"00", X"24", X"03", X"ff", X"fd", 
  X"8c", X"46", X"10", X"04", X"8c", X"47", X"10", X"00", 
  X"30", X"c6", X"00", X"01", X"34", X"e7", X"00", X"02", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"00", 
  X"00", X"06", X"30", X"40", X"00", X"e3", X"38", X"24", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"03", X"30", X"c6", X"00", X"ff", 
  X"24", X"c6", X"00", X"01", X"30", X"c6", X"00", X"ff", 
  X"8c", X"47", X"10", X"00", X"00", X"06", X"30", X"40", 
  X"34", X"e7", X"00", X"02", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"e3", X"38", X"24", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"04", X"00", X"00", X"00", X"00", 
  X"30", X"e7", X"00", X"01", X"10", X"e0", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"24", X"c6", X"00", X"01", 
  X"30", X"c6", X"00", X"ff", X"8c", X"47", X"10", X"00", 
  X"00", X"06", X"30", X"40", X"34", X"e7", X"00", X"02", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"00", 
  X"30", X"c6", X"00", X"ff", X"00", X"e3", X"38", X"24", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"24", X"c6", X"00", X"01", X"30", X"c6", X"00", X"ff", 
  X"8c", X"47", X"10", X"00", X"00", X"06", X"30", X"40", 
  X"34", X"e7", X"00", X"02", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"00", X"30", X"c6", X"00", X"ff", 
  X"00", X"e3", X"38", X"24", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"04", X"00", X"00", X"00", X"00", 
  X"30", X"e7", X"00", X"01", X"10", X"e0", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"24", X"c6", X"00", X"01", 
  X"30", X"c6", X"00", X"ff", X"8c", X"47", X"10", X"00", 
  X"00", X"06", X"30", X"40", X"34", X"e7", X"00", X"02", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"00", 
  X"30", X"c6", X"00", X"ff", X"00", X"e3", X"38", X"24", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"24", X"c6", X"00", X"01", X"30", X"c6", X"00", X"ff", 
  X"8c", X"47", X"10", X"00", X"00", X"06", X"30", X"40", 
  X"34", X"e7", X"00", X"02", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"00", X"30", X"c6", X"00", X"ff", 
  X"00", X"e3", X"38", X"24", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"04", X"00", X"00", X"00", X"00", 
  X"30", X"e7", X"00", X"01", X"10", X"e0", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"24", X"c6", X"00", X"01", 
  X"30", X"c6", X"00", X"ff", X"8c", X"47", X"10", X"00", 
  X"00", X"06", X"30", X"40", X"34", X"e7", X"00", X"02", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"00", 
  X"30", X"c6", X"00", X"ff", X"00", X"e3", X"38", X"24", 
  X"ac", X"47", X"10", X"00", X"8c", X"47", X"10", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"24", X"c6", X"00", X"01", X"30", X"c6", X"00", X"ff", 
  X"8c", X"47", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"34", X"e7", X"00", X"02", X"ac", X"47", X"10", X"00", 
  X"8c", X"47", X"10", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"e3", X"38", X"24", X"ac", X"47", X"10", X"00", 
  X"a0", X"86", X"00", X"00", X"24", X"84", X"00", X"01", 
  X"14", X"85", X"ff", X"8b", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"02", X"20", X"00", X"8c", X"43", X"10", X"00", 
  X"27", X"bd", X"ff", X"e0", X"34", X"63", X"00", X"01", 
  X"af", X"bf", X"00", X"1c", X"27", X"a4", X"00", X"10", 
  X"24", X"05", X"00", X"01", X"ac", X"43", X"10", X"00", 
  X"0f", X"f0", X"03", X"34", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"f8", X"af", X"a0", X"00", X"00", 
  X"00", X"04", X"18", X"c0", X"8f", X"a2", X"00", X"00", 
  X"00", X"04", X"21", X"40", X"00", X"64", X"20", X"21", 
  X"00", X"44", X"10", X"2b", X"10", X"40", X"00", X"0f", 
  X"00", X"00", X"00", X"00", X"3c", X"03", X"00", X"08", 
  X"8f", X"a2", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"24", X"42", X"00", X"07", X"ac", X"62", X"c0", X"00", 
  X"8f", X"a2", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"24", X"42", X"00", X"01", X"af", X"a2", X"00", X"00", 
  X"8f", X"a2", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"00", X"44", X"10", X"2b", X"14", X"40", X"ff", X"f4", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"08", X"27", X"bd", X"ff", X"d8", 
  X"af", X"b1", X"00", X"20", X"af", X"b0", X"00", X"1c", 
  X"af", X"bf", X"00", X"24", X"24", X"10", X"13", X"88", 
  X"0b", X"f0", X"03", X"e4", X"24", X"11", X"00", X"ff", 
  X"0f", X"f0", X"03", X"c0", X"26", X"10", X"ff", X"ff", 
  X"12", X"00", X"00", X"0e", X"00", X"00", X"10", X"21", 
  X"27", X"a4", X"00", X"10", X"0f", X"f0", X"03", X"34", 
  X"24", X"05", X"00", X"01", X"93", X"a2", X"00", X"10", 
  X"00", X"00", X"00", X"00", X"14", X"51", X"ff", X"f6", 
  X"24", X"04", X"00", X"64", X"8f", X"bf", X"00", X"24", 
  X"00", X"10", X"10", X"2b", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"8f", X"bf", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"3c", X"02", X"20", X"00", X"8c", X"44", X"10", X"00", 
  X"24", X"03", X"ff", X"fe", X"27", X"bd", X"ff", X"e0", 
  X"00", X"83", X"18", X"24", X"af", X"bf", X"00", X"1c", 
  X"27", X"a4", X"00", X"10", X"24", X"05", X"00", X"01", 
  X"ac", X"43", X"10", X"00", X"0f", X"f0", X"03", X"34", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"03", X"d9", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"05", 
  X"24", X"02", X"00", X"01", X"8f", X"bf", X"00", X"1c", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"0f", X"f0", X"03", X"b2", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"00", X"00", X"10", X"21", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"00", X"04", X"16", X"00", 
  X"27", X"bd", X"ff", X"d0", X"00", X"02", X"16", X"03", 
  X"af", X"b1", X"00", X"28", X"af", X"b0", X"00", X"24", 
  X"af", X"bf", X"00", X"2c", X"00", X"80", X"80", X"21", 
  X"04", X"40", X"00", X"44", X"00", X"a0", X"88", X"21", 
  X"0f", X"f0", X"03", X"b2", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"03", X"f6", X"00", X"00", X"00", X"00", 
  X"10", X"40", X"00", X"2b", X"36", X"05", X"00", X"40", 
  X"00", X"11", X"26", X"02", X"00", X"11", X"1c", X"02", 
  X"00", X"11", X"12", X"02", X"a3", X"a5", X"00", X"14", 
  X"a3", X"a4", X"00", X"15", X"a3", X"a3", X"00", X"16", 
  X"a3", X"a2", X"00", X"17", X"16", X"00", X"00", X"18", 
  X"a3", X"b1", X"00", X"18", X"24", X"02", X"ff", X"95", 
  X"27", X"a4", X"00", X"14", X"24", X"05", X"00", X"06", 
  X"a3", X"a2", X"00", X"19", X"0f", X"f0", X"02", X"4f", 
  X"27", X"b1", X"00", X"10", X"24", X"10", X"00", X"0a", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"03", X"34", 
  X"24", X"05", X"00", X"01", X"93", X"a2", X"00", X"10", 
  X"26", X"10", X"ff", X"ff", X"00", X"02", X"1e", X"00", 
  X"00", X"03", X"1e", X"03", X"04", X"61", X"00", X"03", 
  X"32", X"10", X"00", X"ff", X"16", X"00", X"ff", X"f7", 
  X"02", X"20", X"20", X"21", X"8f", X"bf", X"00", X"2c", 
  X"8f", X"b1", X"00", X"28", X"8f", X"b0", X"00", X"24", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"24", X"02", X"00", X"08", X"16", X"02", X"00", X"0e", 
  X"24", X"02", X"ff", X"87", X"27", X"a4", X"00", X"14", 
  X"24", X"05", X"00", X"06", X"a3", X"a2", X"00", X"19", 
  X"0f", X"f0", X"02", X"4f", X"27", X"b1", X"00", X"10", 
  X"0b", X"f0", X"04", X"2e", X"24", X"10", X"00", X"0a", 
  X"8f", X"bf", X"00", X"2c", X"24", X"02", X"00", X"ff", 
  X"8f", X"b1", X"00", X"28", X"8f", X"b0", X"00", X"24", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"24", X"02", X"00", X"01", X"27", X"a4", X"00", X"14", 
  X"24", X"05", X"00", X"06", X"0f", X"f0", X"02", X"4f", 
  X"a3", X"a2", X"00", X"19", X"24", X"02", X"00", X"0c", 
  X"16", X"02", X"ff", X"d8", X"27", X"b1", X"00", X"10", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"03", X"34", 
  X"24", X"05", X"00", X"01", X"0b", X"f0", X"04", X"2e", 
  X"24", X"10", X"00", X"0a", X"24", X"04", X"00", X"37", 
  X"0f", X"f0", X"04", X"0f", X"00", X"00", X"28", X"21", 
  X"2c", X"43", X"00", X"02", X"10", X"60", X"ff", X"d9", 
  X"32", X"10", X"00", X"7f", X"0b", X"f0", X"04", X"18", 
  X"00", X"00", X"00", X"00", X"27", X"bd", X"ff", X"d8", 
  X"30", X"84", X"00", X"ff", X"af", X"bf", X"00", X"24", 
  X"af", X"b1", X"00", X"20", X"14", X"80", X"00", X"0e", 
  X"af", X"b0", X"00", X"1c", X"3c", X"11", X"00", X"08", 
  X"92", X"30", X"bf", X"fc", X"00", X"00", X"00", X"00", 
  X"32", X"02", X"00", X"01", X"10", X"40", X"00", X"0f", 
  X"24", X"04", X"00", X"0d", X"8f", X"bf", X"00", X"24", 
  X"a2", X"30", X"bf", X"fc", X"02", X"00", X"10", X"21", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"8f", X"bf", X"00", X"24", X"24", X"10", X"00", X"01", 
  X"02", X"00", X"10", X"21", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"0f", X"f0", X"04", X"0f", 
  X"00", X"00", X"28", X"21", X"10", X"40", X"00", X"02", 
  X"27", X"a4", X"00", X"10", X"24", X"10", X"00", X"01", 
  X"0f", X"f0", X"03", X"34", X"24", X"05", X"00", X"01", 
  X"0f", X"f0", X"03", X"b2", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"04", X"6f", X"00", X"00", X"00", X"00", 
  X"27", X"bd", X"ff", X"d8", X"af", X"b1", X"00", X"20", 
  X"af", X"b0", X"00", X"1c", X"af", X"bf", X"00", X"24", 
  X"00", X"80", X"88", X"21", X"0f", X"f0", X"03", X"d9", 
  X"00", X"a0", X"80", X"21", X"14", X"40", X"00", X"06", 
  X"00", X"00", X"10", X"21", X"8f", X"bf", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"27", X"a4", X"00", X"10", X"24", X"05", X"00", X"01", 
  X"0f", X"f0", X"02", X"4f", X"a3", X"b0", X"00", X"10", 
  X"24", X"02", X"00", X"fd", X"12", X"02", X"00", X"12", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"02", X"4f", 
  X"24", X"05", X"02", X"00", X"27", X"a4", X"00", X"10", 
  X"0f", X"f0", X"03", X"34", X"24", X"05", X"00", X"02", 
  X"27", X"a4", X"00", X"10", X"0f", X"f0", X"03", X"34", 
  X"24", X"05", X"00", X"01", X"93", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"24", X"30", X"42", X"00", X"1f", 
  X"38", X"42", X"00", X"05", X"2c", X"42", X"00", X"01", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"8f", X"bf", X"00", X"24", X"24", X"02", X"00", X"01", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"27", X"bd", X"ff", X"d8", X"30", X"84", X"00", X"ff", 
  X"af", X"b1", X"00", X"20", X"af", X"b0", X"00", X"1c", 
  X"af", X"a6", X"00", X"10", X"af", X"bf", X"00", X"24", 
  X"00", X"a0", X"80", X"21", X"0f", X"f0", X"04", X"63", 
  X"30", X"f1", X"00", X"ff", X"30", X"42", X"00", X"01", 
  X"8f", X"a6", X"00", X"10", X"14", X"40", X"00", X"30", 
  X"24", X"02", X"00", X"03", X"12", X"20", X"00", X"28", 
  X"3c", X"02", X"00", X"08", X"90", X"42", X"c0", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"43", X"00", X"08", 
  X"14", X"60", X"00", X"02", X"24", X"03", X"00", X"01", 
  X"00", X"06", X"32", X"40", X"12", X"23", X"00", X"31", 
  X"30", X"42", X"00", X"06", X"14", X"40", X"00", X"29", 
  X"24", X"04", X"00", X"97", X"24", X"04", X"00", X"19", 
  X"0f", X"f0", X"04", X"0f", X"00", X"c0", X"28", X"21", 
  X"10", X"40", X"00", X"0b", X"02", X"00", X"20", X"21", 
  X"24", X"02", X"00", X"01", X"0f", X"f0", X"03", X"b2", 
  X"af", X"a2", X"00", X"10", X"8f", X"bf", X"00", X"24", 
  X"8f", X"a2", X"00", X"10", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"04", X"88", X"24", X"05", X"00", X"fc", 
  X"10", X"40", X"00", X"04", X"26", X"23", X"ff", X"ff", 
  X"30", X"71", X"00", X"ff", X"16", X"20", X"ff", X"f9", 
  X"26", X"10", X"02", X"00", X"00", X"00", X"20", X"21", 
  X"0f", X"f0", X"04", X"88", X"24", X"05", X"00", X"fd", 
  X"10", X"40", X"ff", X"eb", X"00", X"11", X"10", X"2b", 
  X"0b", X"f0", X"04", X"d3", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"24", X"24", X"02", X"00", X"04", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"8f", X"bf", X"00", X"24", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"02", X"20", X"28", X"21", 
  X"0f", X"f0", X"04", X"0f", X"af", X"a6", X"00", X"10", 
  X"8f", X"a6", X"00", X"10", X"0b", X"f0", X"04", X"ce", 
  X"24", X"04", X"00", X"19", X"24", X"04", X"00", X"18", 
  X"0f", X"f0", X"04", X"0f", X"00", X"c0", X"28", X"21", 
  X"14", X"40", X"ff", X"d3", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"04", X"88", X"24", X"05", X"00", X"fe", 
  X"0b", X"f0", X"04", X"d3", X"2c", X"42", X"00", X"01", 
  X"27", X"bd", X"ff", X"d0", X"af", X"b3", X"00", X"28", 
  X"af", X"b2", X"00", X"24", X"af", X"b1", X"00", X"20", 
  X"af", X"b0", X"00", X"1c", X"af", X"bf", X"00", X"2c", 
  X"00", X"80", X"90", X"21", X"00", X"a0", X"98", X"21", 
  X"24", X"10", X"03", X"e8", X"0b", X"f0", X"05", X"13", 
  X"24", X"11", X"00", X"ff", X"0f", X"f0", X"03", X"c0", 
  X"00", X"00", X"00", X"00", X"12", X"00", X"00", X"20", 
  X"00", X"00", X"00", X"00", X"27", X"a4", X"00", X"10", 
  X"0f", X"f0", X"03", X"34", X"24", X"05", X"00", X"01", 
  X"93", X"a2", X"00", X"10", X"24", X"04", X"00", X"64", 
  X"10", X"51", X"ff", X"f6", X"26", X"10", X"ff", X"ff", 
  X"24", X"03", X"00", X"fe", X"10", X"43", X"00", X"08", 
  X"00", X"00", X"10", X"21", X"8f", X"bf", X"00", X"2c", 
  X"8f", X"b3", X"00", X"28", X"8f", X"b2", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"02", X"60", X"28", X"21", X"0f", X"f0", X"03", X"34", 
  X"02", X"40", X"20", X"21", X"27", X"a4", X"00", X"10", 
  X"0f", X"f0", X"03", X"34", X"24", X"05", X"00", X"02", 
  X"8f", X"bf", X"00", X"2c", X"24", X"02", X"00", X"01", 
  X"8f", X"b3", X"00", X"28", X"8f", X"b2", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"93", X"a2", X"00", X"10", X"0b", X"f0", X"05", X"1b", 
  X"24", X"03", X"00", X"fe", X"27", X"bd", X"ff", X"d0", 
  X"30", X"84", X"00", X"ff", X"af", X"b0", X"00", X"28", 
  X"af", X"a6", X"00", X"20", X"af", X"bf", X"00", X"2c", 
  X"0f", X"f0", X"04", X"63", X"30", X"b0", X"00", X"ff", 
  X"30", X"42", X"00", X"01", X"8f", X"a6", X"00", X"20", 
  X"14", X"40", X"00", X"11", X"24", X"02", X"00", X"01", 
  X"12", X"02", X"00", X"18", X"24", X"04", X"00", X"09", 
  X"16", X"00", X"00", X"12", X"24", X"02", X"00", X"03", 
  X"0f", X"f0", X"03", X"f6", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"00", X"3e", X"00", X"00", X"00", X"00", 
  X"24", X"02", X"00", X"01", X"0f", X"f0", X"03", X"b2", 
  X"af", X"a2", X"00", X"20", X"8f", X"bf", X"00", X"2c", 
  X"8f", X"a2", X"00", X"20", X"8f", X"b0", X"00", X"28", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"8f", X"bf", X"00", X"2c", X"24", X"02", X"00", X"03", 
  X"8f", X"b0", X"00", X"28", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"12", X"02", X"00", X"2b", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"05", X"49", 
  X"24", X"02", X"00", X"04", X"00", X"00", X"28", X"21", 
  X"0f", X"f0", X"04", X"0f", X"af", X"a6", X"00", X"20", 
  X"14", X"40", X"ff", X"ec", X"24", X"02", X"00", X"01", 
  X"27", X"a4", X"00", X"10", X"0f", X"f0", X"05", X"04", 
  X"24", X"05", X"00", X"10", X"8f", X"a6", X"00", X"20", 
  X"10", X"40", X"ff", X"e6", X"24", X"02", X"00", X"01", 
  X"93", X"a2", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"00", X"02", X"11", X"82", X"10", X"50", X"00", X"21", 
  X"00", X"00", X"00", X"00", X"93", X"a8", X"00", X"18", 
  X"93", X"a4", X"00", X"17", X"93", X"a5", X"00", X"1a", 
  X"93", X"a7", X"00", X"15", X"93", X"a2", X"00", X"19", 
  X"93", X"a3", X"00", X"16", X"00", X"08", X"41", X"82", 
  X"00", X"04", X"20", X"80", X"30", X"e7", X"00", X"0f", 
  X"00", X"05", X"29", X"c2", X"30", X"42", X"00", X"03", 
  X"01", X"04", X"20", X"21", X"30", X"63", X"00", X"03", 
  X"00", X"e5", X"28", X"21", X"00", X"02", X"10", X"40", 
  X"24", X"84", X"00", X"01", X"00", X"03", X"1a", X"80", 
  X"00", X"a2", X"10", X"21", X"00", X"83", X"18", X"21", 
  X"24", X"42", X"ff", X"f9", X"00", X"43", X"10", X"04", 
  X"ac", X"c2", X"00", X"00", X"0b", X"f0", X"05", X"49", 
  X"00", X"00", X"10", X"21", X"24", X"02", X"00", X"80", 
  X"ac", X"c2", X"00", X"00", X"0b", X"f0", X"05", X"49", 
  X"00", X"00", X"10", X"21", X"0f", X"f0", X"03", X"b2", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"05", X"49", 
  X"00", X"00", X"10", X"21", X"93", X"a3", X"00", X"17", 
  X"93", X"a2", X"00", X"18", X"93", X"a4", X"00", X"19", 
  X"30", X"63", X"00", X"3f", X"00", X"03", X"1a", X"00", 
  X"00", X"02", X"12", X"00", X"24", X"63", X"00", X"01", 
  X"00", X"44", X"10", X"21", X"00", X"62", X"10", X"21", 
  X"00", X"02", X"12", X"80", X"ac", X"c2", X"00", X"00", 
  X"0b", X"f0", X"05", X"49", X"00", X"00", X"10", X"21", 
  X"27", X"bd", X"ff", X"d8", X"30", X"84", X"00", X"ff", 
  X"af", X"b1", X"00", X"20", X"af", X"b0", X"00", X"1c", 
  X"af", X"a6", X"00", X"10", X"af", X"bf", X"00", X"24", 
  X"00", X"a0", X"80", X"21", X"0f", X"f0", X"04", X"63", 
  X"30", X"f1", X"00", X"ff", X"30", X"42", X"00", X"01", 
  X"8f", X"a6", X"00", X"10", X"14", X"40", X"00", X"2b", 
  X"24", X"02", X"00", X"03", X"12", X"20", X"00", X"23", 
  X"3c", X"02", X"00", X"08", X"90", X"42", X"c0", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"42", X"00", X"08", 
  X"14", X"40", X"00", X"02", X"24", X"02", X"00", X"01", 
  X"00", X"06", X"32", X"40", X"12", X"22", X"00", X"26", 
  X"24", X"04", X"00", X"12", X"0f", X"f0", X"04", X"0f", 
  X"00", X"c0", X"28", X"21", X"10", X"40", X"00", X"0b", 
  X"02", X"00", X"20", X"21", X"24", X"02", X"00", X"01", 
  X"0f", X"f0", X"03", X"b2", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"24", X"8f", X"a2", X"00", X"10", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"02", X"00", X"20", X"21", X"0f", X"f0", X"05", X"04", 
  X"24", X"05", X"02", X"00", X"10", X"40", X"00", X"04", 
  X"26", X"23", X"ff", X"ff", X"30", X"71", X"00", X"ff", 
  X"16", X"20", X"ff", X"f9", X"26", X"10", X"02", X"00", 
  X"24", X"04", X"00", X"0c", X"0f", X"f0", X"04", X"0f", 
  X"00", X"00", X"28", X"21", X"0b", X"f0", X"05", X"b2", 
  X"00", X"11", X"10", X"2b", X"8f", X"bf", X"00", X"24", 
  X"24", X"02", X"00", X"04", X"8f", X"b1", X"00", X"20", 
  X"8f", X"b0", X"00", X"1c", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"8f", X"bf", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"24", X"04", X"00", X"11", X"0f", X"f0", X"04", X"0f", 
  X"00", X"c0", X"28", X"21", X"14", X"40", X"ff", X"db", 
  X"02", X"00", X"20", X"21", X"0f", X"f0", X"05", X"04", 
  X"24", X"05", X"02", X"00", X"0b", X"f0", X"05", X"b2", 
  X"2c", X"42", X"00", X"01", X"27", X"bd", X"ff", X"d0", 
  X"30", X"84", X"00", X"ff", X"af", X"bf", X"00", X"2c", 
  X"af", X"b2", X"00", X"28", X"af", X"b1", X"00", X"24", 
  X"14", X"80", X"00", X"22", X"af", X"b0", X"00", X"20", 
  X"24", X"03", X"00", X"05", X"3c", X"02", X"20", X"00", 
  X"ac", X"43", X"10", X"00", X"24", X"10", X"00", X"0a", 
  X"26", X"10", X"ff", X"ff", X"27", X"a4", X"00", X"10", 
  X"24", X"05", X"00", X"01", X"0f", X"f0", X"03", X"34", 
  X"32", X"10", X"00", X"ff", X"16", X"00", X"ff", X"fb", 
  X"26", X"10", X"ff", X"ff", X"00", X"00", X"20", X"21", 
  X"0f", X"f0", X"04", X"0f", X"00", X"00", X"28", X"21", 
  X"00", X"40", X"80", X"21", X"24", X"02", X"00", X"01", 
  X"12", X"02", X"00", X"17", X"24", X"04", X"00", X"08", 
  X"24", X"02", X"00", X"01", X"00", X"00", X"88", X"21", 
  X"3c", X"03", X"00", X"08", X"a0", X"71", X"c0", X"04", 
  X"3c", X"03", X"00", X"08", X"af", X"a2", X"00", X"18", 
  X"0f", X"f0", X"03", X"b2", X"a0", X"62", X"bf", X"fc", 
  X"8f", X"bf", X"00", X"2c", X"8f", X"a2", X"00", X"18", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"8f", X"bf", X"00", X"2c", 
  X"24", X"02", X"00", X"03", X"8f", X"b2", X"00", X"28", 
  X"8f", X"b1", X"00", X"24", X"8f", X"b0", X"00", X"20", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"30", 
  X"0f", X"f0", X"04", X"0f", X"24", X"05", X"01", X"aa", 
  X"10", X"50", X"00", X"1e", X"24", X"04", X"00", X"a9", 
  X"0f", X"f0", X"04", X"0f", X"00", X"00", X"28", X"21", 
  X"2c", X"42", X"00", X"02", X"14", X"40", X"00", X"16", 
  X"00", X"00", X"00", X"00", X"24", X"12", X"00", X"01", 
  X"24", X"11", X"00", X"01", X"0b", X"f0", X"06", X"1b", 
  X"24", X"10", X"03", X"e8", X"0f", X"f0", X"03", X"c0", 
  X"00", X"00", X"00", X"00", X"12", X"00", X"ff", X"db", 
  X"24", X"02", X"00", X"01", X"02", X"40", X"20", X"21", 
  X"0f", X"f0", X"04", X"0f", X"00", X"00", X"28", X"21", 
  X"26", X"10", X"ff", X"ff", X"14", X"40", X"ff", X"f7", 
  X"24", X"04", X"03", X"e8", X"24", X"04", X"00", X"10", 
  X"0f", X"f0", X"04", X"0f", X"24", X"05", X"02", X"00", 
  X"14", X"40", X"ff", X"cf", X"3c", X"03", X"00", X"08", 
  X"0b", X"f0", X"05", X"f8", X"a0", X"71", X"c0", X"04", 
  X"24", X"12", X"00", X"a9", X"0b", X"f0", X"06", X"15", 
  X"24", X"11", X"00", X"02", X"27", X"a4", X"00", X"10", 
  X"24", X"05", X"00", X"04", X"0f", X"f0", X"03", X"34", 
  X"af", X"a2", X"00", X"18", X"93", X"a3", X"00", X"12", 
  X"8f", X"a2", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"14", X"62", X"ff", X"c2", X"24", X"02", X"00", X"01", 
  X"93", X"a3", X"00", X"13", X"24", X"02", X"00", X"aa", 
  X"14", X"62", X"ff", X"be", X"24", X"02", X"00", X"01", 
  X"0b", X"f0", X"06", X"3e", X"24", X"10", X"03", X"e8", 
  X"0f", X"f0", X"03", X"c0", X"00", X"00", X"00", X"00", 
  X"12", X"00", X"ff", X"b8", X"24", X"02", X"00", X"01", 
  X"24", X"04", X"00", X"a9", X"0f", X"f0", X"04", X"0f", 
  X"3c", X"05", X"40", X"00", X"26", X"10", X"ff", X"ff", 
  X"14", X"40", X"ff", X"f7", X"24", X"04", X"03", X"e8", 
  X"24", X"04", X"00", X"3a", X"0f", X"f0", X"04", X"0f", 
  X"00", X"00", X"28", X"21", X"14", X"40", X"ff", X"ad", 
  X"24", X"02", X"00", X"01", X"27", X"a4", X"00", X"10", 
  X"0f", X"f0", X"03", X"34", X"24", X"05", X"00", X"04", 
  X"93", X"a2", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"30", X"42", X"00", X"40", X"10", X"40", X"00", X"03", 
  X"00", X"00", X"10", X"21", X"0b", X"f0", X"05", X"f6", 
  X"24", X"11", X"00", X"0c", X"0b", X"f0", X"05", X"f6", 
  X"24", X"11", X"00", X"04", X"03", X"e0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"8c", X"82", X"00", X"00", 
  X"27", X"bd", X"ff", X"e8", X"10", X"40", X"00", X"0a", 
  X"af", X"bf", X"00", X"14", X"90", X"43", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"00", X"06", 
  X"00", X"00", X"00", X"00", X"94", X"45", X"00", X"06", 
  X"94", X"83", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"10", X"a3", X"00", X"06", X"00", X"00", X"00", X"00", 
  X"24", X"02", X"00", X"09", X"8f", X"bf", X"00", X"14", 
  X"00", X"00", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"18", X"90", X"44", X"00", X"01", 
  X"0f", X"f0", X"04", X"63", X"00", X"00", X"00", X"00", 
  X"30", X"42", X"00", X"01", X"14", X"40", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"06", X"65", 
  X"00", X"00", X"10", X"21", X"0b", X"f0", X"06", X"65", 
  X"24", X"02", X"00", X"03", X"8c", X"82", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"18", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"1c", 
  X"00", X"80", X"88", X"21", X"10", X"45", X"00", X"03", 
  X"00", X"a0", X"80", X"21", X"14", X"a0", X"00", X"07", 
  X"26", X"25", X"00", X"24", X"8f", X"bf", X"00", X"1c", 
  X"00", X"00", X"10", X"21", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"90", X"84", X"00", X"01", 
  X"02", X"00", X"30", X"21", X"0f", X"f0", X"05", X"96", 
  X"24", X"07", X"00", X"01", X"14", X"40", X"00", X"07", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"ae", X"30", X"00", X"20", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8f", X"bf", X"00", X"1c", 
  X"24", X"02", X"00", X"01", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"27", X"bd", X"ff", X"e8", 
  X"af", X"b0", X"00", X"10", X"af", X"bf", X"00", X"14", 
  X"00", X"80", X"80", X"21", X"90", X"84", X"00", X"01", 
  X"00", X"a0", X"30", X"21", X"24", X"07", X"00", X"01", 
  X"0f", X"f0", X"05", X"96", X"26", X"05", X"00", X"24", 
  X"14", X"40", X"00", X"30", X"24", X"02", X"00", X"03", 
  X"92", X"03", X"02", X"23", X"92", X"02", X"02", X"22", 
  X"00", X"03", X"1a", X"00", X"00", X"62", X"18", X"25", 
  X"00", X"03", X"1c", X"00", X"00", X"03", X"1c", X"03", 
  X"24", X"02", X"aa", X"55", X"10", X"62", X"00", X"05", 
  X"24", X"02", X"00", X"02", X"8f", X"bf", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"18", X"92", X"05", X"00", X"5d", 
  X"92", X"04", X"00", X"5c", X"92", X"03", X"00", X"5a", 
  X"00", X"04", X"24", X"00", X"00", X"05", X"2e", X"00", 
  X"92", X"02", X"00", X"5b", X"00", X"a4", X"28", X"25", 
  X"00", X"a3", X"28", X"25", X"00", X"02", X"12", X"00", 
  X"3c", X"04", X"00", X"ff", X"00", X"a2", X"28", X"25", 
  X"34", X"84", X"ff", X"ff", X"3c", X"03", X"00", X"54", 
  X"00", X"a4", X"28", X"24", X"24", X"63", X"41", X"46", 
  X"10", X"a3", X"ff", X"ec", X"00", X"00", X"10", X"21", 
  X"92", X"07", X"00", X"79", X"92", X"02", X"00", X"78", 
  X"92", X"06", X"00", X"76", X"92", X"05", X"00", X"77", 
  X"00", X"07", X"3e", X"00", X"00", X"02", X"14", X"00", 
  X"00", X"e2", X"10", X"25", X"00", X"46", X"10", X"25", 
  X"00", X"05", X"2a", X"00", X"00", X"45", X"10", X"25", 
  X"00", X"44", X"10", X"24", X"8f", X"bf", X"00", X"14", 
  X"00", X"43", X"10", X"23", X"00", X"02", X"10", X"2b", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"18", X"8f", X"bf", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"18", X"90", X"a2", X"00", X"1b", 
  X"90", X"a3", X"00", X"1a", X"00", X"02", X"12", X"00", 
  X"00", X"43", X"10", X"25", X"24", X"03", X"00", X"03", 
  X"10", X"83", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"90", X"a3", X"00", X"15", X"90", X"a4", X"00", X"14", 
  X"00", X"03", X"1a", X"00", X"00", X"64", X"18", X"25", 
  X"00", X"03", X"1c", X"00", X"03", X"e0", X"00", X"08", 
  X"00", X"43", X"10", X"25", X"27", X"bd", X"ff", X"e0", 
  X"8c", X"82", X"00", X"00", X"af", X"bf", X"00", X"1c", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"90", X"43", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"24", X"63", X"ff", X"d0", X"2c", X"66", X"00", X"0a", 
  X"10", X"c0", X"00", X"05", X"24", X"06", X"00", X"3a", 
  X"90", X"47", X"00", X"01", X"00", X"00", X"00", X"00", 
  X"10", X"e6", X"00", X"2d", X"24", X"42", X"00", X"02", 
  X"ac", X"a0", X"00", X"00", X"3c", X"02", X"00", X"08", 
  X"8c", X"50", X"c0", X"08", X"00", X"00", X"00", X"00", 
  X"12", X"00", X"00", X"0d", X"24", X"02", X"00", X"0c", 
  X"ac", X"b0", X"00", X"00", X"92", X"02", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"14", X"40", X"00", X"1a", 
  X"00", X"00", X"00", X"00", X"a2", X"00", X"00", X"00", 
  X"a2", X"00", X"00", X"01", X"0f", X"f0", X"05", X"db", 
  X"00", X"00", X"20", X"21", X"30", X"42", X"00", X"01", 
  X"10", X"40", X"00", X"06", X"24", X"02", X"00", X"03", 
  X"8f", X"bf", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"06", X"95", X"00", X"00", X"28", X"21", 
  X"92", X"02", X"01", X"e6", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"1c", X"24", X"02", X"00", X"0d", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"92", X"04", X"00", X"01", X"0f", X"f0", X"04", X"63", 
  X"00", X"00", X"00", X"00", X"30", X"42", X"00", X"01", 
  X"14", X"40", X"ff", X"e2", X"00", X"00", X"10", X"21", 
  X"0b", X"f0", X"07", X"04", X"00", X"00", X"00", X"00", 
  X"ac", X"82", X"00", X"00", X"10", X"60", X"ff", X"d3", 
  X"ac", X"a0", X"00", X"00", X"8f", X"bf", X"00", X"1c", 
  X"24", X"02", X"00", X"0b", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"92", X"11", X"01", X"ed", 
  X"92", X"04", X"01", X"ec", X"92", X"03", X"01", X"ea", 
  X"00", X"04", X"24", X"00", X"92", X"02", X"01", X"eb", 
  X"00", X"11", X"8e", X"00", X"02", X"24", X"88", X"25", 
  X"02", X"23", X"88", X"25", X"00", X"02", X"12", X"00", 
  X"02", X"22", X"88", X"25", X"02", X"00", X"20", X"21", 
  X"0f", X"f0", X"06", X"95", X"02", X"20", X"28", X"21", 
  X"24", X"03", X"00", X"03", X"14", X"43", X"00", X"03", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"07", X"04", 
  X"24", X"02", X"00", X"01", X"14", X"40", X"ff", X"d6", 
  X"00", X"00", X"00", X"00", X"92", X"03", X"00", X"30", 
  X"92", X"02", X"00", X"2f", X"00", X"03", X"1a", X"00", 
  X"00", X"62", X"18", X"25", X"00", X"03", X"1c", X"00", 
  X"00", X"03", X"1c", X"03", X"24", X"02", X"02", X"00", 
  X"14", X"62", X"ff", X"cd", X"00", X"00", X"00", X"00", 
  X"92", X"02", X"00", X"3b", X"92", X"03", X"00", X"3a", 
  X"00", X"02", X"12", X"00", X"00", X"43", X"10", X"25", 
  X"14", X"40", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"92", X"05", X"00", X"4b", X"92", X"02", X"00", X"4a", 
  X"00", X"05", X"2e", X"00", X"00", X"02", X"14", X"00", 
  X"92", X"04", X"00", X"48", X"92", X"03", X"00", X"49", 
  X"00", X"a2", X"10", X"25", X"00", X"44", X"10", X"25", 
  X"00", X"03", X"1a", X"00", X"00", X"43", X"10", X"25", 
  X"92", X"08", X"00", X"34", X"ae", X"02", X"00", X"10", 
  X"25", X"03", X"ff", X"ff", X"30", X"63", X"00", X"ff", 
  X"2c", X"63", X"00", X"02", X"10", X"60", X"ff", X"b6", 
  X"a2", X"08", X"00", X"03", X"92", X"03", X"00", X"31", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"ff", X"b2", 
  X"a2", X"03", X"00", X"02", X"24", X"64", X"ff", X"ff", 
  X"00", X"83", X"20", X"24", X"14", X"80", X"ff", X"ae", 
  X"00", X"00", X"00", X"00", X"92", X"04", X"00", X"36", 
  X"92", X"05", X"00", X"35", X"00", X"04", X"22", X"00", 
  X"00", X"85", X"20", X"25", X"30", X"85", X"00", X"0f", 
  X"14", X"a0", X"ff", X"a7", X"a6", X"04", X"00", X"08", 
  X"92", X"05", X"00", X"38", X"92", X"06", X"00", X"37", 
  X"00", X"05", X"2a", X"00", X"00", X"a6", X"28", X"25", 
  X"14", X"a0", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"92", X"09", X"00", X"47", X"92", X"06", X"00", X"46", 
  X"00", X"09", X"4e", X"00", X"00", X"06", X"34", X"00", 
  X"92", X"07", X"00", X"44", X"92", X"05", X"00", X"45", 
  X"01", X"26", X"30", X"25", X"00", X"c7", X"30", X"25", 
  X"00", X"05", X"2a", X"00", X"00", X"c5", X"28", X"25", 
  X"92", X"06", X"00", X"33", X"92", X"07", X"00", X"32", 
  X"00", X"06", X"32", X"00", X"00", X"c7", X"30", X"25", 
  X"10", X"c0", X"ff", X"91", X"00", X"48", X"00", X"18", 
  X"00", X"04", X"39", X"02", X"00", X"e6", X"38", X"21", 
  X"00", X"00", X"40", X"12", X"00", X"e8", X"38", X"21", 
  X"00", X"a7", X"48", X"2b", X"15", X"20", X"ff", X"8a", 
  X"00", X"00", X"00", X"00", X"00", X"a7", X"28", X"23", 
  X"14", X"60", X"00", X"02", X"00", X"a3", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"00", X"00", X"18", X"12", 
  X"10", X"60", X"ff", X"83", X"00", X"00", X"00", X"00", 
  X"2c", X"65", X"0f", X"f6", X"14", X"a0", X"00", X"27", 
  X"24", X"05", X"00", X"01", X"34", X"05", X"ff", X"f6", 
  X"00", X"65", X"28", X"2b", X"14", X"a0", X"00", X"23", 
  X"24", X"05", X"00", X"02", X"24", X"63", X"00", X"02", 
  X"00", X"f1", X"38", X"21", X"00", X"d1", X"30", X"21", 
  X"ae", X"03", X"00", X"0c", X"ae", X"07", X"00", X"1c", 
  X"14", X"80", X"ff", X"75", X"ae", X"06", X"00", X"14", 
  X"92", X"07", X"00", X"53", X"92", X"05", X"00", X"52", 
  X"00", X"07", X"3e", X"00", X"00", X"05", X"2c", X"00", 
  X"92", X"06", X"00", X"50", X"92", X"04", X"00", X"51", 
  X"00", X"e5", X"28", X"25", X"00", X"a6", X"28", X"25", 
  X"00", X"04", X"22", X"00", X"00", X"a4", X"20", X"25", 
  X"ae", X"04", X"00", X"18", X"00", X"03", X"18", X"80", 
  X"24", X"05", X"00", X"03", X"24", X"63", X"01", X"ff", 
  X"00", X"03", X"1a", X"42", X"00", X"43", X"10", X"2b", 
  X"14", X"40", X"ff", X"63", X"3c", X"03", X"00", X"08", 
  X"a2", X"05", X"00", X"00", X"94", X"62", X"c0", X"0c", 
  X"ae", X"00", X"00", X"20", X"24", X"42", X"00", X"01", 
  X"a4", X"62", X"c0", X"0c", X"a6", X"02", X"00", X"06", 
  X"a2", X"00", X"00", X"04", X"0b", X"f0", X"07", X"04", 
  X"00", X"00", X"10", X"21", X"24", X"63", X"00", X"02", 
  X"00", X"f1", X"38", X"21", X"00", X"d1", X"30", X"21", 
  X"ae", X"03", X"00", X"0c", X"ae", X"07", X"00", X"1c", 
  X"10", X"80", X"ff", X"53", X"ae", X"06", X"00", X"14", 
  X"01", X"06", X"30", X"21", X"24", X"04", X"00", X"02", 
  X"10", X"a4", X"00", X"09", X"ae", X"06", X"00", X"18", 
  X"24", X"04", X"00", X"03", X"00", X"64", X"00", X"18", 
  X"30", X"63", X"00", X"01", X"24", X"05", X"00", X"01", 
  X"00", X"00", X"20", X"12", X"00", X"04", X"20", X"42", 
  X"0b", X"f0", X"07", X"a9", X"00", X"83", X"18", X"21", 
  X"0b", X"f0", X"07", X"a9", X"00", X"03", X"18", X"40", 
  X"8c", X"83", X"00", X"0c", X"24", X"a5", X"ff", X"fe", 
  X"24", X"63", X"ff", X"fe", X"00", X"a3", X"18", X"2b", 
  X"10", X"60", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"90", X"83", X"00", X"02", X"8c", X"82", X"00", X"1c", 
  X"00", X"a3", X"00", X"18", X"00", X"00", X"28", X"12", 
  X"03", X"e0", X"00", X"08", X"00", X"a2", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"27", X"bd", X"ff", X"d8", X"2c", X"a2", X"00", X"02", 
  X"af", X"b1", X"00", X"18", X"af", X"b0", X"00", X"14", 
  X"af", X"bf", X"00", X"24", X"af", X"b3", X"00", X"20", 
  X"af", X"b2", X"00", X"1c", X"00", X"a0", X"80", X"21", 
  X"14", X"40", X"00", X"16", X"00", X"80", X"88", X"21", 
  X"8c", X"82", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"a2", X"10", X"2b", X"10", X"40", X"00", X"11", 
  X"24", X"03", X"00", X"02", X"90", X"82", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"43", X"00", X"15", 
  X"24", X"03", X"00", X"03", X"10", X"43", X"00", X"3b", 
  X"24", X"03", X"00", X"01", X"10", X"43", X"00", X"1f", 
  X"00", X"05", X"90", X"42", X"24", X"02", X"ff", X"ff", 
  X"8f", X"bf", X"00", X"24", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"8f", X"bf", X"00", X"24", 
  X"24", X"02", X"00", X"01", X"8f", X"b3", X"00", X"20", 
  X"8f", X"b2", X"00", X"1c", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"28", X"8c", X"82", X"00", X"14", 
  X"00", X"05", X"2a", X"02", X"0f", X"f0", X"06", X"73", 
  X"00", X"a2", X"28", X"21", X"14", X"40", X"ff", X"eb", 
  X"00", X"10", X"80", X"40", X"32", X"10", X"01", X"ff", 
  X"02", X"30", X"10", X"21", X"00", X"40", X"80", X"21", 
  X"90", X"42", X"00", X"25", X"92", X"03", X"00", X"24", 
  X"00", X"02", X"12", X"00", X"0b", X"f0", X"07", X"f2", 
  X"00", X"43", X"10", X"25", X"02", X"45", X"90", X"21", 
  X"8c", X"82", X"00", X"14", X"00", X"12", X"2a", X"42", 
  X"0f", X"f0", X"06", X"73", X"00", X"a2", X"28", X"21", 
  X"14", X"40", X"ff", X"dd", X"24", X"02", X"ff", X"ff", 
  X"26", X"53", X"00", X"01", X"8e", X"22", X"00", X"14", 
  X"32", X"52", X"01", X"ff", X"00", X"13", X"2a", X"42", 
  X"02", X"32", X"90", X"21", X"02", X"20", X"20", X"21", 
  X"92", X"52", X"00", X"24", X"0f", X"f0", X"06", X"73", 
  X"00", X"a2", X"28", X"21", X"14", X"40", X"ff", X"d1", 
  X"32", X"73", X"01", X"ff", X"02", X"33", X"88", X"21", 
  X"92", X"22", X"00", X"24", X"32", X"10", X"00", X"01", 
  X"00", X"02", X"12", X"00", X"12", X"00", X"00", X"1a", 
  X"00", X"52", X"10", X"25", X"0b", X"f0", X"07", X"f2", 
  X"00", X"02", X"11", X"02", X"8c", X"82", X"00", X"14", 
  X"00", X"05", X"29", X"c2", X"0f", X"f0", X"06", X"73", 
  X"00", X"a2", X"28", X"21", X"14", X"40", X"ff", X"c3", 
  X"00", X"10", X"80", X"80", X"32", X"10", X"01", X"ff", 
  X"02", X"30", X"10", X"21", X"90", X"43", X"00", X"26", 
  X"90", X"45", X"00", X"27", X"90", X"44", X"00", X"25", 
  X"00", X"03", X"1c", X"00", X"00", X"05", X"16", X"00", 
  X"02", X"30", X"80", X"21", X"00", X"62", X"10", X"25", 
  X"00", X"04", X"22", X"00", X"92", X"03", X"00", X"24", 
  X"00", X"44", X"10", X"25", X"00", X"43", X"10", X"25", 
  X"3c", X"03", X"0f", X"ff", X"34", X"63", X"ff", X"ff", 
  X"0b", X"f0", X"07", X"f2", X"00", X"43", X"10", X"24", 
  X"0b", X"f0", X"07", X"f2", X"30", X"42", X"0f", X"ff", 
  X"27", X"bd", X"ff", X"e0", X"af", X"b1", X"00", X"14", 
  X"94", X"91", X"00", X"06", X"af", X"b0", X"00", X"10", 
  X"26", X"31", X"00", X"01", X"32", X"31", X"ff", X"ff", 
  X"af", X"bf", X"00", X"1c", X"af", X"b2", X"00", X"18", 
  X"12", X"20", X"00", X"1f", X"00", X"80", X"80", X"21", 
  X"8c", X"82", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"10", X"40", X"00", X"1b", X"32", X"32", X"00", X"0f", 
  X"12", X"40", X"00", X"0e", X"24", X"42", X"00", X"01", 
  X"8c", X"84", X"00", X"00", X"00", X"12", X"91", X"40", 
  X"24", X"84", X"00", X"24", X"8f", X"bf", X"00", X"1c", 
  X"00", X"92", X"20", X"21", X"a6", X"11", X"00", X"06", 
  X"ae", X"04", X"00", X"14", X"00", X"00", X"10", X"21", 
  X"8f", X"b2", X"00", X"18", X"8f", X"b1", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8c", X"85", X"00", X"0c", 
  X"00", X"00", X"00", X"00", X"14", X"a0", X"00", X"0f", 
  X"ac", X"82", X"00", X"10", X"8c", X"84", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"94", X"82", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"02", X"22", X"10", X"2b", 
  X"14", X"40", X"ff", X"eb", X"00", X"12", X"91", X"40", 
  X"24", X"02", X"00", X"04", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b2", X"00", X"18", X"8f", X"b1", X"00", X"14", 
  X"8f", X"b0", X"00", X"10", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8c", X"84", X"00", X"00", 
  X"00", X"11", X"19", X"02", X"90", X"82", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"24", X"42", X"ff", X"ff", 
  X"00", X"43", X"10", X"24", X"14", X"40", X"ff", X"db", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"07", X"da", 
  X"00", X"00", X"00", X"00", X"2c", X"43", X"00", X"02", 
  X"14", X"60", X"00", X"18", X"24", X"03", X"ff", X"ff", 
  X"10", X"43", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"8e", X"04", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"8c", X"83", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"43", X"28", X"2b", X"10", X"a0", X"ff", X"e4", 
  X"24", X"63", X"ff", X"fe", X"24", X"45", X"ff", X"fe", 
  X"00", X"a3", X"18", X"2b", X"10", X"60", X"00", X"08", 
  X"ae", X"02", X"00", X"0c", X"90", X"83", X"00", X"02", 
  X"8c", X"82", X"00", X"1c", X"00", X"a3", X"00", X"18", 
  X"00", X"00", X"28", X"12", X"00", X"a2", X"10", X"21", 
  X"0b", X"f0", X"08", X"53", X"ae", X"02", X"00", X"10", 
  X"00", X"00", X"10", X"21", X"0b", X"f0", X"08", X"53", 
  X"ae", X"02", X"00", X"10", X"0b", X"f0", X"08", X"6b", 
  X"24", X"02", X"00", X"02", X"0b", X"f0", X"08", X"6b", 
  X"24", X"02", X"00", X"01", X"8c", X"82", X"00", X"08", 
  X"27", X"bd", X"ff", X"e0", X"24", X"03", X"00", X"01", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"1c", 
  X"af", X"b1", X"00", X"18", X"00", X"80", X"80", X"21", 
  X"10", X"43", X"00", X"1f", X"a4", X"80", X"00", X"06", 
  X"8c", X"84", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"8c", X"83", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"43", X"28", X"2b", X"10", X"a0", X"00", X"18", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"1c", 
  X"00", X"00", X"00", X"00", X"90", X"85", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"14", X"a0", X"00", X"31", 
  X"24", X"11", X"ff", X"ff", X"0b", X"f0", X"08", X"ba", 
  X"00", X"00", X"00", X"00", X"14", X"60", X"00", X"0e", 
  X"00", X"00", X"00", X"00", X"8e", X"04", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"8c", X"83", X"00", X"0c", 
  X"00", X"00", X"00", X"00", X"00", X"43", X"18", X"2b", 
  X"10", X"60", X"00", X"07", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"07", X"da", X"00", X"40", X"28", X"21", 
  X"14", X"51", X"ff", X"f4", X"2c", X"43", X"00", X"02", 
  X"0b", X"f0", X"08", X"c1", X"24", X"02", X"00", X"01", 
  X"24", X"02", X"00", X"02", X"8f", X"bf", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"90", X"85", X"00", X"00", X"24", X"02", X"00", X"03", 
  X"10", X"a2", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"94", X"82", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"10", X"40", X"ff", X"f3", X"ae", X"00", X"00", X"0c", 
  X"8c", X"82", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"ae", X"02", X"00", X"10", X"8f", X"bf", X"00", X"1c", 
  X"24", X"84", X"00", X"24", X"ae", X"04", X"00", X"14", 
  X"00", X"00", X"10", X"21", X"8f", X"b1", X"00", X"18", 
  X"8f", X"b0", X"00", X"14", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"20", X"8c", X"82", X"00", X"18", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"ff", X"ee", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"08", X"ab", 
  X"00", X"00", X"00", X"00", X"24", X"45", X"ff", X"fe", 
  X"24", X"63", X"ff", X"fe", X"00", X"a3", X"18", X"2b", 
  X"10", X"60", X"00", X"08", X"ae", X"02", X"00", X"0c", 
  X"90", X"83", X"00", X"02", X"8c", X"82", X"00", X"1c", 
  X"00", X"a3", X"00", X"18", X"00", X"00", X"28", X"12", 
  X"00", X"a2", X"10", X"21", X"0b", X"f0", X"08", X"d1", 
  X"ae", X"02", X"00", X"10", X"00", X"00", X"10", X"21", 
  X"0b", X"f0", X"08", X"d1", X"ae", X"02", X"00", X"10", 
  X"27", X"bd", X"ff", X"c8", X"af", X"b2", X"00", X"1c", 
  X"af", X"b0", X"00", X"14", X"af", X"bf", X"00", X"34", 
  X"af", X"b7", X"00", X"30", X"af", X"b6", X"00", X"2c", 
  X"af", X"b5", X"00", X"28", X"af", X"b4", X"00", X"24", 
  X"af", X"b3", X"00", X"20", X"af", X"b1", X"00", X"18", 
  X"90", X"a2", X"00", X"00", X"24", X"03", X"00", X"2f", 
  X"00", X"a0", X"80", X"21", X"10", X"43", X"00", X"de", 
  X"00", X"80", X"90", X"21", X"24", X"03", X"00", X"5c", 
  X"10", X"43", X"00", X"db", X"00", X"00", X"00", X"00", 
  X"ae", X"40", X"00", X"08", X"92", X"02", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"2c", X"43", X"00", X"20", 
  X"14", X"60", X"00", X"dc", X"00", X"00", X"00", X"00", 
  X"8e", X"55", X"00", X"18", X"24", X"11", X"00", X"2f", 
  X"24", X"13", X"00", X"5c", X"24", X"14", X"00", X"20", 
  X"24", X"16", X"00", X"2e", X"3c", X"17", X"bf", X"c0", 
  X"10", X"51", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"14", X"53", X"00", X"05", X"26", X"a3", X"00", X"0b", 
  X"26", X"10", X"00", X"01", X"92", X"02", X"00", X"00", 
  X"0b", X"f0", X"09", X"0c", X"00", X"00", X"00", X"00", 
  X"02", X"a0", X"10", X"21", X"a0", X"54", X"00", X"00", 
  X"24", X"42", X"00", X"01", X"14", X"43", X"ff", X"fd", 
  X"00", X"00", X"28", X"21", X"00", X"00", X"18", X"21", 
  X"24", X"04", X"00", X"08", X"00", X"00", X"40", X"21", 
  X"24", X"09", X"00", X"08", X"24", X"0a", X"00", X"22", 
  X"02", X"03", X"10", X"21", X"90", X"42", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"2c", X"46", X"00", X"21", 
  X"14", X"c0", X"00", X"21", X"24", X"63", X"00", X"01", 
  X"10", X"51", X"00", X"9c", X"00", X"00", X"00", X"00", 
  X"10", X"53", X"00", X"9a", X"00", X"00", X"00", X"00", 
  X"10", X"56", X"00", X"03", X"00", X"a4", X"30", X"2b", 
  X"14", X"c0", X"00", X"5b", X"00", X"02", X"36", X"00", 
  X"14", X"89", X"00", X"03", X"00", X"00", X"00", X"00", 
  X"10", X"56", X"00", X"0d", X"02", X"03", X"10", X"21", 
  X"24", X"02", X"00", X"06", X"8f", X"bf", X"00", X"34", 
  X"8f", X"b7", X"00", X"30", X"8f", X"b6", X"00", X"2c", 
  X"8f", X"b5", X"00", X"28", X"8f", X"b4", X"00", X"24", 
  X"8f", X"b3", X"00", X"20", X"8f", X"b2", X"00", X"1c", 
  X"8f", X"b1", X"00", X"18", X"8f", X"b0", X"00", X"14", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"38", 
  X"90", X"42", X"00", X"00", X"00", X"08", X"40", X"80", 
  X"2c", X"46", X"00", X"21", X"31", X"08", X"00", X"ff", 
  X"24", X"05", X"00", X"08", X"24", X"04", X"00", X"0b", 
  X"10", X"c0", X"ff", X"e1", X"24", X"63", X"00", X"01", 
  X"02", X"03", X"80", X"21", X"24", X"02", X"00", X"04", 
  X"10", X"a0", X"ff", X"e9", X"00", X"00", X"00", X"00", 
  X"92", X"a5", X"00", X"00", X"24", X"03", X"00", X"e5", 
  X"10", X"a3", X"00", X"a4", X"24", X"03", X"00", X"08", 
  X"10", X"83", X"00", X"a7", X"31", X"04", X"00", X"03", 
  X"24", X"03", X"00", X"01", X"10", X"83", X"00", X"aa", 
  X"31", X"08", X"00", X"0c", X"24", X"03", X"00", X"04", 
  X"11", X"03", X"00", X"94", X"00", X"00", X"00", X"00", 
  X"a2", X"a2", X"00", X"0b", X"0f", X"f0", X"08", X"99", 
  X"02", X"40", X"20", X"21", X"14", X"40", X"00", X"70", 
  X"00", X"00", X"00", X"00", X"8e", X"44", X"00", X"00", 
  X"8e", X"45", X"00", X"10", X"0f", X"f0", X"06", X"73", 
  X"00", X"00", X"00", X"00", X"14", X"40", X"00", X"6a", 
  X"00", X"00", X"00", X"00", X"8e", X"45", X"00", X"14", 
  X"00", X"00", X"00", X"00", X"90", X"a3", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"00", X"6c", 
  X"00", X"00", X"00", X"00", X"90", X"a9", X"00", X"0b", 
  X"00", X"00", X"00", X"00", X"31", X"23", X"00", X"08", 
  X"14", X"60", X"00", X"5b", X"00", X"a0", X"18", X"21", 
  X"8e", X"55", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"02", X"a0", X"20", X"21", X"24", X"a8", X"00", X"0b", 
  X"90", X"67", X"00", X"00", X"90", X"86", X"00", X"00", 
  X"24", X"63", X"00", X"01", X"14", X"e6", X"00", X"52", 
  X"24", X"84", X"00", X"01", X"14", X"68", X"ff", X"fa", 
  X"00", X"00", X"00", X"00", X"92", X"a3", X"00", X"0b", 
  X"00", X"00", X"00", X"00", X"30", X"63", X"00", X"04", 
  X"14", X"60", X"ff", X"b8", X"00", X"00", X"00", X"00", 
  X"31", X"29", X"00", X"10", X"11", X"20", X"00", X"69", 
  X"00", X"00", X"00", X"00", X"8e", X"42", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"90", X"44", X"00", X"00", 
  X"0f", X"f0", X"06", X"d3", X"00", X"00", X"00", X"00", 
  X"ae", X"42", X"00", X"08", X"92", X"02", X"00", X"00", 
  X"0b", X"f0", X"09", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"06", X"36", X"03", X"04", X"c0", X"00", X"37", 
  X"00", X"00", X"00", X"00", X"24", X"46", X"00", X"7f", 
  X"30", X"c6", X"00", X"ff", X"2c", X"c6", X"00", X"1f", 
  X"14", X"c0", X"00", X"20", X"02", X"03", X"30", X"21", 
  X"24", X"46", X"00", X"20", X"30", X"c6", X"00", X"ff", 
  X"2c", X"c6", X"00", X"1d", X"14", X"c0", X"00", X"1b", 
  X"02", X"03", X"30", X"21", X"10", X"4a", X"ff", X"9c", 
  X"26", X"e6", X"3a", X"14", X"0b", X"f0", X"09", X"99", 
  X"24", X"c6", X"00", X"01", X"10", X"47", X"ff", X"98", 
  X"24", X"c6", X"00", X"01", X"90", X"c7", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"14", X"e0", X"ff", X"fb", 
  X"00", X"00", X"00", X"00", X"24", X"46", X"ff", X"bf", 
  X"30", X"c6", X"00", X"ff", X"2c", X"c6", X"00", X"1a", 
  X"14", X"c0", X"00", X"37", X"24", X"46", X"ff", X"9f", 
  X"30", X"c6", X"00", X"ff", X"2c", X"c6", X"00", X"1a", 
  X"10", X"c0", X"00", X"05", X"02", X"a5", X"30", X"21", 
  X"24", X"42", X"ff", X"e0", X"35", X"08", X"00", X"01", 
  X"30", X"42", X"00", X"ff", X"02", X"a5", X"30", X"21", 
  X"a0", X"c2", X"00", X"00", X"0b", X"f0", X"09", X"1e", 
  X"24", X"a5", X"00", X"01", X"90", X"c6", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"24", X"c7", X"ff", X"c0", 
  X"2c", X"e7", X"00", X"3f", X"14", X"e0", X"00", X"05", 
  X"24", X"87", X"ff", X"ff", X"38", X"c7", X"00", X"80", 
  X"2c", X"e7", X"00", X"7d", X"10", X"e0", X"ff", X"7a", 
  X"24", X"87", X"ff", X"ff", X"00", X"a7", X"38", X"2b", 
  X"10", X"e0", X"ff", X"77", X"02", X"a5", X"58", X"21", 
  X"a1", X"62", X"00", X"00", X"24", X"63", X"00", X"01", 
  X"a1", X"66", X"00", X"01", X"0b", X"f0", X"09", X"1e", 
  X"24", X"a5", X"00", X"02", X"0b", X"f0", X"09", X"89", 
  X"35", X"08", X"00", X"03", X"02", X"03", X"80", X"21", 
  X"0b", X"f0", X"09", X"46", X"00", X"00", X"10", X"21", 
  X"0f", X"f0", X"08", X"42", X"02", X"40", X"20", X"21", 
  X"10", X"40", X"ff", X"92", X"00", X"00", X"00", X"00", 
  X"8e", X"43", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"90", X"64", X"00", X"0b", X"24", X"03", X"00", X"04", 
  X"14", X"43", X"ff", X"64", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"09", X"d5", X"30", X"82", X"00", X"04", 
  X"8e", X"42", X"00", X"18", X"00", X"00", X"00", X"00", 
  X"90", X"44", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"30", X"82", X"00", X"04", X"2c", X"42", X"00", X"01", 
  X"0b", X"f0", X"09", X"31", X"24", X"42", X"00", X"04", 
  X"0b", X"f0", X"09", X"a9", X"35", X"08", X"00", X"02", 
  X"26", X"10", X"00", X"01", X"ae", X"40", X"00", X"08", 
  X"92", X"02", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"2c", X"43", X"00", X"20", X"10", X"60", X"ff", X"26", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"08", X"99", 
  X"02", X"40", X"20", X"21", X"0b", X"f0", X"09", X"31", 
  X"ae", X"40", X"00", X"14", X"0b", X"f0", X"09", X"31", 
  X"24", X"02", X"00", X"05", X"34", X"42", X"00", X"08", 
  X"a2", X"a2", X"00", X"0b", X"0f", X"f0", X"08", X"99", 
  X"02", X"40", X"20", X"21", X"14", X"40", X"ff", X"dc", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"09", X"59", 
  X"00", X"00", X"00", X"00", X"24", X"03", X"00", X"05", 
  X"a2", X"a3", X"00", X"00", X"24", X"03", X"00", X"08", 
  X"14", X"83", X"ff", X"5b", X"31", X"04", X"00", X"03", 
  X"00", X"08", X"40", X"80", X"31", X"08", X"00", X"ff", 
  X"31", X"04", X"00", X"03", X"24", X"03", X"00", X"01", 
  X"14", X"83", X"ff", X"58", X"31", X"08", X"00", X"0c", 
  X"24", X"03", X"00", X"04", X"15", X"03", X"ff", X"58", 
  X"34", X"42", X"00", X"10", X"0b", X"f0", X"09", X"e8", 
  X"34", X"42", X"00", X"08", X"30", X"84", X"00", X"ff", 
  X"14", X"80", X"00", X"0d", X"24", X"02", X"00", X"0b", 
  X"3c", X"02", X"00", X"08", X"8c", X"43", X"c0", X"08", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"a0", X"60", X"00", X"00", 
  X"10", X"a0", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"a0", X"a0", X"00", X"00", X"ac", X"45", X"c0", X"08", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"27", X"bd", X"ff", X"b0", X"af", X"b2", X"00", X"40", 
  X"af", X"b0", X"00", X"38", X"af", X"bf", X"00", X"4c", 
  X"af", X"b4", X"00", X"48", X"af", X"b3", X"00", X"44", 
  X"af", X"b1", X"00", X"3c", X"00", X"80", X"80", X"21", 
  X"af", X"a5", X"00", X"54", X"10", X"80", X"00", X"21", 
  X"00", X"c0", X"90", X"21", X"ac", X"80", X"00", X"00", 
  X"27", X"a5", X"00", X"1c", X"0f", X"f0", X"06", X"e3", 
  X"27", X"a4", X"00", X"54", X"10", X"40", X"00", X"0a", 
  X"00", X"40", X"88", X"21", X"8f", X"bf", X"00", X"4c", 
  X"02", X"20", X"10", X"21", X"8f", X"b4", X"00", X"48", 
  X"8f", X"b3", X"00", X"44", X"8f", X"b2", X"00", X"40", 
  X"8f", X"b1", X"00", X"3c", X"8f", X"b0", X"00", X"38", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"50", 
  X"8f", X"a5", X"00", X"54", X"27", X"a2", X"00", X"10", 
  X"27", X"a4", X"00", X"1c", X"0f", X"f0", X"08", X"ee", 
  X"af", X"a2", X"00", X"34", X"8f", X"b3", X"00", X"30", 
  X"14", X"40", X"ff", X"f0", X"00", X"40", X"88", X"21", 
  X"12", X"60", X"00", X"29", X"00", X"00", X"00", X"00", 
  X"92", X"62", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"30", X"42", X"00", X"10", X"10", X"40", X"00", X"0d", 
  X"32", X"52", X"00", X"01", X"0b", X"f0", X"0a", X"21", 
  X"24", X"11", X"00", X"04", X"8f", X"bf", X"00", X"4c", 
  X"24", X"11", X"00", X"09", X"02", X"20", X"10", X"21", 
  X"8f", X"b4", X"00", X"48", X"8f", X"b3", X"00", X"44", 
  X"8f", X"b2", X"00", X"40", X"8f", X"b1", X"00", X"3c", 
  X"8f", X"b0", X"00", X"38", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"50", X"8f", X"b4", X"00", X"1c", 
  X"a2", X"12", X"00", X"06", X"92", X"84", X"00", X"00", 
  X"0f", X"f0", X"06", X"d3", X"02", X"60", X"28", X"21", 
  X"ae", X"02", X"00", X"10", X"92", X"65", X"00", X"1f", 
  X"92", X"63", X"00", X"1e", X"92", X"62", X"00", X"1c", 
  X"92", X"64", X"00", X"1d", X"00", X"05", X"2e", X"00", 
  X"00", X"03", X"1c", X"00", X"00", X"a3", X"18", X"25", 
  X"00", X"62", X"18", X"25", X"00", X"04", X"22", X"00", 
  X"96", X"82", X"00", X"06", X"00", X"64", X"18", X"25", 
  X"ae", X"03", X"00", X"0c", X"ae", X"00", X"00", X"08", 
  X"ae", X"00", X"00", X"18", X"ae", X"14", X"00", X"00", 
  X"0b", X"f0", X"0a", X"21", X"a6", X"02", X"00", X"04", 
  X"0b", X"f0", X"0a", X"21", X"24", X"11", X"00", X"06", 
  X"27", X"bd", X"ff", X"c0", X"af", X"b5", X"00", X"2c", 
  X"af", X"b3", X"00", X"24", X"af", X"b0", X"00", X"18", 
  X"af", X"bf", X"00", X"3c", X"af", X"be", X"00", X"38", 
  X"af", X"b7", X"00", X"34", X"af", X"b6", X"00", X"30", 
  X"af", X"b4", X"00", X"28", X"af", X"b2", X"00", X"20", 
  X"af", X"b1", X"00", X"1c", X"ac", X"e0", X"00", X"00", 
  X"00", X"e0", X"98", X"21", X"af", X"a5", X"00", X"10", 
  X"af", X"a6", X"00", X"14", X"0f", X"f0", X"06", X"57", 
  X"00", X"80", X"80", X"21", X"8f", X"a5", X"00", X"10", 
  X"8f", X"a6", X"00", X"14", X"14", X"40", X"00", X"2c", 
  X"00", X"40", X"a8", X"21", X"92", X"02", X"00", X"06", 
  X"00", X"00", X"00", X"00", X"00", X"02", X"1e", X"00", 
  X"00", X"03", X"1e", X"03", X"04", X"60", X"00", X"92", 
  X"30", X"42", X"00", X"01", X"10", X"40", X"00", X"31", 
  X"00", X"00", X"00", X"00", X"8e", X"07", X"00", X"08", 
  X"8e", X"02", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"47", X"10", X"23", X"00", X"46", X"18", X"2b", 
  X"14", X"60", X"00", X"81", X"00", X"c0", X"88", X"21", 
  X"12", X"20", X"00", X"1b", X"00", X"a0", X"90", X"21", 
  X"24", X"1e", X"02", X"00", X"26", X"17", X"00", X"1c", 
  X"30", X"e2", X"01", X"ff", X"14", X"40", X"00", X"33", 
  X"03", X"c2", X"a0", X"23", X"8e", X"04", X"00", X"00", 
  X"00", X"07", X"12", X"42", X"90", X"83", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"24", X"63", X"ff", X"ff", 
  X"00", X"43", X"18", X"24", X"30", X"63", X"00", X"ff", 
  X"10", X"60", X"00", X"41", X"00", X"00", X"00", X"00", 
  X"8e", X"02", X"00", X"14", X"8c", X"85", X"00", X"0c", 
  X"24", X"56", X"ff", X"fe", X"24", X"a2", X"ff", X"fe", 
  X"02", X"c2", X"10", X"2b", X"14", X"40", X"00", X"4c", 
  X"00", X"00", X"00", X"00", X"92", X"03", X"00", X"06", 
  X"24", X"02", X"ff", X"80", X"00", X"62", X"10", X"25", 
  X"a2", X"02", X"00", X"06", X"24", X"15", X"00", X"02", 
  X"8f", X"bf", X"00", X"3c", X"02", X"a0", X"10", X"21", 
  X"8f", X"be", X"00", X"38", X"8f", X"b7", X"00", X"34", 
  X"8f", X"b6", X"00", X"30", X"8f", X"b5", X"00", X"2c", 
  X"8f", X"b4", X"00", X"28", X"8f", X"b3", X"00", X"24", 
  X"8f", X"b2", X"00", X"20", X"8f", X"b1", X"00", X"1c", 
  X"8f", X"b0", X"00", X"18", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"40", X"0b", X"f0", X"0a", X"9e", 
  X"24", X"15", X"00", X"07", X"8e", X"02", X"00", X"18", 
  X"00", X"00", X"00", X"00", X"10", X"56", X"00", X"07", 
  X"02", X"e0", X"28", X"21", X"90", X"84", X"00", X"01", 
  X"02", X"c0", X"30", X"21", X"0f", X"f0", X"05", X"96", 
  X"24", X"07", X"00", X"01", X"14", X"40", X"00", X"56", 
  X"00", X"00", X"00", X"00", X"8e", X"07", X"00", X"08", 
  X"ae", X"16", X"00", X"18", X"30", X"e2", X"01", X"ff", 
  X"03", X"c2", X"a0", X"23", X"02", X"34", X"18", X"2b", 
  X"10", X"60", X"00", X"02", X"00", X"00", X"00", X"00", 
  X"02", X"20", X"a0", X"21", X"12", X"80", X"00", X"09", 
  X"02", X"e2", X"10", X"21", X"00", X"54", X"28", X"21", 
  X"02", X"40", X"18", X"21", X"90", X"44", X"00", X"00", 
  X"24", X"42", X"00", X"01", X"a0", X"64", X"00", X"00", 
  X"14", X"45", X"ff", X"fc", X"24", X"63", X"00", X"01", 
  X"8e", X"07", X"00", X"08", X"8e", X"62", X"00", X"00", 
  X"00", X"f4", X"38", X"21", X"00", X"54", X"10", X"21", 
  X"02", X"34", X"88", X"23", X"ae", X"07", X"00", X"08", 
  X"12", X"20", X"ff", X"cf", X"ae", X"62", X"00", X"00", 
  X"0b", X"f0", X"0a", X"86", X"02", X"54", X"90", X"21", 
  X"14", X"e0", X"00", X"31", X"00", X"00", X"00", X"00", 
  X"8e", X"02", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"2c", X"44", X"00", X"02", X"14", X"80", X"00", X"3a", 
  X"00", X"00", X"00", X"00", X"24", X"04", X"ff", X"ff", 
  X"10", X"44", X"00", X"31", X"24", X"56", X"ff", X"fe", 
  X"8e", X"04", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"8c", X"85", X"00", X"0c", X"ae", X"02", X"00", X"14", 
  X"24", X"a2", X"ff", X"fe", X"02", X"c2", X"10", X"2b", 
  X"10", X"40", X"ff", X"b6", X"00", X"00", X"00", X"00", 
  X"90", X"82", X"00", X"02", X"8c", X"85", X"00", X"1c", 
  X"02", X"c2", X"00", X"18", X"00", X"00", X"b0", X"12", 
  X"02", X"c5", X"b0", X"21", X"12", X"c0", X"ff", X"af", 
  X"00", X"11", X"a2", X"42", X"12", X"80", X"ff", X"c1", 
  X"02", X"c3", X"b0", X"21", X"00", X"74", X"28", X"21", 
  X"00", X"45", X"28", X"2b", X"10", X"a0", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"00", X"43", X"a0", X"23", 
  X"90", X"84", X"00", X"01", X"02", X"40", X"28", X"21", 
  X"02", X"c0", X"30", X"21", X"0f", X"f0", X"05", X"96", 
  X"32", X"87", X"00", X"ff", X"14", X"40", X"00", X"04", 
  X"00", X"14", X"a2", X"40", X"8e", X"07", X"00", X"08", 
  X"0b", X"f0", X"0a", X"c9", X"00", X"00", X"00", X"00", 
  X"92", X"03", X"00", X"06", X"24", X"02", X"ff", X"80", 
  X"00", X"62", X"10", X"25", X"a2", X"02", X"00", X"06", 
  X"0b", X"f0", X"0a", X"9e", X"24", X"15", X"00", X"01", 
  X"0b", X"f0", X"0a", X"82", X"00", X"40", X"88", X"21", 
  X"8e", X"05", X"00", X"14", X"0f", X"f0", X"07", X"da", 
  X"af", X"a3", X"00", X"10", X"8f", X"a3", X"00", X"10", 
  X"0b", X"f0", X"0a", X"d7", X"2c", X"44", X"00", X"02", 
  X"0b", X"f0", X"0a", X"9e", X"24", X"15", X"00", X"02", 
  X"92", X"03", X"00", X"06", X"24", X"02", X"ff", X"80", 
  X"00", X"62", X"10", X"25", X"a2", X"02", X"00", X"06", 
  X"0b", X"f0", X"0a", X"9e", X"24", X"15", X"00", X"01", 
  X"92", X"03", X"00", X"06", X"24", X"02", X"ff", X"80", 
  X"00", X"62", X"10", X"25", X"a2", X"02", X"00", X"06", 
  X"0b", X"f0", X"0a", X"9e", X"24", X"15", X"00", X"02", 
  X"27", X"bd", X"ff", X"e8", X"af", X"b0", X"00", X"10", 
  X"af", X"bf", X"00", X"14", X"0f", X"f0", X"06", X"57", 
  X"00", X"80", X"80", X"21", X"14", X"40", X"00", X"02", 
  X"00", X"00", X"00", X"00", X"ae", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"18", 
  X"27", X"bd", X"ff", X"c8", X"af", X"b1", X"00", X"20", 
  X"af", X"b0", X"00", X"1c", X"af", X"a5", X"00", X"10", 
  X"af", X"bf", X"00", X"34", X"af", X"b5", X"00", X"30", 
  X"af", X"b4", X"00", X"2c", X"af", X"b3", X"00", X"28", 
  X"af", X"b2", X"00", X"24", X"0f", X"f0", X"06", X"57", 
  X"00", X"80", X"80", X"21", X"8f", X"a5", X"00", X"10", 
  X"14", X"40", X"00", X"49", X"00", X"40", X"88", X"21", 
  X"82", X"02", X"00", X"06", X"00", X"00", X"00", X"00", 
  X"04", X"40", X"00", X"6a", X"00", X"00", X"00", X"00", 
  X"8e", X"02", X"00", X"0c", X"00", X"00", X"00", X"00", 
  X"00", X"45", X"18", X"2b", X"14", X"60", X"00", X"4a", 
  X"00", X"a0", X"90", X"21", X"8e", X"02", X"00", X"08", 
  X"12", X"40", X"00", X"3d", X"ae", X"00", X"00", X"08", 
  X"8e", X"04", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"90", X"93", X"00", X"02", X"10", X"40", X"00", X"48", 
  X"00", X"13", X"9a", X"40", X"26", X"43", X"ff", X"ff", 
  X"16", X"60", X"00", X"02", X"00", X"73", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"24", X"42", X"ff", X"ff", 
  X"00", X"00", X"18", X"12", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"16", X"60", X"00", X"02", 
  X"00", X"53", X"00", X"1b", X"00", X"07", X"00", X"0d", 
  X"00", X"00", X"28", X"12", X"00", X"65", X"18", X"2b", 
  X"14", X"60", X"00", X"39", X"00", X"13", X"18", X"23", 
  X"00", X"62", X"10", X"24", X"ae", X"02", X"00", X"08", 
  X"02", X"42", X"90", X"23", X"8e", X"02", X"00", X"14", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"36", 
  X"00", X"00", X"00", X"00", X"02", X"72", X"18", X"2b", 
  X"10", X"60", X"00", X"4c", X"00", X"13", X"a8", X"23", 
  X"02", X"53", X"90", X"23", X"0b", X"f0", X"0b", X"6e", 
  X"24", X"14", X"ff", X"ff", X"14", X"80", X"00", X"41", 
  X"00", X"00", X"00", X"00", X"8e", X"04", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"8c", X"86", X"00", X"0c", 
  X"00", X"00", X"00", X"00", X"00", X"46", X"30", X"2b", 
  X"10", X"c0", X"00", X"3a", X"00", X"00", X"00", X"00", 
  X"8e", X"06", X"00", X"08", X"ae", X"02", X"00", X"14", 
  X"02", X"66", X"30", X"21", X"10", X"60", X"00", X"3d", 
  X"ae", X"06", X"00", X"08", X"00", X"a0", X"90", X"21", 
  X"0f", X"f0", X"07", X"da", X"00", X"40", X"28", X"21", 
  X"02", X"55", X"28", X"21", X"00", X"b3", X"18", X"21", 
  X"2c", X"44", X"00", X"02", X"14", X"54", X"ff", X"eb", 
  X"02", X"63", X"18", X"2b", X"92", X"03", X"00", X"06", 
  X"24", X"02", X"ff", X"80", X"00", X"62", X"10", X"25", 
  X"a2", X"02", X"00", X"06", X"24", X"11", X"00", X"01", 
  X"8f", X"bf", X"00", X"34", X"02", X"20", X"10", X"21", 
  X"8f", X"b5", X"00", X"30", X"8f", X"b4", X"00", X"2c", 
  X"8f", X"b3", X"00", X"28", X"8f", X"b2", X"00", X"24", 
  X"8f", X"b1", X"00", X"20", X"8f", X"b0", X"00", X"1c", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"38", 
  X"00", X"40", X"90", X"21", X"8e", X"02", X"00", X"08", 
  X"12", X"40", X"ff", X"f3", X"ae", X"00", X"00", X"08", 
  X"0b", X"f0", X"0b", X"3e", X"00", X"00", X"00", X"00", 
  X"8e", X"02", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"ff", X"cc", X"ae", X"02", X"00", X"14", 
  X"8e", X"03", X"00", X"08", X"00", X"00", X"90", X"21", 
  X"30", X"63", X"01", X"ff", X"10", X"60", X"ff", X"e8", 
  X"00", X"00", X"00", X"00", X"8e", X"02", X"00", X"18", 
  X"00", X"00", X"00", X"00", X"10", X"52", X"ff", X"e4", 
  X"02", X"40", X"30", X"21", X"90", X"84", X"00", X"01", 
  X"26", X"05", X"00", X"1c", X"0f", X"f0", X"05", X"96", 
  X"24", X"07", X"00", X"01", X"14", X"40", X"ff", X"d9", 
  X"00", X"00", X"00", X"00", X"0b", X"f0", X"0b", X"7a", 
  X"ae", X"12", X"00", X"18", X"0b", X"f0", X"0b", X"7a", 
  X"24", X"11", X"00", X"02", X"92", X"03", X"00", X"06", 
  X"24", X"02", X"ff", X"80", X"00", X"62", X"10", X"25", 
  X"a2", X"02", X"00", X"06", X"0b", X"f0", X"0b", X"7a", 
  X"24", X"11", X"00", X"02", X"8e", X"06", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"00", X"d2", X"18", X"21", 
  X"32", X"45", X"01", X"ff", X"10", X"a0", X"00", X"10", 
  X"ae", X"03", X"00", X"08", X"8c", X"85", X"00", X"0c", 
  X"24", X"42", X"ff", X"fe", X"24", X"a5", X"ff", X"fe", 
  X"00", X"45", X"28", X"2b", X"10", X"a0", X"ff", X"ef", 
  X"00", X"00", X"00", X"00", X"90", X"86", X"00", X"02", 
  X"8c", X"85", X"00", X"1c", X"00", X"46", X"00", X"18", 
  X"00", X"00", X"10", X"12", X"00", X"45", X"28", X"21", 
  X"10", X"a0", X"ff", X"e8", X"00", X"12", X"92", X"42", 
  X"0b", X"f0", X"0b", X"90", X"00", X"b2", X"90", X"21", 
  X"0b", X"f0", X"0b", X"90", X"00", X"00", X"90", X"21", 
  X"27", X"bd", X"ff", X"d0", X"af", X"b0", X"00", X"24", 
  X"af", X"bf", X"00", X"2c", X"af", X"b1", X"00", X"28", 
  X"00", X"80", X"80", X"21", X"10", X"80", X"00", X"2f", 
  X"af", X"a5", X"00", X"34", X"27", X"a4", X"00", X"34", 
  X"0f", X"f0", X"06", X"e3", X"02", X"00", X"28", X"21", 
  X"8e", X"11", X"00", X"00", X"10", X"40", X"00", X"07", 
  X"00", X"00", X"00", X"00", X"8f", X"bf", X"00", X"2c", 
  X"ae", X"00", X"00", X"00", X"8f", X"b1", X"00", X"28", 
  X"8f", X"b0", X"00", X"24", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"27", X"a2", X"00", X"10", 
  X"8f", X"a5", X"00", X"34", X"ae", X"02", X"00", X"18", 
  X"0f", X"f0", X"08", X"ee", X"02", X"00", X"20", X"21", 
  X"14", X"40", X"00", X"13", X"24", X"03", X"00", X"04", 
  X"8e", X"05", X"00", X"14", X"00", X"00", X"00", X"00", 
  X"10", X"a0", X"00", X"0a", X"00", X"00", X"00", X"00", 
  X"90", X"a2", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"30", X"42", X"00", X"10", X"10", X"40", X"ff", X"eb", 
  X"24", X"02", X"00", X"05", X"92", X"24", X"00", X"00", 
  X"0f", X"f0", X"06", X"d3", X"00", X"00", X"00", X"00", 
  X"ae", X"02", X"00", X"08", X"96", X"22", X"00", X"06", 
  X"02", X"00", X"20", X"21", X"0f", X"f0", X"08", X"99", 
  X"a6", X"02", X"00", X"04", X"24", X"03", X"00", X"04", 
  X"10", X"43", X"00", X"0e", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"ff", X"de", X"00", X"00", X"00", X"00", 
  X"8f", X"bf", X"00", X"2c", X"8f", X"b1", X"00", X"28", 
  X"8f", X"b0", X"00", X"24", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"8f", X"bf", X"00", X"2c", 
  X"24", X"02", X"00", X"09", X"8f", X"b1", X"00", X"28", 
  X"8f", X"b0", X"00", X"24", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"30", X"0b", X"f0", X"0b", X"cb", 
  X"24", X"02", X"00", X"05", X"27", X"bd", X"ff", X"c8", 
  X"af", X"b4", X"00", X"30", X"af", X"b2", X"00", X"28", 
  X"af", X"b0", X"00", X"20", X"af", X"bf", X"00", X"34", 
  X"af", X"b3", X"00", X"2c", X"af", X"b1", X"00", X"24", 
  X"00", X"80", X"80", X"21", X"0f", X"f0", X"06", X"57", 
  X"00", X"a0", X"a0", X"21", X"14", X"40", X"00", X"2e", 
  X"00", X"40", X"90", X"21", X"12", X"80", X"00", X"88", 
  X"27", X"a2", X"00", X"10", X"ae", X"02", X"00", X"18", 
  X"24", X"11", X"00", X"e5", X"24", X"02", X"00", X"04", 
  X"24", X"13", X"00", X"2e", X"8e", X"03", X"00", X"10", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"00", X"37", 
  X"00", X"60", X"28", X"21", X"8e", X"04", X"00", X"00", 
  X"0f", X"f0", X"06", X"73", X"00", X"00", X"00", X"00", 
  X"14", X"40", X"00", X"14", X"02", X"00", X"20", X"21", 
  X"8e", X"03", X"00", X"14", X"00", X"00", X"00", X"00", 
  X"90", X"62", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"10", X"40", X"00", X"6e", X"00", X"00", X"00", X"00", 
  X"10", X"51", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"10", X"53", X"00", X"06", X"00", X"00", X"00", X"00", 
  X"90", X"62", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"30", X"42", X"00", X"08", X"10", X"40", X"00", X"69", 
  X"00", X"00", X"00", X"00", X"0f", X"f0", X"08", X"42", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"ff", X"e5", 
  X"00", X"00", X"00", X"00", X"24", X"03", X"00", X"04", 
  X"14", X"43", X"00", X"12", X"ae", X"00", X"00", X"10", 
  X"26", X"82", X"00", X"09", X"a0", X"40", X"00", X"00", 
  X"0f", X"f0", X"08", X"42", X"02", X"00", X"20", X"21", 
  X"24", X"03", X"00", X"04", X"14", X"43", X"00", X"0b", 
  X"00", X"00", X"00", X"00", X"ae", X"00", X"00", X"10", 
  X"8f", X"bf", X"00", X"34", X"02", X"40", X"10", X"21", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"8f", X"bf", X"00", X"34", 
  X"00", X"40", X"90", X"21", X"02", X"40", X"10", X"21", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"14", X"40", X"ff", X"e1", 
  X"00", X"00", X"00", X"00", X"10", X"60", X"00", X"4a", 
  X"26", X"84", X"00", X"09", X"8e", X"05", X"00", X"14", 
  X"00", X"00", X"18", X"21", X"24", X"06", X"00", X"20", 
  X"24", X"08", X"00", X"05", X"0b", X"f0", X"0c", X"54", 
  X"24", X"07", X"00", X"08", X"a0", X"82", X"00", X"00", 
  X"10", X"67", X"00", X"0c", X"24", X"84", X"00", X"01", 
  X"00", X"a3", X"10", X"21", X"90", X"42", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"46", X"00", X"07", 
  X"24", X"63", X"00", X"01", X"14", X"48", X"ff", X"f7", 
  X"00", X"00", X"00", X"00", X"24", X"02", X"00", X"e5", 
  X"a0", X"82", X"00", X"00", X"14", X"67", X"ff", X"f6", 
  X"24", X"84", X"00", X"01", X"90", X"a3", X"00", X"08", 
  X"24", X"02", X"00", X"20", X"10", X"62", X"00", X"29", 
  X"00", X"a0", X"18", X"21", X"24", X"02", X"00", X"2e", 
  X"a0", X"82", X"00", X"00", X"24", X"82", X"00", X"01", 
  X"24", X"07", X"00", X"20", X"24", X"84", X"00", X"04", 
  X"90", X"66", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"10", X"c7", X"00", X"05", X"24", X"63", X"00", X"01", 
  X"a0", X"46", X"00", X"00", X"24", X"42", X"00", X"01", 
  X"14", X"44", X"ff", X"f9", X"00", X"00", X"00", X"00", 
  X"90", X"a3", X"00", X"0b", X"00", X"00", X"00", X"00", 
  X"a2", X"83", X"00", X"08", X"90", X"a7", X"00", X"1f", 
  X"90", X"a3", X"00", X"1e", X"90", X"a6", X"00", X"1c", 
  X"90", X"a4", X"00", X"1d", X"00", X"07", X"3e", X"00", 
  X"00", X"03", X"1c", X"00", X"00", X"e3", X"18", X"25", 
  X"00", X"04", X"22", X"00", X"00", X"66", X"18", X"25", 
  X"00", X"64", X"18", X"25", X"ae", X"83", X"00", X"00", 
  X"90", X"a3", X"00", X"19", X"90", X"a4", X"00", X"18", 
  X"00", X"03", X"1a", X"00", X"00", X"64", X"18", X"25", 
  X"a6", X"83", X"00", X"04", X"90", X"a3", X"00", X"17", 
  X"90", X"a4", X"00", X"16", X"00", X"03", X"1a", X"00", 
  X"00", X"64", X"18", X"25", X"0b", X"f0", X"0c", X"2d", 
  X"a6", X"83", X"00", X"06", X"0b", X"f0", X"0c", X"29", 
  X"24", X"02", X"00", X"04", X"0b", X"f0", X"0c", X"70", 
  X"00", X"80", X"10", X"21", X"8e", X"03", X"00", X"10", 
  X"0b", X"f0", X"0c", X"49", X"00", X"00", X"00", X"00", 
  X"0f", X"f0", X"08", X"99", X"02", X"00", X"20", X"21", 
  X"0b", X"f0", X"0c", X"34", X"00", X"40", X"90", X"21", 
  X"0b", X"f0", X"0c", X"2d", X"00", X"80", X"10", X"21", 
  X"10", X"80", X"00", X"09", X"00", X"00", X"00", X"00", 
  X"8c", X"82", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"a0", X"45", X"00", X"00", X"8c", X"82", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"24", X"42", X"00", X"01", 
  X"03", X"e0", X"00", X"08", X"ac", X"82", X"00", X"00", 
  X"0b", X"f0", X"0e", X"2a", X"00", X"a0", X"20", X"21", 
  X"27", X"bd", X"ff", X"d8", X"af", X"b2", X"00", X"18", 
  X"af", X"b1", X"00", X"14", X"af", X"b0", X"00", X"10", 
  X"af", X"bf", X"00", X"24", X"af", X"b4", X"00", X"20", 
  X"af", X"b3", X"00", X"1c", X"00", X"c0", X"90", X"21", 
  X"00", X"80", X"88", X"21", X"18", X"c0", X"00", X"32", 
  X"00", X"a0", X"80", X"21", X"90", X"a2", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"40", X"00", X"3d", 
  X"00", X"a0", X"10", X"21", X"00", X"00", X"18", X"21", 
  X"24", X"42", X"00", X"01", X"90", X"44", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"14", X"80", X"ff", X"fc", 
  X"24", X"63", X"00", X"01", X"00", X"72", X"10", X"2a", 
  X"14", X"40", X"00", X"02", X"02", X"43", X"90", X"23", 
  X"00", X"00", X"90", X"21", X"30", X"e2", X"00", X"02", 
  X"10", X"40", X"00", X"22", X"30", X"e7", X"00", X"01", 
  X"10", X"e0", X"00", X"22", X"24", X"14", X"00", X"30", 
  X"00", X"00", X"98", X"21", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"a0", X"00", X"08", 
  X"00", X"00", X"00", X"00", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"0c", X"96", X"26", X"10", X"00", X"01", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"fa", X"26", X"73", X"00", X"01", 
  X"1a", X"40", X"00", X"08", X"02", X"40", X"80", X"21", 
  X"26", X"10", X"ff", X"ff", X"02", X"20", X"20", X"21", 
  X"0f", X"f0", X"0c", X"96", X"02", X"80", X"28", X"21", 
  X"16", X"00", X"ff", X"fc", X"26", X"10", X"ff", X"ff", 
  X"02", X"72", X"98", X"21", X"8f", X"bf", X"00", X"24", 
  X"02", X"60", X"10", X"21", X"8f", X"b4", X"00", X"20", 
  X"8f", X"b3", X"00", X"1c", X"8f", X"b2", X"00", X"18", 
  X"8f", X"b1", X"00", X"14", X"8f", X"b0", X"00", X"10", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"28", 
  X"30", X"e7", X"00", X"01", X"14", X"e0", X"ff", X"e0", 
  X"24", X"14", X"00", X"20", X"1a", X"40", X"ff", X"de", 
  X"02", X"40", X"98", X"21", X"26", X"73", X"ff", X"ff", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"0c", X"96", 
  X"02", X"80", X"28", X"21", X"16", X"60", X"ff", X"fc", 
  X"26", X"73", X"ff", X"ff", X"26", X"73", X"00", X"01", 
  X"02", X"40", X"98", X"21", X"0b", X"f0", X"0c", X"c1", 
  X"00", X"00", X"90", X"21", X"00", X"00", X"18", X"21", 
  X"0b", X"f0", X"0c", X"bb", X"02", X"43", X"90", X"23", 
  X"27", X"bd", X"ff", X"c8", X"af", X"b4", X"00", X"30", 
  X"af", X"b2", X"00", X"28", X"af", X"b1", X"00", X"24", 
  X"af", X"bf", X"00", X"34", X"af", X"b3", X"00", X"2c", 
  X"af", X"b0", X"00", X"20", X"00", X"a0", X"10", X"21", 
  X"8f", X"b4", X"00", X"48", X"8f", X"b2", X"00", X"4c", 
  X"10", X"a0", X"00", X"3f", X"00", X"80", X"88", X"21", 
  X"14", X"e0", X"00", X"31", X"24", X"03", X"00", X"0a", 
  X"00", X"00", X"38", X"21", X"10", X"40", X"00", X"49", 
  X"a3", X"a0", X"00", X"1b", X"8f", X"a5", X"00", X"50", 
  X"27", X"b3", X"00", X"1b", X"24", X"a5", X"ff", X"c6", 
  X"14", X"c0", X"00", X"02", X"00", X"46", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"00", X"00", X"18", X"10", 
  X"28", X"64", X"00", X"0a", X"00", X"00", X"00", X"00", 
  X"14", X"c0", X"00", X"02", X"00", X"46", X"00", X"1b", 
  X"00", X"07", X"00", X"0d", X"00", X"00", X"10", X"12", 
  X"14", X"80", X"00", X"02", X"26", X"73", X"ff", X"ff", 
  X"00", X"65", X"18", X"21", X"24", X"63", X"00", X"30", 
  X"14", X"40", X"ff", X"f1", X"a2", X"63", X"00", X"00", 
  X"14", X"e0", X"00", X"10", X"00", X"00", X"00", X"00", 
  X"00", X"00", X"80", X"21", X"02", X"20", X"20", X"21", 
  X"02", X"60", X"28", X"21", X"02", X"80", X"30", X"21", 
  X"0f", X"f0", X"0c", X"a2", X"02", X"40", X"38", X"21", 
  X"8f", X"bf", X"00", X"34", X"00", X"50", X"10", X"21", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"12", X"80", X"00", X"0f", 
  X"32", X"42", X"00", X"02", X"10", X"40", X"00", X"0d", 
  X"02", X"20", X"20", X"21", X"0f", X"f0", X"0c", X"96", 
  X"24", X"05", X"00", X"2d", X"26", X"94", X"ff", X"ff", 
  X"0b", X"f0", X"0d", X"17", X"24", X"10", X"00", X"01", 
  X"14", X"c3", X"ff", X"d0", X"00", X"00", X"38", X"21", 
  X"04", X"a1", X"ff", X"ce", X"00", X"00", X"00", X"00", 
  X"00", X"05", X"10", X"23", X"0b", X"f0", X"0c", X"ff", 
  X"24", X"07", X"00", X"01", X"26", X"73", X"ff", X"ff", 
  X"24", X"02", X"00", X"2d", X"a2", X"62", X"00", X"00", 
  X"0b", X"f0", X"0d", X"17", X"00", X"00", X"80", X"21", 
  X"27", X"a5", X"00", X"10", X"02", X"80", X"30", X"21", 
  X"02", X"40", X"38", X"21", X"24", X"02", X"00", X"30", 
  X"a3", X"a2", X"00", X"10", X"0f", X"f0", X"0c", X"a2", 
  X"a3", X"a0", X"00", X"11", X"8f", X"bf", X"00", X"34", 
  X"8f", X"b4", X"00", X"30", X"8f", X"b3", X"00", X"2c", 
  X"8f", X"b2", X"00", X"28", X"8f", X"b1", X"00", X"24", 
  X"8f", X"b0", X"00", X"20", X"03", X"e0", X"00", X"08", 
  X"27", X"bd", X"00", X"38", X"10", X"e0", X"ff", X"cc", 
  X"27", X"b3", X"00", X"1b", X"0b", X"f0", X"0d", X"25", 
  X"00", X"00", X"00", X"00", X"27", X"bd", X"ff", X"b8", 
  X"af", X"b4", X"00", X"38", X"af", X"b0", X"00", X"28", 
  X"af", X"bf", X"00", X"44", X"af", X"b6", X"00", X"40", 
  X"af", X"b5", X"00", X"3c", X"af", X"b3", X"00", X"34", 
  X"af", X"b2", X"00", X"30", X"af", X"b1", X"00", X"2c", 
  X"00", X"a0", X"80", X"21", X"90", X"a5", X"00", X"00", 
  X"00", X"80", X"a0", X"21", X"10", X"a0", X"00", X"a0", 
  X"af", X"a6", X"00", X"50", X"00", X"00", X"90", X"21", 
  X"24", X"13", X"00", X"25", X"24", X"15", X"00", X"2d", 
  X"24", X"11", X"00", X"30", X"3c", X"16", X"bf", X"c0", 
  X"14", X"b3", X"00", X"53", X"00", X"00", X"00", X"00", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"a0", X"00", X"3e", 
  X"00", X"00", X"00", X"00", X"10", X"b3", X"00", X"4c", 
  X"00", X"00", X"00", X"00", X"10", X"b5", X"00", X"54", 
  X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"21", 
  X"14", X"b1", X"00", X"07", X"24", X"a2", X"ff", X"d0", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"10", X"b1", X"ff", X"fc", 
  X"34", X"63", X"00", X"02", X"24", X"a2", X"ff", X"d0", 
  X"30", X"42", X"00", X"ff", X"2c", X"42", X"00", X"0a", 
  X"10", X"40", X"00", X"0d", X"00", X"00", X"10", X"21", 
  X"00", X"02", X"20", X"40", X"00", X"02", X"10", X"c0", 
  X"00", X"82", X"10", X"21", X"26", X"10", X"00", X"01", 
  X"00", X"45", X"10", X"21", X"92", X"05", X"00", X"00", 
  X"00", X"00", X"00", X"00", X"24", X"a4", X"ff", X"d0", 
  X"30", X"84", X"00", X"ff", X"2c", X"84", X"00", X"0a", 
  X"14", X"80", X"ff", X"f5", X"24", X"42", X"ff", X"d0", 
  X"24", X"04", X"00", X"73", X"10", X"a4", X"00", X"3c", 
  X"24", X"04", X"00", X"64", X"10", X"a4", X"00", X"46", 
  X"02", X"80", X"20", X"21", X"24", X"04", X"00", X"78", 
  X"10", X"a4", X"00", X"51", X"02", X"80", X"20", X"21", 
  X"24", X"04", X"00", X"58", X"10", X"a4", X"00", X"55", 
  X"02", X"80", X"20", X"21", X"24", X"04", X"00", X"75", 
  X"10", X"a4", X"00", X"60", X"02", X"80", X"20", X"21", 
  X"24", X"04", X"00", X"63", X"14", X"a4", X"00", X"24", 
  X"26", X"10", X"00", X"01", X"8f", X"a9", X"00", X"50", 
  X"27", X"a5", X"00", X"20", X"8d", X"28", X"00", X"00", 
  X"02", X"80", X"20", X"21", X"25", X"29", X"00", X"04", 
  X"00", X"40", X"30", X"21", X"00", X"60", X"38", X"21", 
  X"af", X"a9", X"00", X"50", X"a3", X"a8", X"00", X"20", 
  X"0f", X"f0", X"0c", X"a2", X"a3", X"a0", X"00", X"21", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"bd", X"02", X"42", X"90", X"21", 
  X"12", X"80", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"8e", X"82", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"a0", X"40", X"00", X"00", X"8f", X"bf", X"00", X"44", 
  X"02", X"40", X"10", X"21", X"8f", X"b6", X"00", X"40", 
  X"8f", X"b5", X"00", X"3c", X"8f", X"b4", X"00", X"38", 
  X"8f", X"b3", X"00", X"34", X"8f", X"b2", X"00", X"30", 
  X"8f", X"b1", X"00", X"2c", X"8f", X"b0", X"00", X"28", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"48", 
  X"0f", X"f0", X"0c", X"96", X"02", X"80", X"20", X"21", 
  X"26", X"52", X"00", X"01", X"26", X"10", X"00", X"01", 
  X"92", X"05", X"00", X"00", X"00", X"00", X"00", X"00", 
  X"14", X"a0", X"ff", X"a5", X"00", X"00", X"00", X"00", 
  X"0b", X"f0", X"0d", X"a4", X"00", X"00", X"00", X"00", 
  X"26", X"10", X"00", X"01", X"92", X"05", X"00", X"00", 
  X"0b", X"f0", X"0d", X"6c", X"24", X"03", X"00", X"01", 
  X"8f", X"a4", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8c", X"85", X"00", X"00", X"24", X"84", X"00", X"04", 
  X"10", X"a0", X"00", X"31", X"af", X"a4", X"00", X"50", 
  X"02", X"80", X"20", X"21", X"00", X"40", X"30", X"21", 
  X"0f", X"f0", X"0c", X"a2", X"00", X"60", X"38", X"21", 
  X"0b", X"f0", X"0d", X"b7", X"02", X"42", X"90", X"21", 
  X"8f", X"a8", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8d", X"05", X"00", X"00", X"24", X"06", X"00", X"0a", 
  X"25", X"08", X"00", X"04", X"24", X"07", X"00", X"01", 
  X"af", X"a2", X"00", X"10", X"24", X"02", X"00", X"61", 
  X"af", X"a8", X"00", X"50", X"af", X"a3", X"00", X"14", 
  X"0f", X"f0", X"0c", X"f0", X"af", X"a2", X"00", X"18", 
  X"0b", X"f0", X"0d", X"b7", X"02", X"42", X"90", X"21", 
  X"8f", X"a8", X"00", X"50", X"00", X"00", X"00", X"00", 
  X"8d", X"05", X"00", X"00", X"24", X"06", X"00", X"10", 
  X"25", X"08", X"00", X"04", X"0b", X"f0", X"0d", X"d4", 
  X"00", X"00", X"38", X"21", X"8f", X"a8", X"00", X"50", 
  X"00", X"00", X"00", X"00", X"8d", X"05", X"00", X"00", 
  X"24", X"06", X"00", X"10", X"25", X"08", X"00", X"04", 
  X"af", X"a2", X"00", X"10", X"00", X"00", X"38", X"21", 
  X"24", X"02", X"00", X"41", X"af", X"a8", X"00", X"50", 
  X"af", X"a3", X"00", X"14", X"0f", X"f0", X"0c", X"f0", 
  X"af", X"a2", X"00", X"18", X"0b", X"f0", X"0d", X"b7", 
  X"02", X"42", X"90", X"21", X"8f", X"a8", X"00", X"50", 
  X"00", X"00", X"00", X"00", X"8d", X"05", X"00", X"00", 
  X"24", X"06", X"00", X"0a", X"25", X"08", X"00", X"04", 
  X"0b", X"f0", X"0d", X"d4", X"00", X"00", X"38", X"21", 
  X"0b", X"f0", X"0d", X"c8", X"26", X"c5", X"3a", X"24", 
  X"0b", X"f0", X"0d", X"a4", X"00", X"00", X"90", X"21", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"24", 
  X"00", X"80", X"18", X"21", X"af", X"a5", X"00", X"24", 
  X"af", X"a6", X"00", X"28", X"00", X"00", X"20", X"21", 
  X"00", X"60", X"28", X"21", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"0d", X"4d", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"28", 
  X"af", X"a4", X"00", X"20", X"af", X"a6", X"00", X"28", 
  X"27", X"a4", X"00", X"20", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"0d", X"4d", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"27", X"bd", X"ff", X"e0", X"27", X"a2", X"00", X"2c", 
  X"af", X"a4", X"00", X"20", X"00", X"c0", X"28", X"21", 
  X"27", X"a4", X"00", X"20", X"00", X"40", X"30", X"21", 
  X"af", X"bf", X"00", X"1c", X"af", X"a7", X"00", X"2c", 
  X"0f", X"f0", X"0d", X"4d", X"af", X"a2", X"00", X"10", 
  X"8f", X"bf", X"00", X"1c", X"00", X"00", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"27", X"bd", X"00", X"20", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"10", X"21", 
  X"00", X"80", X"10", X"21", X"3c", X"05", X"20", X"00", 
  X"8c", X"a3", X"00", X"04", X"00", X"00", X"00", X"00", 
  X"30", X"63", X"00", X"01", X"10", X"60", X"ff", X"fc", 
  X"3c", X"03", X"20", X"00", X"ac", X"62", X"00", X"00", 
  X"03", X"e0", X"00", X"08", X"00", X"00", X"00", X"00", 
  X"3c", X"03", X"20", X"00", X"8c", X"62", X"00", X"04", 
  X"00", X"00", X"00", X"00", X"30", X"42", X"00", X"02", 
  X"10", X"40", X"ff", X"fc", X"3c", X"02", X"20", X"00", 
  X"8c", X"42", X"00", X"00", X"03", X"e0", X"00", X"08", 
  X"30", X"42", X"00", X"ff", X"44", X"69", X"73", X"6b", 
  X"20", X"61", X"62", X"73", X"65", X"6e", X"74", X"2e", 
  X"00", X"00", X"00", X"00", X"4c", X"6f", X"77", X"20", 
  X"6c", X"65", X"76", X"65", X"6c", X"20", X"64", X"69", 
  X"73", X"6b", X"20", X"69", X"2f", X"6f", X"20", X"65", 
  X"72", X"72", X"6f", X"72", X"2e", X"00", X"00", X"00", 
  X"4e", X"6f", X"20", X"76", X"61", X"6c", X"69", X"64", 
  X"20", X"66", X"69", X"6c", X"65", X"73", X"79", X"73", 
  X"74", X"65", X"6d", X"20", X"69", X"6e", X"20", X"64", 
  X"72", X"69", X"76", X"65", X"2e", X"00", X"00", X"00", 
  X"46", X"69", X"6c", X"65", X"20", X"6e", X"6f", X"74", 
  X"20", X"66", X"6f", X"75", X"6e", X"64", X"2e", X"00", 
  X"46", X"61", X"69", X"6c", X"65", X"64", X"20", X"77", 
  X"69", X"74", X"68", X"20", X"72", X"63", X"3d", X"25", 
  X"75", X"2e", X"00", X"00", X"49", X"4f", X"4e", X"20", 
  X"53", X"44", X"20", X"6c", X"6f", X"61", X"64", X"65", 
  X"72", X"20", X"2d", X"2d", X"20", X"4e", X"6f", X"76", 
  X"20", X"31", X"35", X"20", X"32", X"30", X"31", X"32", 
  X"0a", X"0a", X"00", X"00", X"43", X"4f", X"44", X"45", 
  X"2e", X"42", X"49", X"4e", X"00", X"00", X"00", X"00", 
  X"4c", X"6f", X"61", X"64", X"69", X"6e", X"67", X"20", 
  X"66", X"69", X"6c", X"65", X"20", X"27", X"2f", X"63", 
  X"6f", X"64", X"65", X"2e", X"62", X"69", X"6e", X"27", 
  X"20", X"6f", X"6e", X"74", X"6f", X"20", X"52", X"41", 
  X"4d", X"20", X"61", X"74", X"20", X"61", X"64", X"64", 
  X"72", X"65", X"73", X"73", X"20", X"30", X"78", X"30", 
  X"30", X"30", X"30", X"30", X"30", X"30", X"30", X"2e", 
  X"2e", X"2e", X"0a", X"00", X"44", X"6f", X"6e", X"65", 
  X"2e", X"20", X"52", X"65", X"61", X"64", X"20", X"25", 
  X"75", X"20", X"62", X"79", X"74", X"65", X"73", X"2e", 
  X"0a", X"00", X"00", X"00", X"54", X"72", X"61", X"6e", 
  X"73", X"66", X"65", X"72", X"72", X"69", X"6e", X"67", 
  X"20", X"63", X"6f", X"6e", X"74", X"72", X"6f", X"6c", 
  X"20", X"74", X"6f", X"20", X"61", X"64", X"64", X"72", 
  X"65", X"73", X"73", X"20", X"30", X"78", X"30", X"30", 
  X"30", X"30", X"30", X"30", X"30", X"30", X"0a", X"0a", 
  X"00", X"00", X"00", X"00", X"22", X"2a", X"2b", X"2c", 
  X"3a", X"3b", X"3c", X"3d", X"3e", X"3f", X"5b", X"5d", 
  X"7c", X"7f", X"00", X"00", X"28", X"6e", X"75", X"6c", 
  X"6c", X"29", X"00", X"00", X"01" );



end package obj_code_pkg;
