-- Rom file for twiddle factors 
-- ../../../rtl/vhdl/WISHBONE_FFT/rom1.vhd contains 1024 points of 16 width 
--  for a 1024 point fft.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;


ENTITY rom1 IS
         GENERIC(
        data_width : integer :=16;
        address_width : integer :=10
    );
    PORT(
        clk :in std_logic;
        address :in std_logic_vector (9      downto 0);
        datar : OUT std_logic_vector (data_width-1 DOWNTO 0) ;
        datai : OUT std_logic_vector (data_width-1 DOWNTO 0)
    );
end rom1;
ARCHITECTURE behavior OF rom1 IS

 BEGIN

process (address,clk)
begin
    	if(rising_edge(clk)) then 
 case address is
        when "0000000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "0000000001" => datar <= "0111111111111101";datai <= "1111111001101110"; --2
        when "0000000010" => datar <= "0111111111110101";datai <= "1111110011011100"; --4
        when "0000000011" => datar <= "0111111111101001";datai <= "1111101101001010"; --6
        when "0000000100" => datar <= "0111111111011000";datai <= "1111100110111000"; --8
        when "0000000101" => datar <= "0111111111000001";datai <= "1111100000100111"; --10
        when "0000000110" => datar <= "0111111110100110";datai <= "1111011010010110"; --12
        when "0000000111" => datar <= "0111111110000110";datai <= "1111010100000101"; --14
        when "0000001000" => datar <= "0111111101100001";datai <= "1111001101110100"; --16
        when "0000001001" => datar <= "0111111100110111";datai <= "1111000111100100"; --18
        when "0000001010" => datar <= "0111111100001001";datai <= "1111000001010101"; --20
        when "0000001011" => datar <= "0111111011010101";datai <= "1110111011000110"; --22
        when "0000001100" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "0000001101" => datar <= "0111111001011111";datai <= "1110101110101011"; --26
        when "0000001110" => datar <= "0111111000011101";datai <= "1110101000011110"; --28
        when "0000001111" => datar <= "0111110111010101";datai <= "1110100010010010"; --30
        when "0000010000" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "0000010001" => datar <= "0111110100111001";datai <= "1110010101111110"; --34
        when "0000010010" => datar <= "0111110011100011";datai <= "1110001111110101"; --36
        when "0000010011" => datar <= "0111110010001000";datai <= "1110001001101101"; --38
        when "0000010100" => datar <= "0111110000101001";datai <= "1110000011100110"; --40
        when "0000010101" => datar <= "0111101111000101";datai <= "1101111101100001"; --42
        when "0000010110" => datar <= "0111101101011100";datai <= "1101110111011101"; --44
        when "0000010111" => datar <= "0111101011101110";datai <= "1101110001011010"; --46
        when "0000011000" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "0000011001" => datar <= "0111101000000101";datai <= "1101100101011000"; --50
        when "0000011010" => datar <= "0111100110001001";datai <= "1101011111011010"; --52
        when "0000011011" => datar <= "0111100100001001";datai <= "1101011001011101"; --54
        when "0000011100" => datar <= "0111100010000100";datai <= "1101010011100001"; --56
        when "0000011101" => datar <= "0111011111111010";datai <= "1101001101100111"; --58
        when "0000011110" => datar <= "0111011101101011";datai <= "1101000111101111"; --60
        when "0000011111" => datar <= "0111011011011000";datai <= "1101000001111001"; --62
        when "0000100000" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "0000100001" => datar <= "0111010110100101";datai <= "1100110110010010"; --66
        when "0000100010" => datar <= "0111010100000100";datai <= "1100110000100001"; --68
        when "0000100011" => datar <= "0111010001011111";datai <= "1100101010110011"; --70
        when "0000100100" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "0000100101" => datar <= "0111001100000111";datai <= "1100011111011100"; --74
        when "0000100110" => datar <= "0111001001010100";datai <= "1100011001110100"; --76
        when "0000100111" => datar <= "0111000110011101";datai <= "1100010100001110"; --78
        when "0000101000" => datar <= "0111000011100010";datai <= "1100001110101010"; --80
        when "0000101001" => datar <= "0111000000100010";datai <= "1100001001001000"; --82
        when "0000101010" => datar <= "0110111101011110";datai <= "1100000011101001"; --84
        when "0000101011" => datar <= "0110111010010110";datai <= "1011111110001101"; --86
        when "0000101100" => datar <= "0110110111001001";datai <= "1011111000110010"; --88
        when "0000101101" => datar <= "0110110011111000";datai <= "1011110011011011"; --90
        when "0000101110" => datar <= "0110110000100011";datai <= "1011101110000110"; --92
        when "0000101111" => datar <= "0110101101001010";datai <= "1011101000110011"; --94
        when "0000110000" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "0000110001" => datar <= "0110100110001011";datai <= "1011011110010111"; --98
        when "0000110010" => datar <= "0110100010100110";datai <= "1011011001001100"; --100
        when "0000110011" => datar <= "0110011110111100";datai <= "1011010100000101"; --102
        when "0000110100" => datar <= "0110011011001111";datai <= "1011001111000001"; --104
        when "0000110101" => datar <= "0110010111011101";datai <= "1011001001111111"; --106
        when "0000110110" => datar <= "0110010011101000";datai <= "1011000101000001"; --108
        when "0000110111" => datar <= "0110001111101110";datai <= "1011000000000101"; --110
        when "0000111000" => datar <= "0110001011110001";datai <= "1010111011001101"; --112
        when "0000111001" => datar <= "0110000111110000";datai <= "1010110110011000"; --114
        when "0000111010" => datar <= "0110000011101011";datai <= "1010110001100101"; --116
        when "0000111011" => datar <= "0101111111100011";datai <= "1010101100110111"; --118
        when "0000111100" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "0000111101" => datar <= "0101110111000111";datai <= "1010100011100011"; --122
        when "0000111110" => datar <= "0101110010110011";datai <= "1010011110111110"; --124
        when "0000111111" => datar <= "0101101110011100";datai <= "1010011010011100"; --126
        when "0001000000" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "0001000001" => datar <= "0101100101100100";datai <= "1010010001100100"; --130
        when "0001000010" => datar <= "0101100001000010";datai <= "1010001101001101"; --132
        when "0001000011" => datar <= "0101011100011101";datai <= "1010001000111001"; --134
        when "0001000100" => datar <= "0101010111110101";datai <= "1010000100101001"; --136
        when "0001000101" => datar <= "0101010011001001";datai <= "1010000000011101"; --138
        when "0001000110" => datar <= "0101001110011011";datai <= "1001111100010101"; --140
        when "0001000111" => datar <= "0101001001101000";datai <= "1001111000010000"; --142
        when "0001001000" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "0001001001" => datar <= "0100111111111011";datai <= "1001110000010010"; --146
        when "0001001010" => datar <= "0100111010111111";datai <= "1001101100011000"; --148
        when "0001001011" => datar <= "0100110110000001";datai <= "1001101000100011"; --150
        when "0001001100" => datar <= "0100110000111111";datai <= "1001100100110001"; --152
        when "0001001101" => datar <= "0100101011111011";datai <= "1001100001000100"; --154
        when "0001001110" => datar <= "0100100110110100";datai <= "1001011101011010"; --156
        when "0001001111" => datar <= "0100100001101001";datai <= "1001011001110101"; --158
        when "0001010000" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "0001010001" => datar <= "0100010111001101";datai <= "1001010010110110"; --162
        when "0001010010" => datar <= "0100010001111010";datai <= "1001001111011101"; --164
        when "0001010011" => datar <= "0100001100100101";datai <= "1001001100001000"; --166
        when "0001010100" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "0001010101" => datar <= "0100000001110011";datai <= "1001000101101010"; --170
        when "0001010110" => datar <= "0011111100010111";datai <= "1001000010100010"; --172
        when "0001010111" => datar <= "0011110110111000";datai <= "1000111111011110"; --174
        when "0001011000" => datar <= "0011110001010110";datai <= "1000111100011110"; --176
        when "0001011001" => datar <= "0011101011110010";datai <= "1000111001100011"; --178
        when "0001011010" => datar <= "0011100110001100";datai <= "1000110110101100"; --180
        when "0001011011" => datar <= "0011100000100100";datai <= "1000110011111001"; --182
        when "0001011100" => datar <= "0011011010111010";datai <= "1000110001001011"; --184
        when "0001011101" => datar <= "0011010101001101";datai <= "1000101110100001"; --186
        when "0001011110" => datar <= "0011001111011111";datai <= "1000101011111100"; --188
        when "0001011111" => datar <= "0011001001101110";datai <= "1000101001011011"; --190
        when "0001100000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "0001100001" => datar <= "0010111110000111";datai <= "1000100100101000"; --194
        when "0001100010" => datar <= "0010111000010001";datai <= "1000100010010101"; --196
        when "0001100011" => datar <= "0010110010011001";datai <= "1000100000000110"; --198
        when "0001100100" => datar <= "0010101100011111";datai <= "1000011101111100"; --200
        when "0001100101" => datar <= "0010100110100011";datai <= "1000011011110111"; --202
        when "0001100110" => datar <= "0010100000100110";datai <= "1000011001110111"; --204
        when "0001100111" => datar <= "0010011010101000";datai <= "1000010111111011"; --206
        when "0001101000" => datar <= "0010010100101000";datai <= "1000010110000100"; --208
        when "0001101001" => datar <= "0010001110100110";datai <= "1000010100010010"; --210
        when "0001101010" => datar <= "0010001000100011";datai <= "1000010010100100"; --212
        when "0001101011" => datar <= "0010000010011111";datai <= "1000010000111011"; --214
        when "0001101100" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "0001101101" => datar <= "0001110110010011";datai <= "1000001101111000"; --218
        when "0001101110" => datar <= "0001110000001011";datai <= "1000001100011101"; --220
        when "0001101111" => datar <= "0001101010000010";datai <= "1000001011000111"; --222
        when "0001110000" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "0001110001" => datar <= "0001011101101110";datai <= "1000001000101011"; --226
        when "0001110010" => datar <= "0001010111100010";datai <= "1000000111100011"; --228
        when "0001110011" => datar <= "0001010001010101";datai <= "1000000110100001"; --230
        when "0001110100" => datar <= "0001001011001000";datai <= "1000000101100100"; --232
        when "0001110101" => datar <= "0001000100111010";datai <= "1000000100101011"; --234
        when "0001110110" => datar <= "0000111110101011";datai <= "1000000011110111"; --236
        when "0001110111" => datar <= "0000111000011100";datai <= "1000000011001001"; --238
        when "0001111000" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "0001111001" => datar <= "0000101011111011";datai <= "1000000001111010"; --242
        when "0001111010" => datar <= "0000100101101010";datai <= "1000000001011010"; --244
        when "0001111011" => datar <= "0000011111011001";datai <= "1000000000111111"; --246
        when "0001111100" => datar <= "0000011001001000";datai <= "1000000000101000"; --248
        when "0001111101" => datar <= "0000010010110110";datai <= "1000000000010111"; --250
        when "0001111110" => datar <= "0000001100100100";datai <= "1000000000001011"; --252
        when "0001111111" => datar <= "0000000110010010";datai <= "1000000000000011"; --254
        when "0010000000" => datar <= "0000000000000000";datai <= "1000000000000001"; --256
        when "0010000001" => datar <= "1111111001101110";datai <= "1000000000000011"; --258
        when "0010000010" => datar <= "1111110011011100";datai <= "1000000000001011"; --260
        when "0010000011" => datar <= "1111101101001010";datai <= "1000000000010111"; --262
        when "0010000100" => datar <= "1111100110111000";datai <= "1000000000101000"; --264
        when "0010000101" => datar <= "1111100000100111";datai <= "1000000000111111"; --266
        when "0010000110" => datar <= "1111011010010110";datai <= "1000000001011010"; --268
        when "0010000111" => datar <= "1111010100000101";datai <= "1000000001111010"; --270
        when "0010001000" => datar <= "1111001101110100";datai <= "1000000010011111"; --272
        when "0010001001" => datar <= "1111000111100100";datai <= "1000000011001001"; --274
        when "0010001010" => datar <= "1111000001010101";datai <= "1000000011110111"; --276
        when "0010001011" => datar <= "1110111011000110";datai <= "1000000100101011"; --278
        when "0010001100" => datar <= "1110110100111000";datai <= "1000000101100100"; --280
        when "0010001101" => datar <= "1110101110101011";datai <= "1000000110100001"; --282
        when "0010001110" => datar <= "1110101000011110";datai <= "1000000111100011"; --284
        when "0010001111" => datar <= "1110100010010010";datai <= "1000001000101011"; --286
        when "0010010000" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "0010010001" => datar <= "1110010101111110";datai <= "1000001011000111"; --290
        when "0010010010" => datar <= "1110001111110101";datai <= "1000001100011101"; --292
        when "0010010011" => datar <= "1110001001101101";datai <= "1000001101111000"; --294
        when "0010010100" => datar <= "1110000011100110";datai <= "1000001111010111"; --296
        when "0010010101" => datar <= "1101111101100001";datai <= "1000010000111011"; --298
        when "0010010110" => datar <= "1101110111011101";datai <= "1000010010100100"; --300
        when "0010010111" => datar <= "1101110001011010";datai <= "1000010100010010"; --302
        when "0010011000" => datar <= "1101101011011000";datai <= "1000010110000100"; --304
        when "0010011001" => datar <= "1101100101011000";datai <= "1000010111111011"; --306
        when "0010011010" => datar <= "1101011111011010";datai <= "1000011001110111"; --308
        when "0010011011" => datar <= "1101011001011101";datai <= "1000011011110111"; --310
        when "0010011100" => datar <= "1101010011100001";datai <= "1000011101111100"; --312
        when "0010011101" => datar <= "1101001101100111";datai <= "1000100000000110"; --314
        when "0010011110" => datar <= "1101000111101111";datai <= "1000100010010101"; --316
        when "0010011111" => datar <= "1101000001111001";datai <= "1000100100101000"; --318
        when "0010100000" => datar <= "1100111100000101";datai <= "1000100110111111"; --320
        when "0010100001" => datar <= "1100110110010010";datai <= "1000101001011011"; --322
        when "0010100010" => datar <= "1100110000100001";datai <= "1000101011111100"; --324
        when "0010100011" => datar <= "1100101010110011";datai <= "1000101110100001"; --326
        when "0010100100" => datar <= "1100100101000110";datai <= "1000110001001011"; --328
        when "0010100101" => datar <= "1100011111011100";datai <= "1000110011111001"; --330
        when "0010100110" => datar <= "1100011001110100";datai <= "1000110110101100"; --332
        when "0010100111" => datar <= "1100010100001110";datai <= "1000111001100011"; --334
        when "0010101000" => datar <= "1100001110101010";datai <= "1000111100011110"; --336
        when "0010101001" => datar <= "1100001001001000";datai <= "1000111111011110"; --338
        when "0010101010" => datar <= "1100000011101001";datai <= "1001000010100010"; --340
        when "0010101011" => datar <= "1011111110001101";datai <= "1001000101101010"; --342
        when "0010101100" => datar <= "1011111000110010";datai <= "1001001000110111"; --344
        when "0010101101" => datar <= "1011110011011011";datai <= "1001001100001000"; --346
        when "0010101110" => datar <= "1011101110000110";datai <= "1001001111011101"; --348
        when "0010101111" => datar <= "1011101000110011";datai <= "1001010010110110"; --350
        when "0010110000" => datar <= "1011100011100100";datai <= "1001010110010011"; --352
        when "0010110001" => datar <= "1011011110010111";datai <= "1001011001110101"; --354
        when "0010110010" => datar <= "1011011001001100";datai <= "1001011101011010"; --356
        when "0010110011" => datar <= "1011010100000101";datai <= "1001100001000100"; --358
        when "0010110100" => datar <= "1011001111000001";datai <= "1001100100110001"; --360
        when "0010110101" => datar <= "1011001001111111";datai <= "1001101000100011"; --362
        when "0010110110" => datar <= "1011000101000001";datai <= "1001101100011000"; --364
        when "0010110111" => datar <= "1011000000000101";datai <= "1001110000010010"; --366
        when "0010111000" => datar <= "1010111011001101";datai <= "1001110100001111"; --368
        when "0010111001" => datar <= "1010110110011000";datai <= "1001111000010000"; --370
        when "0010111010" => datar <= "1010110001100101";datai <= "1001111100010101"; --372
        when "0010111011" => datar <= "1010101100110111";datai <= "1010000000011101"; --374
        when "0010111100" => datar <= "1010101000001011";datai <= "1010000100101001"; --376
        when "0010111101" => datar <= "1010100011100011";datai <= "1010001000111001"; --378
        when "0010111110" => datar <= "1010011110111110";datai <= "1010001101001101"; --380
        when "0010111111" => datar <= "1010011010011100";datai <= "1010010001100100"; --382
        when "0011000000" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "0011000001" => datar <= "1010010001100100";datai <= "1010011010011100"; --386
        when "0011000010" => datar <= "1010001101001101";datai <= "1010011110111110"; --388
        when "0011000011" => datar <= "1010001000111001";datai <= "1010100011100011"; --390
        when "0011000100" => datar <= "1010000100101001";datai <= "1010101000001011"; --392
        when "0011000101" => datar <= "1010000000011101";datai <= "1010101100110111"; --394
        when "0011000110" => datar <= "1001111100010101";datai <= "1010110001100101"; --396
        when "0011000111" => datar <= "1001111000010000";datai <= "1010110110011000"; --398
        when "0011001000" => datar <= "1001110100001111";datai <= "1010111011001101"; --400
        when "0011001001" => datar <= "1001110000010010";datai <= "1011000000000101"; --402
        when "0011001010" => datar <= "1001101100011000";datai <= "1011000101000001"; --404
        when "0011001011" => datar <= "1001101000100011";datai <= "1011001001111111"; --406
        when "0011001100" => datar <= "1001100100110001";datai <= "1011001111000001"; --408
        when "0011001101" => datar <= "1001100001000100";datai <= "1011010100000101"; --410
        when "0011001110" => datar <= "1001011101011010";datai <= "1011011001001100"; --412
        when "0011001111" => datar <= "1001011001110101";datai <= "1011011110010111"; --414
        when "0011010000" => datar <= "1001010110010011";datai <= "1011100011100100"; --416
        when "0011010001" => datar <= "1001010010110110";datai <= "1011101000110011"; --418
        when "0011010010" => datar <= "1001001111011101";datai <= "1011101110000110"; --420
        when "0011010011" => datar <= "1001001100001000";datai <= "1011110011011011"; --422
        when "0011010100" => datar <= "1001001000110111";datai <= "1011111000110010"; --424
        when "0011010101" => datar <= "1001000101101010";datai <= "1011111110001101"; --426
        when "0011010110" => datar <= "1001000010100010";datai <= "1100000011101001"; --428
        when "0011010111" => datar <= "1000111111011110";datai <= "1100001001001000"; --430
        when "0011011000" => datar <= "1000111100011110";datai <= "1100001110101010"; --432
        when "0011011001" => datar <= "1000111001100011";datai <= "1100010100001110"; --434
        when "0011011010" => datar <= "1000110110101100";datai <= "1100011001110100"; --436
        when "0011011011" => datar <= "1000110011111001";datai <= "1100011111011100"; --438
        when "0011011100" => datar <= "1000110001001011";datai <= "1100100101000110"; --440
        when "0011011101" => datar <= "1000101110100001";datai <= "1100101010110011"; --442
        when "0011011110" => datar <= "1000101011111100";datai <= "1100110000100001"; --444
        when "0011011111" => datar <= "1000101001011011";datai <= "1100110110010010"; --446
        when "0011100000" => datar <= "1000100110111111";datai <= "1100111100000101"; --448
        when "0011100001" => datar <= "1000100100101000";datai <= "1101000001111001"; --450
        when "0011100010" => datar <= "1000100010010101";datai <= "1101000111101111"; --452
        when "0011100011" => datar <= "1000100000000110";datai <= "1101001101100111"; --454
        when "0011100100" => datar <= "1000011101111100";datai <= "1101010011100001"; --456
        when "0011100101" => datar <= "1000011011110111";datai <= "1101011001011101"; --458
        when "0011100110" => datar <= "1000011001110111";datai <= "1101011111011010"; --460
        when "0011100111" => datar <= "1000010111111011";datai <= "1101100101011000"; --462
        when "0011101000" => datar <= "1000010110000100";datai <= "1101101011011000"; --464
        when "0011101001" => datar <= "1000010100010010";datai <= "1101110001011010"; --466
        when "0011101010" => datar <= "1000010010100100";datai <= "1101110111011101"; --468
        when "0011101011" => datar <= "1000010000111011";datai <= "1101111101100001"; --470
        when "0011101100" => datar <= "1000001111010111";datai <= "1110000011100110"; --472
        when "0011101101" => datar <= "1000001101111000";datai <= "1110001001101101"; --474
        when "0011101110" => datar <= "1000001100011101";datai <= "1110001111110101"; --476
        when "0011101111" => datar <= "1000001011000111";datai <= "1110010101111110"; --478
        when "0011110000" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "0011110001" => datar <= "1000001000101011";datai <= "1110100010010010"; --482
        when "0011110010" => datar <= "1000000111100011";datai <= "1110101000011110"; --484
        when "0011110011" => datar <= "1000000110100001";datai <= "1110101110101011"; --486
        when "0011110100" => datar <= "1000000101100100";datai <= "1110110100111000"; --488
        when "0011110101" => datar <= "1000000100101011";datai <= "1110111011000110"; --490
        when "0011110110" => datar <= "1000000011110111";datai <= "1111000001010101"; --492
        when "0011110111" => datar <= "1000000011001001";datai <= "1111000111100100"; --494
        when "0011111000" => datar <= "1000000010011111";datai <= "1111001101110100"; --496
        when "0011111001" => datar <= "1000000001111010";datai <= "1111010100000101"; --498
        when "0011111010" => datar <= "1000000001011010";datai <= "1111011010010110"; --500
        when "0011111011" => datar <= "1000000000111111";datai <= "1111100000100111"; --502
        when "0011111100" => datar <= "1000000000101000";datai <= "1111100110111000"; --504
        when "0011111101" => datar <= "1000000000010111";datai <= "1111101101001010"; --506
        when "0011111110" => datar <= "1000000000001011";datai <= "1111110011011100"; --508
        when "0011111111" => datar <= "1000000000000011";datai <= "1111111001101110"; --510
        when "0100000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "0100000001" => datar <= "0111111111111110";datai <= "1111111100110111"; --1
        when "0100000010" => datar <= "0111111111111101";datai <= "1111111001101110"; --2
        when "0100000011" => datar <= "0111111111111001";datai <= "1111110110100101"; --3
        when "0100000100" => datar <= "0111111111110101";datai <= "1111110011011100"; --4
        when "0100000101" => datar <= "0111111111110000";datai <= "1111110000010011"; --5
        when "0100000110" => datar <= "0111111111101001";datai <= "1111101101001010"; --6
        when "0100000111" => datar <= "0111111111100001";datai <= "1111101010000001"; --7
        when "0100001000" => datar <= "0111111111011000";datai <= "1111100110111000"; --8
        when "0100001001" => datar <= "0111111111001101";datai <= "1111100011101111"; --9
        when "0100001010" => datar <= "0111111111000001";datai <= "1111100000100111"; --10
        when "0100001011" => datar <= "0111111110110100";datai <= "1111011101011110"; --11
        when "0100001100" => datar <= "0111111110100110";datai <= "1111011010010110"; --12
        when "0100001101" => datar <= "0111111110010111";datai <= "1111010111001101"; --13
        when "0100001110" => datar <= "0111111110000110";datai <= "1111010100000101"; --14
        when "0100001111" => datar <= "0111111101110100";datai <= "1111010000111100"; --15
        when "0100010000" => datar <= "0111111101100001";datai <= "1111001101110100"; --16
        when "0100010001" => datar <= "0111111101001101";datai <= "1111001010101100"; --17
        when "0100010010" => datar <= "0111111100110111";datai <= "1111000111100100"; --18
        when "0100010011" => datar <= "0111111100100001";datai <= "1111000100011101"; --19
        when "0100010100" => datar <= "0111111100001001";datai <= "1111000001010101"; --20
        when "0100010101" => datar <= "0111111011101111";datai <= "1110111110001110"; --21
        when "0100010110" => datar <= "0111111011010101";datai <= "1110111011000110"; --22
        when "0100010111" => datar <= "0111111010111001";datai <= "1110110111111111"; --23
        when "0100011000" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "0100011001" => datar <= "0111111001111110";datai <= "1110110001110001"; --25
        when "0100011010" => datar <= "0111111001011111";datai <= "1110101110101011"; --26
        when "0100011011" => datar <= "0111111000111110";datai <= "1110101011100100"; --27
        when "0100011100" => datar <= "0111111000011101";datai <= "1110101000011110"; --28
        when "0100011101" => datar <= "0111110111111010";datai <= "1110100101011000"; --29
        when "0100011110" => datar <= "0111110111010101";datai <= "1110100010010010"; --30
        when "0100011111" => datar <= "0111110110110000";datai <= "1110011111001101"; --31
        when "0100100000" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "0100100001" => datar <= "0111110101100010";datai <= "1110011001000010"; --33
        when "0100100010" => datar <= "0111110100111001";datai <= "1110010101111110"; --34
        when "0100100011" => datar <= "0111110100001110";datai <= "1110010010111001"; --35
        when "0100100100" => datar <= "0111110011100011";datai <= "1110001111110101"; --36
        when "0100100101" => datar <= "0111110010110110";datai <= "1110001100110001"; --37
        when "0100100110" => datar <= "0111110010001000";datai <= "1110001001101101"; --38
        when "0100100111" => datar <= "0111110001011001";datai <= "1110000110101001"; --39
        when "0100101000" => datar <= "0111110000101001";datai <= "1110000011100110"; --40
        when "0100101001" => datar <= "0111101111111000";datai <= "1110000000100011"; --41
        when "0100101010" => datar <= "0111101111000101";datai <= "1101111101100001"; --42
        when "0100101011" => datar <= "0111101110010001";datai <= "1101111010011111"; --43
        when "0100101100" => datar <= "0111101101011100";datai <= "1101110111011101"; --44
        when "0100101101" => datar <= "0111101100100110";datai <= "1101110100011011"; --45
        when "0100101110" => datar <= "0111101011101110";datai <= "1101110001011010"; --46
        when "0100101111" => datar <= "0111101010110110";datai <= "1101101110011001"; --47
        when "0100110000" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "0100110001" => datar <= "0111101001000001";datai <= "1101101000011000"; --49
        when "0100110010" => datar <= "0111101000000101";datai <= "1101100101011000"; --50
        when "0100110011" => datar <= "0111100111001000";datai <= "1101100010011001"; --51
        when "0100110100" => datar <= "0111100110001001";datai <= "1101011111011010"; --52
        when "0100110101" => datar <= "0111100101001010";datai <= "1101011100011011"; --53
        when "0100110110" => datar <= "0111100100001001";datai <= "1101011001011101"; --54
        when "0100110111" => datar <= "0111100011000111";datai <= "1101010110011111"; --55
        when "0100111000" => datar <= "0111100010000100";datai <= "1101010011100001"; --56
        when "0100111001" => datar <= "0111100000111111";datai <= "1101010000100100"; --57
        when "0100111010" => datar <= "0111011111111010";datai <= "1101001101100111"; --58
        when "0100111011" => datar <= "0111011110110011";datai <= "1101001010101011"; --59
        when "0100111100" => datar <= "0111011101101011";datai <= "1101000111101111"; --60
        when "0100111101" => datar <= "0111011100100010";datai <= "1101000100110100"; --61
        when "0100111110" => datar <= "0111011011011000";datai <= "1101000001111001"; --62
        when "0100111111" => datar <= "0111011010001101";datai <= "1100111110111111"; --63
        when "0101000000" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "0101000001" => datar <= "0111010111110011";datai <= "1100111001001011"; --65
        when "0101000010" => datar <= "0111010110100101";datai <= "1100110110010010"; --66
        when "0101000011" => datar <= "0111010101010101";datai <= "1100110011011010"; --67
        when "0101000100" => datar <= "0111010100000100";datai <= "1100110000100001"; --68
        when "0101000101" => datar <= "0111010010110010";datai <= "1100101101101010"; --69
        when "0101000110" => datar <= "0111010001011111";datai <= "1100101010110011"; --70
        when "0101000111" => datar <= "0111010000001010";datai <= "1100100111111100"; --71
        when "0101001000" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "0101001001" => datar <= "0111001101011110";datai <= "1100100010010001"; --73
        when "0101001010" => datar <= "0111001100000111";datai <= "1100011111011100"; --74
        when "0101001011" => datar <= "0111001010101110";datai <= "1100011100100111"; --75
        when "0101001100" => datar <= "0111001001010100";datai <= "1100011001110100"; --76
        when "0101001101" => datar <= "0111000111111001";datai <= "1100010111000000"; --77
        when "0101001110" => datar <= "0111000110011101";datai <= "1100010100001110"; --78
        when "0101001111" => datar <= "0111000101000000";datai <= "1100010001011011"; --79
        when "0101010000" => datar <= "0111000011100010";datai <= "1100001110101010"; --80
        when "0101010001" => datar <= "0111000010000011";datai <= "1100001011111001"; --81
        when "0101010010" => datar <= "0111000000100010";datai <= "1100001001001000"; --82
        when "0101010011" => datar <= "0110111111000001";datai <= "1100000110011000"; --83
        when "0101010100" => datar <= "0110111101011110";datai <= "1100000011101001"; --84
        when "0101010101" => datar <= "0110111011111011";datai <= "1100000000111011"; --85
        when "0101010110" => datar <= "0110111010010110";datai <= "1011111110001101"; --86
        when "0101010111" => datar <= "0110111000110000";datai <= "1011111011011111"; --87
        when "0101011000" => datar <= "0110110111001001";datai <= "1011111000110010"; --88
        when "0101011001" => datar <= "0110110101100001";datai <= "1011110110000110"; --89
        when "0101011010" => datar <= "0110110011111000";datai <= "1011110011011011"; --90
        when "0101011011" => datar <= "0110110010001110";datai <= "1011110000110000"; --91
        when "0101011100" => datar <= "0110110000100011";datai <= "1011101110000110"; --92
        when "0101011101" => datar <= "0110101110110111";datai <= "1011101011011100"; --93
        when "0101011110" => datar <= "0110101101001010";datai <= "1011101000110011"; --94
        when "0101011111" => datar <= "0110101011011100";datai <= "1011100110001011"; --95
        when "0101100000" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "0101100001" => datar <= "0110100111111101";datai <= "1011100000111101"; --97
        when "0101100010" => datar <= "0110100110001011";datai <= "1011011110010111"; --98
        when "0101100011" => datar <= "0110100100011001";datai <= "1011011011110001"; --99
        when "0101100100" => datar <= "0110100010100110";datai <= "1011011001001100"; --100
        when "0101100101" => datar <= "0110100000110010";datai <= "1011010110101000"; --101
        when "0101100110" => datar <= "0110011110111100";datai <= "1011010100000101"; --102
        when "0101100111" => datar <= "0110011101000110";datai <= "1011010001100011"; --103
        when "0101101000" => datar <= "0110011011001111";datai <= "1011001111000001"; --104
        when "0101101001" => datar <= "0110011001010110";datai <= "1011001100100000"; --105
        when "0101101010" => datar <= "0110010111011101";datai <= "1011001001111111"; --106
        when "0101101011" => datar <= "0110010101100011";datai <= "1011000111100000"; --107
        when "0101101100" => datar <= "0110010011101000";datai <= "1011000101000001"; --108
        when "0101101101" => datar <= "0110010001101100";datai <= "1011000010100011"; --109
        when "0101101110" => datar <= "0110001111101110";datai <= "1011000000000101"; --110
        when "0101101111" => datar <= "0110001101110000";datai <= "1010111101101001"; --111
        when "0101110000" => datar <= "0110001011110001";datai <= "1010111011001101"; --112
        when "0101110001" => datar <= "0110001001110001";datai <= "1010111000110010"; --113
        when "0101110010" => datar <= "0110000111110000";datai <= "1010110110011000"; --114
        when "0101110011" => datar <= "0110000101101110";datai <= "1010110011111110"; --115
        when "0101110100" => datar <= "0110000011101011";datai <= "1010110001100101"; --116
        when "0101110101" => datar <= "0110000001101000";datai <= "1010101111001110"; --117
        when "0101110110" => datar <= "0101111111100011";datai <= "1010101100110111"; --118
        when "0101110111" => datar <= "0101111101011101";datai <= "1010101010100000"; --119
        when "0101111000" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "0101111001" => datar <= "0101111001001111";datai <= "1010100101110110"; --121
        when "0101111010" => datar <= "0101110111000111";datai <= "1010100011100011"; --122
        when "0101111011" => datar <= "0101110100111110";datai <= "1010100001010000"; --123
        when "0101111100" => datar <= "0101110010110011";datai <= "1010011110111110"; --124
        when "0101111101" => datar <= "0101110000101000";datai <= "1010011100101101"; --125
        when "0101111110" => datar <= "0101101110011100";datai <= "1010011010011100"; --126
        when "0101111111" => datar <= "0101101100001111";datai <= "1010011000001101"; --127
        when "0110000000" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "0110000001" => datar <= "0101100111110011";datai <= "1010010011110001"; --129
        when "0110000010" => datar <= "0101100101100100";datai <= "1010010001100100"; --130
        when "0110000011" => datar <= "0101100011010011";datai <= "1010001111011000"; --131
        when "0110000100" => datar <= "0101100001000010";datai <= "1010001101001101"; --132
        when "0110000101" => datar <= "0101011110110000";datai <= "1010001011000010"; --133
        when "0110000110" => datar <= "0101011100011101";datai <= "1010001000111001"; --134
        when "0110000111" => datar <= "0101011010001010";datai <= "1010000110110001"; --135
        when "0110001000" => datar <= "0101010111110101";datai <= "1010000100101001"; --136
        when "0110001001" => datar <= "0101010101100000";datai <= "1010000010100011"; --137
        when "0110001010" => datar <= "0101010011001001";datai <= "1010000000011101"; --138
        when "0110001011" => datar <= "0101010000110010";datai <= "1001111110011000"; --139
        when "0110001100" => datar <= "0101001110011011";datai <= "1001111100010101"; --140
        when "0110001101" => datar <= "0101001100000010";datai <= "1001111010010010"; --141
        when "0110001110" => datar <= "0101001001101000";datai <= "1001111000010000"; --142
        when "0110001111" => datar <= "0101000111001110";datai <= "1001110110001111"; --143
        when "0110010000" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "0110010001" => datar <= "0101000010010111";datai <= "1001110010010000"; --145
        when "0110010010" => datar <= "0100111111111011";datai <= "1001110000010010"; --146
        when "0110010011" => datar <= "0100111101011101";datai <= "1001101110010100"; --147
        when "0110010100" => datar <= "0100111010111111";datai <= "1001101100011000"; --148
        when "0110010101" => datar <= "0100111000100000";datai <= "1001101010011101"; --149
        when "0110010110" => datar <= "0100110110000001";datai <= "1001101000100011"; --150
        when "0110010111" => datar <= "0100110011100000";datai <= "1001100110101010"; --151
        when "0110011000" => datar <= "0100110000111111";datai <= "1001100100110001"; --152
        when "0110011001" => datar <= "0100101110011101";datai <= "1001100010111010"; --153
        when "0110011010" => datar <= "0100101011111011";datai <= "1001100001000100"; --154
        when "0110011011" => datar <= "0100101001011000";datai <= "1001011111001110"; --155
        when "0110011100" => datar <= "0100100110110100";datai <= "1001011101011010"; --156
        when "0110011101" => datar <= "0100100100001111";datai <= "1001011011100111"; --157
        when "0110011110" => datar <= "0100100001101001";datai <= "1001011001110101"; --158
        when "0110011111" => datar <= "0100011111000011";datai <= "1001011000000011"; --159
        when "0110100000" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "0110100001" => datar <= "0100011001110101";datai <= "1001010100100100"; --161
        when "0110100010" => datar <= "0100010111001101";datai <= "1001010010110110"; --162
        when "0110100011" => datar <= "0100010100100100";datai <= "1001010001001001"; --163
        when "0110100100" => datar <= "0100010001111010";datai <= "1001001111011101"; --164
        when "0110100101" => datar <= "0100001111010000";datai <= "1001001101110010"; --165
        when "0110100110" => datar <= "0100001100100101";datai <= "1001001100001000"; --166
        when "0110100111" => datar <= "0100001001111010";datai <= "1001001010011111"; --167
        when "0110101000" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "0110101001" => datar <= "0100000100100001";datai <= "1001000111010000"; --169
        when "0110101010" => datar <= "0100000001110011";datai <= "1001000101101010"; --170
        when "0110101011" => datar <= "0011111111000101";datai <= "1001000100000101"; --171
        when "0110101100" => datar <= "0011111100010111";datai <= "1001000010100010"; --172
        when "0110101101" => datar <= "0011111001101000";datai <= "1001000000111111"; --173
        when "0110101110" => datar <= "0011110110111000";datai <= "1000111111011110"; --174
        when "0110101111" => datar <= "0011110100000111";datai <= "1000111101111101"; --175
        when "0110110000" => datar <= "0011110001010110";datai <= "1000111100011110"; --176
        when "0110110001" => datar <= "0011101110100101";datai <= "1000111011000000"; --177
        when "0110110010" => datar <= "0011101011110010";datai <= "1000111001100011"; --178
        when "0110110011" => datar <= "0011101001000000";datai <= "1000111000000111"; --179
        when "0110110100" => datar <= "0011100110001100";datai <= "1000110110101100"; --180
        when "0110110101" => datar <= "0011100011011001";datai <= "1000110101010010"; --181
        when "0110110110" => datar <= "0011100000100100";datai <= "1000110011111001"; --182
        when "0110110111" => datar <= "0011011101101111";datai <= "1000110010100010"; --183
        when "0110111000" => datar <= "0011011010111010";datai <= "1000110001001011"; --184
        when "0110111001" => datar <= "0011011000000100";datai <= "1000101111110110"; --185
        when "0110111010" => datar <= "0011010101001101";datai <= "1000101110100001"; --186
        when "0110111011" => datar <= "0011010010010110";datai <= "1000101101001110"; --187
        when "0110111100" => datar <= "0011001111011111";datai <= "1000101011111100"; --188
        when "0110111101" => datar <= "0011001100100110";datai <= "1000101010101011"; --189
        when "0110111110" => datar <= "0011001001101110";datai <= "1000101001011011"; --190
        when "0110111111" => datar <= "0011000110110101";datai <= "1000101000001101"; --191
        when "0111000000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "0111000001" => datar <= "0011000001000001";datai <= "1000100101110011"; --193
        when "0111000010" => datar <= "0010111110000111";datai <= "1000100100101000"; --194
        when "0111000011" => datar <= "0010111011001100";datai <= "1000100011011110"; --195
        when "0111000100" => datar <= "0010111000010001";datai <= "1000100010010101"; --196
        when "0111000101" => datar <= "0010110101010101";datai <= "1000100001001101"; --197
        when "0111000110" => datar <= "0010110010011001";datai <= "1000100000000110"; --198
        when "0111000111" => datar <= "0010101111011100";datai <= "1000011111000001"; --199
        when "0111001000" => datar <= "0010101100011111";datai <= "1000011101111100"; --200
        when "0111001001" => datar <= "0010101001100001";datai <= "1000011100111001"; --201
        when "0111001010" => datar <= "0010100110100011";datai <= "1000011011110111"; --202
        when "0111001011" => datar <= "0010100011100101";datai <= "1000011010110110"; --203
        when "0111001100" => datar <= "0010100000100110";datai <= "1000011001110111"; --204
        when "0111001101" => datar <= "0010011101100111";datai <= "1000011000111000"; --205
        when "0111001110" => datar <= "0010011010101000";datai <= "1000010111111011"; --206
        when "0111001111" => datar <= "0010010111101000";datai <= "1000010110111111"; --207
        when "0111010000" => datar <= "0010010100101000";datai <= "1000010110000100"; --208
        when "0111010001" => datar <= "0010010001100111";datai <= "1000010101001010"; --209
        when "0111010010" => datar <= "0010001110100110";datai <= "1000010100010010"; --210
        when "0111010011" => datar <= "0010001011100101";datai <= "1000010011011010"; --211
        when "0111010100" => datar <= "0010001000100011";datai <= "1000010010100100"; --212
        when "0111010101" => datar <= "0010000101100001";datai <= "1000010001101111"; --213
        when "0111010110" => datar <= "0010000010011111";datai <= "1000010000111011"; --214
        when "0111010111" => datar <= "0001111111011101";datai <= "1000010000001000"; --215
        when "0111011000" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "0111011001" => datar <= "0001111001010111";datai <= "1000001110100111"; --217
        when "0111011010" => datar <= "0001110110010011";datai <= "1000001101111000"; --218
        when "0111011011" => datar <= "0001110011001111";datai <= "1000001101001010"; --219
        when "0111011100" => datar <= "0001110000001011";datai <= "1000001100011101"; --220
        when "0111011101" => datar <= "0001101101000111";datai <= "1000001011110010"; --221
        when "0111011110" => datar <= "0001101010000010";datai <= "1000001011000111"; --222
        when "0111011111" => datar <= "0001100110111110";datai <= "1000001010011110"; --223
        when "0111100000" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "0111100001" => datar <= "0001100000110011";datai <= "1000001001010000"; --225
        when "0111100010" => datar <= "0001011101101110";datai <= "1000001000101011"; --226
        when "0111100011" => datar <= "0001011010101000";datai <= "1000001000000110"; --227
        when "0111100100" => datar <= "0001010111100010";datai <= "1000000111100011"; --228
        when "0111100101" => datar <= "0001010100011100";datai <= "1000000111000010"; --229
        when "0111100110" => datar <= "0001010001010101";datai <= "1000000110100001"; --230
        when "0111100111" => datar <= "0001001110001111";datai <= "1000000110000010"; --231
        when "0111101000" => datar <= "0001001011001000";datai <= "1000000101100100"; --232
        when "0111101001" => datar <= "0001001000000001";datai <= "1000000101000111"; --233
        when "0111101010" => datar <= "0001000100111010";datai <= "1000000100101011"; --234
        when "0111101011" => datar <= "0001000001110010";datai <= "1000000100010001"; --235
        when "0111101100" => datar <= "0000111110101011";datai <= "1000000011110111"; --236
        when "0111101101" => datar <= "0000111011100011";datai <= "1000000011011111"; --237
        when "0111101110" => datar <= "0000111000011100";datai <= "1000000011001001"; --238
        when "0111101111" => datar <= "0000110101010100";datai <= "1000000010110011"; --239
        when "0111110000" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "0111110001" => datar <= "0000101111000100";datai <= "1000000010001100"; --241
        when "0111110010" => datar <= "0000101011111011";datai <= "1000000001111010"; --242
        when "0111110011" => datar <= "0000101000110011";datai <= "1000000001101001"; --243
        when "0111110100" => datar <= "0000100101101010";datai <= "1000000001011010"; --244
        when "0111110101" => datar <= "0000100010100010";datai <= "1000000001001100"; --245
        when "0111110110" => datar <= "0000011111011001";datai <= "1000000000111111"; --246
        when "0111110111" => datar <= "0000011100010001";datai <= "1000000000110011"; --247
        when "0111111000" => datar <= "0000011001001000";datai <= "1000000000101000"; --248
        when "0111111001" => datar <= "0000010101111111";datai <= "1000000000011111"; --249
        when "0111111010" => datar <= "0000010010110110";datai <= "1000000000010111"; --250
        when "0111111011" => datar <= "0000001111101101";datai <= "1000000000010000"; --251
        when "0111111100" => datar <= "0000001100100100";datai <= "1000000000001011"; --252
        when "0111111101" => datar <= "0000001001011011";datai <= "1000000000000111"; --253
        when "0111111110" => datar <= "0000000110010010";datai <= "1000000000000011"; --254
        when "0111111111" => datar <= "0000000011001001";datai <= "1000000000000010"; --255
        when "1000000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "1000000001" => datar <= "0111111111111001";datai <= "1111110110100101"; --3
        when "1000000010" => datar <= "0111111111101001";datai <= "1111101101001010"; --6
        when "1000000011" => datar <= "0111111111001101";datai <= "1111100011101111"; --9
        when "1000000100" => datar <= "0111111110100110";datai <= "1111011010010110"; --12
        when "1000000101" => datar <= "0111111101110100";datai <= "1111010000111100"; --15
        when "1000000110" => datar <= "0111111100110111";datai <= "1111000111100100"; --18
        when "1000000111" => datar <= "0111111011101111";datai <= "1110111110001110"; --21
        when "1000001000" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "1000001001" => datar <= "0111111000111110";datai <= "1110101011100100"; --27
        when "1000001010" => datar <= "0111110111010101";datai <= "1110100010010010"; --30
        when "1000001011" => datar <= "0111110101100010";datai <= "1110011001000010"; --33
        when "1000001100" => datar <= "0111110011100011";datai <= "1110001111110101"; --36
        when "1000001101" => datar <= "0111110001011001";datai <= "1110000110101001"; --39
        when "1000001110" => datar <= "0111101111000101";datai <= "1101111101100001"; --42
        when "1000001111" => datar <= "0111101100100110";datai <= "1101110100011011"; --45
        when "1000010000" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "1000010001" => datar <= "0111100111001000";datai <= "1101100010011001"; --51
        when "1000010010" => datar <= "0111100100001001";datai <= "1101011001011101"; --54
        when "1000010011" => datar <= "0111100000111111";datai <= "1101010000100100"; --57
        when "1000010100" => datar <= "0111011101101011";datai <= "1101000111101111"; --60
        when "1000010101" => datar <= "0111011010001101";datai <= "1100111110111111"; --63
        when "1000010110" => datar <= "0111010110100101";datai <= "1100110110010010"; --66
        when "1000010111" => datar <= "0111010010110010";datai <= "1100101101101010"; --69
        when "1000011000" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "1000011001" => datar <= "0111001010101110";datai <= "1100011100100111"; --75
        when "1000011010" => datar <= "0111000110011101";datai <= "1100010100001110"; --78
        when "1000011011" => datar <= "0111000010000011";datai <= "1100001011111001"; --81
        when "1000011100" => datar <= "0110111101011110";datai <= "1100000011101001"; --84
        when "1000011101" => datar <= "0110111000110000";datai <= "1011111011011111"; --87
        when "1000011110" => datar <= "0110110011111000";datai <= "1011110011011011"; --90
        when "1000011111" => datar <= "0110101110110111";datai <= "1011101011011100"; --93
        when "1000100000" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "1000100001" => datar <= "0110100100011001";datai <= "1011011011110001"; --99
        when "1000100010" => datar <= "0110011110111100";datai <= "1011010100000101"; --102
        when "1000100011" => datar <= "0110011001010110";datai <= "1011001100100000"; --105
        when "1000100100" => datar <= "0110010011101000";datai <= "1011000101000001"; --108
        when "1000100101" => datar <= "0110001101110000";datai <= "1010111101101001"; --111
        when "1000100110" => datar <= "0110000111110000";datai <= "1010110110011000"; --114
        when "1000100111" => datar <= "0110000001101000";datai <= "1010101111001110"; --117
        when "1000101000" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "1000101001" => datar <= "0101110100111110";datai <= "1010100001010000"; --123
        when "1000101010" => datar <= "0101101110011100";datai <= "1010011010011100"; --126
        when "1000101011" => datar <= "0101100111110011";datai <= "1010010011110001"; --129
        when "1000101100" => datar <= "0101100001000010";datai <= "1010001101001101"; --132
        when "1000101101" => datar <= "0101011010001010";datai <= "1010000110110001"; --135
        when "1000101110" => datar <= "0101010011001001";datai <= "1010000000011101"; --138
        when "1000101111" => datar <= "0101001100000010";datai <= "1001111010010010"; --141
        when "1000110000" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "1000110001" => datar <= "0100111101011101";datai <= "1001101110010100"; --147
        when "1000110010" => datar <= "0100110110000001";datai <= "1001101000100011"; --150
        when "1000110011" => datar <= "0100101110011101";datai <= "1001100010111010"; --153
        when "1000110100" => datar <= "0100100110110100";datai <= "1001011101011010"; --156
        when "1000110101" => datar <= "0100011111000011";datai <= "1001011000000011"; --159
        when "1000110110" => datar <= "0100010111001101";datai <= "1001010010110110"; --162
        when "1000110111" => datar <= "0100001111010000";datai <= "1001001101110010"; --165
        when "1000111000" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "1000111001" => datar <= "0011111111000101";datai <= "1001000100000101"; --171
        when "1000111010" => datar <= "0011110110111000";datai <= "1000111111011110"; --174
        when "1000111011" => datar <= "0011101110100101";datai <= "1000111011000000"; --177
        when "1000111100" => datar <= "0011100110001100";datai <= "1000110110101100"; --180
        when "1000111101" => datar <= "0011011101101111";datai <= "1000110010100010"; --183
        when "1000111110" => datar <= "0011010101001101";datai <= "1000101110100001"; --186
        when "1000111111" => datar <= "0011001100100110";datai <= "1000101010101011"; --189
        when "1001000000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "1001000001" => datar <= "0010111011001100";datai <= "1000100011011110"; --195
        when "1001000010" => datar <= "0010110010011001";datai <= "1000100000000110"; --198
        when "1001000011" => datar <= "0010101001100001";datai <= "1000011100111001"; --201
        when "1001000100" => datar <= "0010100000100110";datai <= "1000011001110111"; --204
        when "1001000101" => datar <= "0010010111101000";datai <= "1000010110111111"; --207
        when "1001000110" => datar <= "0010001110100110";datai <= "1000010100010010"; --210
        when "1001000111" => datar <= "0010000101100001";datai <= "1000010001101111"; --213
        when "1001001000" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "1001001001" => datar <= "0001110011001111";datai <= "1000001101001010"; --219
        when "1001001010" => datar <= "0001101010000010";datai <= "1000001011000111"; --222
        when "1001001011" => datar <= "0001100000110011";datai <= "1000001001010000"; --225
        when "1001001100" => datar <= "0001010111100010";datai <= "1000000111100011"; --228
        when "1001001101" => datar <= "0001001110001111";datai <= "1000000110000010"; --231
        when "1001001110" => datar <= "0001000100111010";datai <= "1000000100101011"; --234
        when "1001001111" => datar <= "0000111011100011";datai <= "1000000011011111"; --237
        when "1001010000" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "1001010001" => datar <= "0000101000110011";datai <= "1000000001101001"; --243
        when "1001010010" => datar <= "0000011111011001";datai <= "1000000000111111"; --246
        when "1001010011" => datar <= "0000010101111111";datai <= "1000000000011111"; --249
        when "1001010100" => datar <= "0000001100100100";datai <= "1000000000001011"; --252
        when "1001010101" => datar <= "0000000011001001";datai <= "1000000000000010"; --255
        when "1001010110" => datar <= "1111111001101110";datai <= "1000000000000011"; --258
        when "1001010111" => datar <= "1111110000010011";datai <= "1000000000010000"; --261
        when "1001011000" => datar <= "1111100110111000";datai <= "1000000000101000"; --264
        when "1001011001" => datar <= "1111011101011110";datai <= "1000000001001100"; --267
        when "1001011010" => datar <= "1111010100000101";datai <= "1000000001111010"; --270
        when "1001011011" => datar <= "1111001010101100";datai <= "1000000010110011"; --273
        when "1001011100" => datar <= "1111000001010101";datai <= "1000000011110111"; --276
        when "1001011101" => datar <= "1110110111111111";datai <= "1000000101000111"; --279
        when "1001011110" => datar <= "1110101110101011";datai <= "1000000110100001"; --282
        when "1001011111" => datar <= "1110100101011000";datai <= "1000001000000110"; --285
        when "1001100000" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "1001100001" => datar <= "1110010010111001";datai <= "1000001011110010"; --291
        when "1001100010" => datar <= "1110001001101101";datai <= "1000001101111000"; --294
        when "1001100011" => datar <= "1110000000100011";datai <= "1000010000001000"; --297
        when "1001100100" => datar <= "1101110111011101";datai <= "1000010010100100"; --300
        when "1001100101" => datar <= "1101101110011001";datai <= "1000010101001010"; --303
        when "1001100110" => datar <= "1101100101011000";datai <= "1000010111111011"; --306
        when "1001100111" => datar <= "1101011100011011";datai <= "1000011010110110"; --309
        when "1001101000" => datar <= "1101010011100001";datai <= "1000011101111100"; --312
        when "1001101001" => datar <= "1101001010101011";datai <= "1000100001001101"; --315
        when "1001101010" => datar <= "1101000001111001";datai <= "1000100100101000"; --318
        when "1001101011" => datar <= "1100111001001011";datai <= "1000101000001101"; --321
        when "1001101100" => datar <= "1100110000100001";datai <= "1000101011111100"; --324
        when "1001101101" => datar <= "1100100111111100";datai <= "1000101111110110"; --327
        when "1001101110" => datar <= "1100011111011100";datai <= "1000110011111001"; --330
        when "1001101111" => datar <= "1100010111000000";datai <= "1000111000000111"; --333
        when "1001110000" => datar <= "1100001110101010";datai <= "1000111100011110"; --336
        when "1001110001" => datar <= "1100000110011000";datai <= "1001000000111111"; --339
        when "1001110010" => datar <= "1011111110001101";datai <= "1001000101101010"; --342
        when "1001110011" => datar <= "1011110110000110";datai <= "1001001010011111"; --345
        when "1001110100" => datar <= "1011101110000110";datai <= "1001001111011101"; --348
        when "1001110101" => datar <= "1011100110001011";datai <= "1001010100100100"; --351
        when "1001110110" => datar <= "1011011110010111";datai <= "1001011001110101"; --354
        when "1001110111" => datar <= "1011010110101000";datai <= "1001011111001110"; --357
        when "1001111000" => datar <= "1011001111000001";datai <= "1001100100110001"; --360
        when "1001111001" => datar <= "1011000111100000";datai <= "1001101010011101"; --363
        when "1001111010" => datar <= "1011000000000101";datai <= "1001110000010010"; --366
        when "1001111011" => datar <= "1010111000110010";datai <= "1001110110001111"; --369
        when "1001111100" => datar <= "1010110001100101";datai <= "1001111100010101"; --372
        when "1001111101" => datar <= "1010101010100000";datai <= "1010000010100011"; --375
        when "1001111110" => datar <= "1010100011100011";datai <= "1010001000111001"; --378
        when "1001111111" => datar <= "1010011100101101";datai <= "1010001111011000"; --381
        when "1010000000" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "1010000001" => datar <= "1010001111011000";datai <= "1010011100101101"; --387
        when "1010000010" => datar <= "1010001000111001";datai <= "1010100011100011"; --390
        when "1010000011" => datar <= "1010000010100011";datai <= "1010101010100000"; --393
        when "1010000100" => datar <= "1001111100010101";datai <= "1010110001100101"; --396
        when "1010000101" => datar <= "1001110110001111";datai <= "1010111000110010"; --399
        when "1010000110" => datar <= "1001110000010010";datai <= "1011000000000101"; --402
        when "1010000111" => datar <= "1001101010011101";datai <= "1011000111100000"; --405
        when "1010001000" => datar <= "1001100100110001";datai <= "1011001111000001"; --408
        when "1010001001" => datar <= "1001011111001110";datai <= "1011010110101000"; --411
        when "1010001010" => datar <= "1001011001110101";datai <= "1011011110010111"; --414
        when "1010001011" => datar <= "1001010100100100";datai <= "1011100110001011"; --417
        when "1010001100" => datar <= "1001001111011101";datai <= "1011101110000110"; --420
        when "1010001101" => datar <= "1001001010011111";datai <= "1011110110000110"; --423
        when "1010001110" => datar <= "1001000101101010";datai <= "1011111110001101"; --426
        when "1010001111" => datar <= "1001000000111111";datai <= "1100000110011000"; --429
        when "1010010000" => datar <= "1000111100011110";datai <= "1100001110101010"; --432
        when "1010010001" => datar <= "1000111000000111";datai <= "1100010111000000"; --435
        when "1010010010" => datar <= "1000110011111001";datai <= "1100011111011100"; --438
        when "1010010011" => datar <= "1000101111110110";datai <= "1100100111111100"; --441
        when "1010010100" => datar <= "1000101011111100";datai <= "1100110000100001"; --444
        when "1010010101" => datar <= "1000101000001101";datai <= "1100111001001011"; --447
        when "1010010110" => datar <= "1000100100101000";datai <= "1101000001111001"; --450
        when "1010010111" => datar <= "1000100001001101";datai <= "1101001010101011"; --453
        when "1010011000" => datar <= "1000011101111100";datai <= "1101010011100001"; --456
        when "1010011001" => datar <= "1000011010110110";datai <= "1101011100011011"; --459
        when "1010011010" => datar <= "1000010111111011";datai <= "1101100101011000"; --462
        when "1010011011" => datar <= "1000010101001010";datai <= "1101101110011001"; --465
        when "1010011100" => datar <= "1000010010100100";datai <= "1101110111011101"; --468
        when "1010011101" => datar <= "1000010000001000";datai <= "1110000000100011"; --471
        when "1010011110" => datar <= "1000001101111000";datai <= "1110001001101101"; --474
        when "1010011111" => datar <= "1000001011110010";datai <= "1110010010111001"; --477
        when "1010100000" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "1010100001" => datar <= "1000001000000110";datai <= "1110100101011000"; --483
        when "1010100010" => datar <= "1000000110100001";datai <= "1110101110101011"; --486
        when "1010100011" => datar <= "1000000101000111";datai <= "1110110111111111"; --489
        when "1010100100" => datar <= "1000000011110111";datai <= "1111000001010101"; --492
        when "1010100101" => datar <= "1000000010110011";datai <= "1111001010101100"; --495
        when "1010100110" => datar <= "1000000001111010";datai <= "1111010100000101"; --498
        when "1010100111" => datar <= "1000000001001100";datai <= "1111011101011110"; --501
        when "1010101000" => datar <= "1000000000101000";datai <= "1111100110111000"; --504
        when "1010101001" => datar <= "1000000000010000";datai <= "1111110000010011"; --507
        when "1010101010" => datar <= "1000000000000011";datai <= "1111111001101110"; --510
        when "1010101011" => datar <= "1000000000000010";datai <= "0000000011001001"; --513
        when "1010101100" => datar <= "1000000000001011";datai <= "0000001100100100"; --516
        when "1010101101" => datar <= "1000000000011111";datai <= "0000010101111111"; --519
        when "1010101110" => datar <= "1000000000111111";datai <= "0000011111011001"; --522
        when "1010101111" => datar <= "1000000001101001";datai <= "0000101000110011"; --525
        when "1010110000" => datar <= "1000000010011111";datai <= "0000110010001100"; --528
        when "1010110001" => datar <= "1000000011011111";datai <= "0000111011100011"; --531
        when "1010110010" => datar <= "1000000100101011";datai <= "0001000100111010"; --534
        when "1010110011" => datar <= "1000000110000010";datai <= "0001001110001111"; --537
        when "1010110100" => datar <= "1000000111100011";datai <= "0001010111100010"; --540
        when "1010110101" => datar <= "1000001001010000";datai <= "0001100000110011"; --543
        when "1010110110" => datar <= "1000001011000111";datai <= "0001101010000010"; --546
        when "1010110111" => datar <= "1000001101001010";datai <= "0001110011001111"; --549
        when "1010111000" => datar <= "1000001111010111";datai <= "0001111100011010"; --552
        when "1010111001" => datar <= "1000010001101111";datai <= "0010000101100001"; --555
        when "1010111010" => datar <= "1000010100010010";datai <= "0010001110100110"; --558
        when "1010111011" => datar <= "1000010110111111";datai <= "0010010111101000"; --561
        when "1010111100" => datar <= "1000011001110111";datai <= "0010100000100110"; --564
        when "1010111101" => datar <= "1000011100111001";datai <= "0010101001100001"; --567
        when "1010111110" => datar <= "1000100000000110";datai <= "0010110010011001"; --570
        when "1010111111" => datar <= "1000100011011110";datai <= "0010111011001100"; --573
        when "1011000000" => datar <= "1000100110111111";datai <= "0011000011111011"; --576
        when "1011000001" => datar <= "1000101010101011";datai <= "0011001100100110"; --579
        when "1011000010" => datar <= "1000101110100001";datai <= "0011010101001101"; --582
        when "1011000011" => datar <= "1000110010100010";datai <= "0011011101101111"; --585
        when "1011000100" => datar <= "1000110110101100";datai <= "0011100110001100"; --588
        when "1011000101" => datar <= "1000111011000000";datai <= "0011101110100101"; --591
        when "1011000110" => datar <= "1000111111011110";datai <= "0011110110111000"; --594
        when "1011000111" => datar <= "1001000100000101";datai <= "0011111111000101"; --597
        when "1011001000" => datar <= "1001001000110111";datai <= "0100000111001110"; --600
        when "1011001001" => datar <= "1001001101110010";datai <= "0100001111010000"; --603
        when "1011001010" => datar <= "1001010010110110";datai <= "0100010111001101"; --606
        when "1011001011" => datar <= "1001011000000011";datai <= "0100011111000011"; --609
        when "1011001100" => datar <= "1001011101011010";datai <= "0100100110110100"; --612
        when "1011001101" => datar <= "1001100010111010";datai <= "0100101110011101"; --615
        when "1011001110" => datar <= "1001101000100011";datai <= "0100110110000001"; --618
        when "1011001111" => datar <= "1001101110010100";datai <= "0100111101011101"; --621
        when "1011010000" => datar <= "1001110100001111";datai <= "0101000100110011"; --624
        when "1011010001" => datar <= "1001111010010010";datai <= "0101001100000010"; --627
        when "1011010010" => datar <= "1010000000011101";datai <= "0101010011001001"; --630
        when "1011010011" => datar <= "1010000110110001";datai <= "0101011010001010"; --633
        when "1011010100" => datar <= "1010001101001101";datai <= "0101100001000010"; --636
        when "1011010101" => datar <= "1010010011110001";datai <= "0101100111110011"; --639
        when "1011010110" => datar <= "1010011010011100";datai <= "0101101110011100"; --642
        when "1011010111" => datar <= "1010100001010000";datai <= "0101110100111110"; --645
        when "1011011000" => datar <= "1010101000001011";datai <= "0101111011010111"; --648
        when "1011011001" => datar <= "1010101111001110";datai <= "0110000001101000"; --651
        when "1011011010" => datar <= "1010110110011000";datai <= "0110000111110000"; --654
        when "1011011011" => datar <= "1010111101101001";datai <= "0110001101110000"; --657
        when "1011011100" => datar <= "1011000101000001";datai <= "0110010011101000"; --660
        when "1011011101" => datar <= "1011001100100000";datai <= "0110011001010110"; --663
        when "1011011110" => datar <= "1011010100000101";datai <= "0110011110111100"; --666
        when "1011011111" => datar <= "1011011011110001";datai <= "0110100100011001"; --669
        when "1011100000" => datar <= "1011100011100100";datai <= "0110101001101101"; --672
        when "1011100001" => datar <= "1011101011011100";datai <= "0110101110110111"; --675
        when "1011100010" => datar <= "1011110011011011";datai <= "0110110011111000"; --678
        when "1011100011" => datar <= "1011111011011111";datai <= "0110111000110000"; --681
        when "1011100100" => datar <= "1100000011101001";datai <= "0110111101011110"; --684
        when "1011100101" => datar <= "1100001011111001";datai <= "0111000010000011"; --687
        when "1011100110" => datar <= "1100010100001110";datai <= "0111000110011101"; --690
        when "1011100111" => datar <= "1100011100100111";datai <= "0111001010101110"; --693
        when "1011101000" => datar <= "1100100101000110";datai <= "0111001110110101"; --696
        when "1011101001" => datar <= "1100101101101010";datai <= "0111010010110010"; --699
        when "1011101010" => datar <= "1100110110010010";datai <= "0111010110100101"; --702
        when "1011101011" => datar <= "1100111110111111";datai <= "0111011010001101"; --705
        when "1011101100" => datar <= "1101000111101111";datai <= "0111011101101011"; --708
        when "1011101101" => datar <= "1101010000100100";datai <= "0111100000111111"; --711
        when "1011101110" => datar <= "1101011001011101";datai <= "0111100100001001"; --714
        when "1011101111" => datar <= "1101100010011001";datai <= "0111100111001000"; --717
        when "1011110000" => datar <= "1101101011011000";datai <= "0111101001111100"; --720
        when "1011110001" => datar <= "1101110100011011";datai <= "0111101100100110"; --723
        when "1011110010" => datar <= "1101111101100001";datai <= "0111101111000101"; --726
        when "1011110011" => datar <= "1110000110101001";datai <= "0111110001011001"; --729
        when "1011110100" => datar <= "1110001111110101";datai <= "0111110011100011"; --732
        when "1011110101" => datar <= "1110011001000010";datai <= "0111110101100010"; --735
        when "1011110110" => datar <= "1110100010010010";datai <= "0111110111010101"; --738
        when "1011110111" => datar <= "1110101011100100";datai <= "0111111000111110"; --741
        when "1011111000" => datar <= "1110110100111000";datai <= "0111111010011100"; --744
        when "1011111001" => datar <= "1110111110001110";datai <= "0111111011101111"; --747
        when "1011111010" => datar <= "1111000111100100";datai <= "0111111100110111"; --750
        when "1011111011" => datar <= "1111010000111100";datai <= "0111111101110100"; --753
        when "1011111100" => datar <= "1111011010010110";datai <= "0111111110100110"; --756
        when "1011111101" => datar <= "1111100011101111";datai <= "0111111111001101"; --759
        when "1011111110" => datar <= "1111101101001010";datai <= "0111111111101001"; --762
        when "1011111111" => datar <= "1111110110100101";datai <= "0111111111111001"; --765
           when "1100000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100000111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100001111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100010111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100011111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100100111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100101111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1100111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101000111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101001111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101010111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101011111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101100111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101101111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1101111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110000111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110001111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110010111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110011111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110100111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110101111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1110111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111000111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111001111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111010111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111011111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111100111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111101111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "1111111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when others => for i in data_width-1 downto 0 loop
            datar(i)<='0';datai(i)<='0';end loop;
    end case;

    end if;

end process;
END behavior;
