000000 => x"cafe",
000001 => x"03d3",
000002 => x"9c97",
000003 => x"6666",
000004 => x"7431",
000005 => x"3238",
000006 => x"2e61",
000007 => x"736d",
000008 => x"bc0b",
000009 => x"bc04",
000010 => x"bc03",
000011 => x"bc02",
000012 => x"bc01",
000013 => x"be73",
000014 => x"c578",
000015 => x"c906",
000016 => x"be7f",
000017 => x"be6f",
000018 => x"bc00",
000019 => x"c724",
000020 => x"cb07",
000021 => x"c114",
000022 => x"c907",
000023 => x"be78",
000024 => x"c47f",
000025 => x"ec0b",
000026 => x"c002",
000027 => x"ec0c",
000028 => x"c400",
000029 => x"c800",
000030 => x"c7e6",
000031 => x"cb82",
000032 => x"3474",
000033 => x"6c6a",
000034 => x"c6f8",
000035 => x"ca83",
000036 => x"c578",
000037 => x"c904",
000038 => x"29b3",
000039 => x"785a",
000040 => x"c080",
000041 => x"526a",
000042 => x"c7c4",
000043 => x"cb82",
000044 => x"3474",
000045 => x"01b1",
000046 => x"c400",
000047 => x"c800",
000048 => x"1838",
000049 => x"85f6",
000050 => x"586a",
000051 => x"2ad5",
000052 => x"ec5a",
000053 => x"c478",
000054 => x"c804",
000055 => x"c480",
000056 => x"c880",
000057 => x"c578",
000058 => x"c902",
000059 => x"be5e",
000060 => x"ee02",
000061 => x"be1a",
000062 => x"be42",
000063 => x"c6f8",
000064 => x"ca84",
000065 => x"c580",
000066 => x"c980",
000067 => x"7a5a",
000068 => x"be13",
000069 => x"c0a0",
000070 => x"be07",
000071 => x"7a5a",
000072 => x"be0f",
000073 => x"be37",
000074 => x"05b9",
000075 => x"85f8",
000076 => x"bc00",
000077 => x"ec22",
000078 => x"dc05",
000079 => x"b9fe",
000080 => x"ed18",
000081 => x"3470",
000082 => x"ec20",
000083 => x"dc8f",
000084 => x"b9fe",
000085 => x"c800",
000086 => x"3470",
000087 => x"6c6a",
000088 => x"6cea",
000089 => x"6d6a",
000090 => x"6dea",
000091 => x"6e6a",
000092 => x"6fea",
000093 => x"3d42",
000094 => x"3d22",
000095 => x"3d22",
000096 => x"3d22",
000097 => x"be15",
000098 => x"bfeb",
000099 => x"3d40",
000100 => x"be12",
000101 => x"bfe8",
000102 => x"3d45",
000103 => x"3d25",
000104 => x"3d25",
000105 => x"3d25",
000106 => x"be0c",
000107 => x"bfe2",
000108 => x"0140",
000109 => x"be09",
000110 => x"bfdf",
000111 => x"5bea",
000112 => x"5a6a",
000113 => x"59ea",
000114 => x"596a",
000115 => x"58ea",
000116 => x"586a",
000117 => x"3470",
000118 => x"c08f",
000119 => x"2121",
000120 => x"c089",
000121 => x"181a",
000122 => x"8803",
000123 => x"c0b0",
000124 => x"bc02",
000125 => x"c0b7",
000126 => x"0892",
000127 => x"3470",
000128 => x"6c6a",
000129 => x"6cea",
000130 => x"6d6a",
000131 => x"6fea",
000132 => x"0170",
000133 => x"c08d",
000134 => x"bfc7",
000135 => x"c08a",
000136 => x"03a0",
000137 => x"bfc4",
000138 => x"5bea",
000139 => x"596a",
000140 => x"58ea",
000141 => x"586a",
000142 => x"3470",
000143 => x"0270",
000144 => x"7829",
000145 => x"c080",
000146 => x"ccff",
000147 => x"2081",
000148 => x"3c98",
000149 => x"8003",
000150 => x"bfb7",
000151 => x"bdf9",
000152 => x"3440",
000153 => x"6eea",
000154 => x"6e6a",
000155 => x"6dea",
000156 => x"6d6a",
000157 => x"6cea",
000158 => x"6c6a",
000159 => x"6fea",
000160 => x"c3b6",
000161 => x"cb82",
000162 => x"447e",
000163 => x"44fa",
000164 => x"457c",
000165 => x"2800",
000166 => x"3c95",
000167 => x"3419",
000168 => x"8003",
000169 => x"0001",
000170 => x"bdfc",
000171 => x"c3b6",
000172 => x"cb82",
000173 => x"5478",
000174 => x"c3b6",
000175 => x"cb82",
000176 => x"c281",
000177 => x"56fa",
000178 => x"56fc",
000179 => x"56fe",
000180 => x"c3be",
000181 => x"cb82",
000182 => x"c280",
000183 => x"56f8",
000184 => x"c3ba",
000185 => x"cb82",
000186 => x"40fa",
000187 => x"5178",
000188 => x"0521",
000189 => x"c204",
000190 => x"3e44",
000191 => x"0499",
000192 => x"85fe",
000193 => x"f124",
000194 => x"557c",
000195 => x"c3b6",
000196 => x"cb82",
000197 => x"427e",
000198 => x"50fa",
000199 => x"517e",
000200 => x"41fc",
000201 => x"0521",
000202 => x"3d24",
000203 => x"3d24",
000204 => x"0932",
000205 => x"c3be",
000206 => x"cb82",
000207 => x"5078",
000208 => x"0804",
000209 => x"c182",
000210 => x"3db4",
000211 => x"0499",
000212 => x"85fe",
000213 => x"0883",
000214 => x"c3c0",
000215 => x"cb82",
000216 => x"5478",
000217 => x"54fa",
000218 => x"557c",
000219 => x"0180",
000220 => x"0210",
000221 => x"02a0",
000222 => x"6dea",
000223 => x"6e6a",
000224 => x"5038",
000225 => x"50ba",
000226 => x"5148",
000227 => x"51ca",
000228 => x"5258",
000229 => x"52da",
000230 => x"be45",
000231 => x"5aea",
000232 => x"5a6a",
000233 => x"5558",
000234 => x"55da",
000235 => x"5448",
000236 => x"54ca",
000237 => x"c3be",
000238 => x"cb82",
000239 => x"5078",
000240 => x"c084",
000241 => x"0801",
000242 => x"5478",
000243 => x"c3b6",
000244 => x"cb82",
000245 => x"507a",
000246 => x"517e",
000247 => x"c081",
000248 => x"0409",
000249 => x"8003",
000250 => x"3c94",
000251 => x"bdfd",
000252 => x"181a",
000253 => x"0121",
000254 => x"557e",
000255 => x"85c4",
000256 => x"c101",
000257 => x"557e",
000258 => x"c3b6",
000259 => x"cb82",
000260 => x"407a",
000261 => x"50fa",
000262 => x"517c",
000263 => x"3c05",
000264 => x"0499",
000265 => x"85fe",
000266 => x"180a",
000267 => x"0121",
000268 => x"557c",
000269 => x"85ab",
000270 => x"c101",
000271 => x"557c",
000272 => x"c3b6",
000273 => x"cb82",
000274 => x"5078",
000275 => x"50fa",
000276 => x"1809",
000277 => x"0091",
000278 => x"54fa",
000279 => x"85a1",
000280 => x"5bea",
000281 => x"586a",
000282 => x"58ea",
000283 => x"596a",
000284 => x"59ea",
000285 => x"5a6a",
000286 => x"5aea",
000287 => x"3470",
000288 => x"0000",
000289 => x"0000",
000290 => x"0000",
000291 => x"0000",
000292 => x"0000",
000293 => x"0000",
000294 => x"0000",
000295 => x"0000",
000296 => x"0000",
000297 => x"0000",
000298 => x"0000",
000299 => x"6fea",
000300 => x"6c6a",
000301 => x"6cea",
000302 => x"c7bc",
000303 => x"cb82",
000304 => x"f042",
000305 => x"f0ca",
000306 => x"3c0c",
000307 => x"3c92",
000308 => x"3c0c",
000309 => x"3c92",
000310 => x"54f8",
000311 => x"f043",
000312 => x"f0cb",
000313 => x"3c0c",
000314 => x"3c92",
000315 => x"3c0c",
000316 => x"3c92",
000317 => x"54fa",
000318 => x"f052",
000319 => x"f0da",
000320 => x"3c0c",
000321 => x"3c92",
000322 => x"3c0c",
000323 => x"3c92",
000324 => x"54fc",
000325 => x"f053",
000326 => x"f0db",
000327 => x"3c0c",
000328 => x"3c92",
000329 => x"3c0c",
000330 => x"3c92",
000331 => x"54fe",
000332 => x"58ea",
000333 => x"586a",
000334 => x"5178",
000335 => x"51fe",
000336 => x"090a",
000337 => x"15a3",
000338 => x"6dea",
000339 => x"517a",
000340 => x"51fc",
000341 => x"091a",
000342 => x"0da3",
000343 => x"6dea",
000344 => x"5178",
000345 => x"51fe",
000346 => x"110a",
000347 => x"0da3",
000348 => x"6dea",
000349 => x"517a",
000350 => x"51fc",
000351 => x"111a",
000352 => x"15a3",
000353 => x"596a",
000354 => x"58ea",
000355 => x"586a",
000356 => x"5bea",
000357 => x"3470",
000358 => x"0000",
000359 => x"0000",
000360 => x"0000",
000361 => x"0000",
000362 => x"6dea",
000363 => x"6e6a",
000364 => x"6eea",
000365 => x"2ad5",
000366 => x"3dbd",
000367 => x"3ed6",
000368 => x"0649",
000369 => x"85fd",
000370 => x"3ed4",
000371 => x"3ed4",
000372 => x"0aa5",
000373 => x"5458",
000374 => x"54da",
000375 => x"5aea",
000376 => x"5a6a",
000377 => x"59ea",
000378 => x"3470",
000379 => x"6cea",
000380 => x"2891",
000381 => x"3c0d",
000382 => x"8003",
000383 => x"0091",
000384 => x"bdfd",
000385 => x"0010",
000386 => x"58ea",
000387 => x"3470",
000388 => x"4000",
000389 => x"0000",
000390 => x"3fec",
000391 => x"0323",
000392 => x"3fb1",
000393 => x"0645",
000394 => x"3f4e",
000395 => x"0964",
000396 => x"3ec5",
000397 => x"0c7c",
000398 => x"3e14",
000399 => x"0f8c",
000400 => x"3d3e",
000401 => x"1294",
000402 => x"3c42",
000403 => x"158f",
000404 => x"3b20",
000405 => x"187d",
000406 => x"39da",
000407 => x"1b5d",
000408 => x"3871",
000409 => x"1e2b",
000410 => x"36e5",
000411 => x"20e7",
000412 => x"3536",
000413 => x"238e",
000414 => x"3367",
000415 => x"261f",
000416 => x"3179",
000417 => x"2899",
000418 => x"2f6b",
000419 => x"2afa",
000420 => x"2d41",
000421 => x"2d41",
000422 => x"2afa",
000423 => x"2f6b",
000424 => x"2899",
000425 => x"3179",
000426 => x"261f",
000427 => x"3367",
000428 => x"238e",
000429 => x"3536",
000430 => x"20e7",
000431 => x"36e5",
000432 => x"1e2b",
000433 => x"3871",
000434 => x"1b5d",
000435 => x"39da",
000436 => x"187d",
000437 => x"3b20",
000438 => x"158f",
000439 => x"3c42",
000440 => x"1294",
000441 => x"3d3e",
000442 => x"0f8c",
000443 => x"3e14",
000444 => x"0c7c",
000445 => x"3ec5",
000446 => x"0964",
000447 => x"3f4e",
000448 => x"0645",
000449 => x"3fb1",
000450 => x"0323",
000451 => x"3fec",
000452 => x"0000",
000453 => x"4000",
000454 => x"fcdd",
000455 => x"3fec",
000456 => x"f9bb",
000457 => x"3fb1",
000458 => x"f69c",
000459 => x"3f4e",
000460 => x"f384",
000461 => x"3ec5",
000462 => x"f074",
000463 => x"3e14",
000464 => x"ed6c",
000465 => x"3d3e",
000466 => x"ea71",
000467 => x"3c42",
000468 => x"e783",
000469 => x"3b20",
000470 => x"e4a3",
000471 => x"39da",
000472 => x"e1d5",
000473 => x"3871",
000474 => x"df19",
000475 => x"36e5",
000476 => x"dc72",
000477 => x"3536",
000478 => x"d9e1",
000479 => x"3367",
000480 => x"d767",
000481 => x"3179",
000482 => x"d506",
000483 => x"2f6b",
000484 => x"d2bf",
000485 => x"2d41",
000486 => x"d095",
000487 => x"2afa",
000488 => x"ce87",
000489 => x"2899",
000490 => x"cc99",
000491 => x"261f",
000492 => x"caca",
000493 => x"238e",
000494 => x"c91b",
000495 => x"20e7",
000496 => x"c78f",
000497 => x"1e2b",
000498 => x"c626",
000499 => x"1b5d",
000500 => x"c4e0",
000501 => x"187d",
000502 => x"c3be",
000503 => x"158f",
000504 => x"c2c2",
000505 => x"1294",
000506 => x"c1ec",
000507 => x"0f8c",
000508 => x"c13b",
000509 => x"0c7c",
000510 => x"c0b2",
000511 => x"0964",
000512 => x"c04f",
000513 => x"0645",
000514 => x"c014",
000515 => x"0323",
000516 => x"0400",
000517 => x"0000",
000518 => x"0000",
000519 => x"0000",
000520 => x"0400",
000521 => x"0000",
000522 => x"0000",
000523 => x"0000",
000524 => x"0400",
000525 => x"0000",
000526 => x"0000",
000527 => x"0000",
000528 => x"0400",
000529 => x"0000",
000530 => x"0000",
000531 => x"0000",
000532 => x"0400",
000533 => x"0000",
000534 => x"0000",
000535 => x"0000",
000536 => x"0400",
000537 => x"0000",
000538 => x"0000",
000539 => x"0000",
000540 => x"0400",
000541 => x"0000",
000542 => x"0000",
000543 => x"0000",
000544 => x"0400",
000545 => x"0000",
000546 => x"0000",
000547 => x"0000",
000548 => x"0400",
000549 => x"0000",
000550 => x"0000",
000551 => x"0000",
000552 => x"0400",
000553 => x"0000",
000554 => x"0000",
000555 => x"0000",
000556 => x"0400",
000557 => x"0000",
000558 => x"0000",
000559 => x"0000",
000560 => x"0400",
000561 => x"0000",
000562 => x"0000",
000563 => x"0000",
000564 => x"0400",
000565 => x"0000",
000566 => x"0000",
000567 => x"0000",
000568 => x"0400",
000569 => x"0000",
000570 => x"0000",
000571 => x"0000",
000572 => x"0400",
000573 => x"0000",
000574 => x"0000",
000575 => x"0000",
000576 => x"0400",
000577 => x"0000",
000578 => x"0000",
000579 => x"0000",
000580 => x"0400",
000581 => x"0000",
000582 => x"0000",
000583 => x"0000",
000584 => x"0400",
000585 => x"0000",
000586 => x"0000",
000587 => x"0000",
000588 => x"0400",
000589 => x"0000",
000590 => x"0000",
000591 => x"0000",
000592 => x"0400",
000593 => x"0000",
000594 => x"0000",
000595 => x"0000",
000596 => x"0400",
000597 => x"0000",
000598 => x"0000",
000599 => x"0000",
000600 => x"0400",
000601 => x"0000",
000602 => x"0000",
000603 => x"0000",
000604 => x"0400",
000605 => x"0000",
000606 => x"0000",
000607 => x"0000",
000608 => x"0400",
000609 => x"0000",
000610 => x"0000",
000611 => x"0000",
000612 => x"0400",
000613 => x"0000",
000614 => x"0000",
000615 => x"0000",
000616 => x"0400",
000617 => x"0000",
000618 => x"0000",
000619 => x"0000",
000620 => x"0400",
000621 => x"0000",
000622 => x"0000",
000623 => x"0000",
000624 => x"0400",
000625 => x"0000",
000626 => x"0000",
000627 => x"0000",
000628 => x"0400",
000629 => x"0000",
000630 => x"0000",
000631 => x"0000",
000632 => x"0400",
000633 => x"0000",
000634 => x"0000",
000635 => x"0000",
000636 => x"0400",
000637 => x"0000",
000638 => x"0000",
000639 => x"0000",
000640 => x"0400",
000641 => x"0000",
000642 => x"0000",
000643 => x"0000",
000644 => x"0000",
000645 => x"0000",
000646 => x"0000",
000647 => x"0000",
000648 => x"0000",
000649 => x"0000",
000650 => x"0000",
000651 => x"0000",
000652 => x"0000",
000653 => x"0000",
000654 => x"0000",
000655 => x"0000",
000656 => x"0000",
000657 => x"0000",
000658 => x"0000",
000659 => x"0000",
000660 => x"0000",
000661 => x"0000",
000662 => x"0000",
000663 => x"0000",
000664 => x"0000",
000665 => x"0000",
000666 => x"0000",
000667 => x"0000",
000668 => x"0000",
000669 => x"0000",
000670 => x"0000",
000671 => x"0000",
000672 => x"0000",
000673 => x"0000",
000674 => x"0000",
000675 => x"0000",
000676 => x"0000",
000677 => x"0000",
000678 => x"0000",
000679 => x"0000",
000680 => x"0000",
000681 => x"0000",
000682 => x"0000",
000683 => x"0000",
000684 => x"0000",
000685 => x"0000",
000686 => x"0000",
000687 => x"0000",
000688 => x"0000",
000689 => x"0000",
000690 => x"0000",
000691 => x"0000",
000692 => x"0000",
000693 => x"0000",
000694 => x"0000",
000695 => x"0000",
000696 => x"0000",
000697 => x"0000",
000698 => x"0000",
000699 => x"0000",
000700 => x"0000",
000701 => x"0000",
000702 => x"0000",
000703 => x"0000",
000704 => x"0000",
000705 => x"0000",
000706 => x"0000",
000707 => x"0000",
000708 => x"0000",
000709 => x"0000",
000710 => x"0000",
000711 => x"0000",
000712 => x"0000",
000713 => x"0000",
000714 => x"0000",
000715 => x"0000",
000716 => x"0000",
000717 => x"0000",
000718 => x"0000",
000719 => x"0000",
000720 => x"0000",
000721 => x"0000",
000722 => x"0000",
000723 => x"0000",
000724 => x"0000",
000725 => x"0000",
000726 => x"0000",
000727 => x"0000",
000728 => x"0000",
000729 => x"0000",
000730 => x"0000",
000731 => x"0000",
000732 => x"0000",
000733 => x"0000",
000734 => x"0000",
000735 => x"0000",
000736 => x"0000",
000737 => x"0000",
000738 => x"0000",
000739 => x"0000",
000740 => x"0000",
000741 => x"0000",
000742 => x"0000",
000743 => x"0000",
000744 => x"0000",
000745 => x"0000",
000746 => x"0000",
000747 => x"0000",
000748 => x"0000",
000749 => x"0000",
000750 => x"0000",
000751 => x"0000",
000752 => x"0000",
000753 => x"0000",
000754 => x"0000",
000755 => x"0000",
000756 => x"0000",
000757 => x"0000",
000758 => x"0000",
000759 => x"0000",
000760 => x"0000",
000761 => x"0000",
000762 => x"0000",
000763 => x"0000",
000764 => x"0000",
000765 => x"0000",
000766 => x"0000",
000767 => x"0000",
000768 => x"0000",
000769 => x"0000",
000770 => x"0000",
000771 => x"0000",
000772 => x"0000",
000773 => x"0000",
000774 => x"0000",
000775 => x"0000",
000776 => x"0000",
000777 => x"0000",
000778 => x"0000",
000779 => x"0000",
000780 => x"0000",
000781 => x"0000",
000782 => x"0000",
000783 => x"0000",
000784 => x"0000",
000785 => x"0000",
000786 => x"0000",
000787 => x"0000",
000788 => x"0000",
000789 => x"0000",
000790 => x"0000",
000791 => x"0000",
000792 => x"0000",
000793 => x"0000",
000794 => x"0000",
000795 => x"0000",
000796 => x"0000",
000797 => x"0000",
000798 => x"0000",
000799 => x"0000",
000800 => x"0000",
000801 => x"0000",
000802 => x"0000",
000803 => x"0000",
000804 => x"0000",
000805 => x"0000",
000806 => x"0000",
000807 => x"0000",
000808 => x"0000",
000809 => x"0000",
000810 => x"0000",
000811 => x"0000",
000812 => x"0000",
000813 => x"0000",
000814 => x"0000",
000815 => x"0000",
000816 => x"0000",
000817 => x"0000",
000818 => x"0000",
000819 => x"0000",
000820 => x"0000",
000821 => x"0000",
000822 => x"0000",
000823 => x"0000",
000824 => x"0000",
000825 => x"0000",
000826 => x"0000",
000827 => x"0000",
000828 => x"0000",
000829 => x"0000",
000830 => x"0000",
000831 => x"0000",
000832 => x"0000",
000833 => x"0000",
000834 => x"0000",
000835 => x"0000",
000836 => x"0000",
000837 => x"0000",
000838 => x"0000",
000839 => x"0000",
000840 => x"0000",
000841 => x"0000",
000842 => x"0000",
000843 => x"0000",
000844 => x"0000",
000845 => x"0000",
000846 => x"0000",
000847 => x"0000",
000848 => x"0000",
000849 => x"0000",
000850 => x"0000",
000851 => x"0000",
000852 => x"0000",
000853 => x"0000",
000854 => x"0000",
000855 => x"0000",
000856 => x"0000",
000857 => x"0000",
000858 => x"0000",
000859 => x"0000",
000860 => x"0000",
000861 => x"0000",
000862 => x"0000",
000863 => x"0000",
000864 => x"0000",
000865 => x"0000",
000866 => x"0000",
000867 => x"0000",
000868 => x"0000",
000869 => x"0000",
000870 => x"0000",
000871 => x"0000",
000872 => x"0000",
000873 => x"0000",
000874 => x"0000",
000875 => x"0000",
000876 => x"0000",
000877 => x"0000",
000878 => x"0000",
000879 => x"0000",
000880 => x"0000",
000881 => x"0000",
000882 => x"0000",
000883 => x"0000",
000884 => x"0000",
000885 => x"0000",
000886 => x"0000",
000887 => x"0000",
000888 => x"0000",
000889 => x"0000",
000890 => x"0000",
000891 => x"0000",
000892 => x"0000",
000893 => x"0000",
000894 => x"0000",
000895 => x"0000",
000896 => x"0000",
000897 => x"0000",
000898 => x"0000",
000899 => x"0000",
000900 => x"4578",
000901 => x"6365",
000902 => x"7074",
000903 => x"696f",
000904 => x"6e2f",
000905 => x"696e",
000906 => x"7465",
000907 => x"7272",
000908 => x"7570",
000909 => x"7420",
000910 => x"6572",
000911 => x"726f",
000912 => x"7221",
000913 => x"0000",
000914 => x"436f",
000915 => x"6d70",
000916 => x"7574",
000917 => x"696e",
000918 => x"6720",
000919 => x"4646",
000920 => x"542e",
000921 => x"2e2e",
000922 => x"2000",
000923 => x"0000",
000924 => x"0000",
000925 => x"0000",
000926 => x"0000",
000927 => x"0000",
000928 => x"0000",
000929 => x"0000",
000930 => x"0000",
000931 => x"0000",
000932 => x"0000",
000933 => x"0000",
000934 => x"0000",
000935 => x"0000",
000936 => x"0000",
000937 => x"0000",
000938 => x"0000",
000939 => x"0000",
000940 => x"0000",
000941 => x"0000",
000942 => x"0000",
000943 => x"0000",
000944 => x"0000",
000945 => x"0000",
000946 => x"0000",
000947 => x"0000",
000948 => x"0000",
000949 => x"0000",
000950 => x"0000",
000951 => x"0000",
000952 => x"0000",
000953 => x"0000",
000954 => x"0000",
000955 => x"0000",
000956 => x"0000",
000957 => x"0000",
000958 => x"0000",
000959 => x"0000",
000960 => x"0000",
000961 => x"0000",
000962 => x"0000",
000963 => x"0000",
000964 => x"0000",
000965 => x"0000",
000966 => x"0000",
000967 => x"0000",
000968 => x"0000",
000969 => x"0000",
000970 => x"0000",
000971 => x"0000",
000972 => x"0000",
000973 => x"0000",
000974 => x"0000",
000975 => x"0000",
000976 => x"0000",
000977 => x"0000",
000978 => x"0000",
000979 => x"0000",
000980 => x"0000",
000981 => x"0000",
000982 => x"0000",
000983 => x"0000",
000984 => x"0000",
000985 => x"0000",
000986 => x"0000",
others => x"0000"