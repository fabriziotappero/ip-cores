-------------------------------------------------------------------------------
--
-- Parametrizable, generic RAM with enable.
--
-- $Id: generic_ram_ena-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration generic_ram_ena_rtl_c0 of generic_ram_ena is

  for rtl
  end for;

end generic_ram_ena_rtl_c0;
