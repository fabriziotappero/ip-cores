-- Rom file for twiddle factors 
-- ../../../rtl/vhdl/WISHBONE_FFT/rom2.vhd contains 256 points of 16 width 
--  for a 1024 point fft.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;


ENTITY rom2 IS
         GENERIC(
        data_width : integer :=16;
        address_width : integer :=8
    );
    PORT(
        clk :in std_logic;
        address :in std_logic_vector (7      downto 0);
        datar : OUT std_logic_vector (data_width-1 DOWNTO 0) ;
        datai : OUT std_logic_vector (data_width-1 DOWNTO 0)
    );
end rom2;
ARCHITECTURE behavior OF rom2 IS

 BEGIN

process (address,clk)
begin
    	if(rising_edge(clk)) then 
 case address is
        when "00000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "00000001" => datar <= "0111111111011000";datai <= "1111100110111000"; --8
        when "00000010" => datar <= "0111111101100001";datai <= "1111001101110100"; --16
        when "00000011" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "00000100" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "00000101" => datar <= "0111110000101001";datai <= "1110000011100110"; --40
        when "00000110" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "00000111" => datar <= "0111100010000100";datai <= "1101010011100001"; --56
        when "00001000" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "00001001" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "00001010" => datar <= "0111000011100010";datai <= "1100001110101010"; --80
        when "00001011" => datar <= "0110110111001001";datai <= "1011111000110010"; --88
        when "00001100" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "00001101" => datar <= "0110011011001111";datai <= "1011001111000001"; --104
        when "00001110" => datar <= "0110001011110001";datai <= "1010111011001101"; --112
        when "00001111" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "00010000" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "00010001" => datar <= "0101010111110101";datai <= "1010000100101001"; --136
        when "00010010" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "00010011" => datar <= "0100110000111111";datai <= "1001100100110001"; --152
        when "00010100" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "00010101" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "00010110" => datar <= "0011110001010110";datai <= "1000111100011110"; --176
        when "00010111" => datar <= "0011011010111010";datai <= "1000110001001011"; --184
        when "00011000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "00011001" => datar <= "0010101100011111";datai <= "1000011101111100"; --200
        when "00011010" => datar <= "0010010100101000";datai <= "1000010110000100"; --208
        when "00011011" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "00011100" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "00011101" => datar <= "0001001011001000";datai <= "1000000101100100"; --232
        when "00011110" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "00011111" => datar <= "0000011001001000";datai <= "1000000000101000"; --248
        when "00100000" => datar <= "0000000000000000";datai <= "1000000000000001"; --256
        when "00100001" => datar <= "1111100110111000";datai <= "1000000000101000"; --264
        when "00100010" => datar <= "1111001101110100";datai <= "1000000010011111"; --272
        when "00100011" => datar <= "1110110100111000";datai <= "1000000101100100"; --280
        when "00100100" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "00100101" => datar <= "1110000011100110";datai <= "1000001111010111"; --296
        when "00100110" => datar <= "1101101011011000";datai <= "1000010110000100"; --304
        when "00100111" => datar <= "1101010011100001";datai <= "1000011101111100"; --312
        when "00101000" => datar <= "1100111100000101";datai <= "1000100110111111"; --320
        when "00101001" => datar <= "1100100101000110";datai <= "1000110001001011"; --328
        when "00101010" => datar <= "1100001110101010";datai <= "1000111100011110"; --336
        when "00101011" => datar <= "1011111000110010";datai <= "1001001000110111"; --344
        when "00101100" => datar <= "1011100011100100";datai <= "1001010110010011"; --352
        when "00101101" => datar <= "1011001111000001";datai <= "1001100100110001"; --360
        when "00101110" => datar <= "1010111011001101";datai <= "1001110100001111"; --368
        when "00101111" => datar <= "1010101000001011";datai <= "1010000100101001"; --376
        when "00110000" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "00110001" => datar <= "1010000100101001";datai <= "1010101000001011"; --392
        when "00110010" => datar <= "1001110100001111";datai <= "1010111011001101"; --400
        when "00110011" => datar <= "1001100100110001";datai <= "1011001111000001"; --408
        when "00110100" => datar <= "1001010110010011";datai <= "1011100011100100"; --416
        when "00110101" => datar <= "1001001000110111";datai <= "1011111000110010"; --424
        when "00110110" => datar <= "1000111100011110";datai <= "1100001110101010"; --432
        when "00110111" => datar <= "1000110001001011";datai <= "1100100101000110"; --440
        when "00111000" => datar <= "1000100110111111";datai <= "1100111100000101"; --448
        when "00111001" => datar <= "1000011101111100";datai <= "1101010011100001"; --456
        when "00111010" => datar <= "1000010110000100";datai <= "1101101011011000"; --464
        when "00111011" => datar <= "1000001111010111";datai <= "1110000011100110"; --472
        when "00111100" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "00111101" => datar <= "1000000101100100";datai <= "1110110100111000"; --488
        when "00111110" => datar <= "1000000010011111";datai <= "1111001101110100"; --496
        when "00111111" => datar <= "1000000000101000";datai <= "1111100110111000"; --504
        when "01000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "01000001" => datar <= "0111111111110101";datai <= "1111110011011100"; --4
        when "01000010" => datar <= "0111111111011000";datai <= "1111100110111000"; --8
        when "01000011" => datar <= "0111111110100110";datai <= "1111011010010110"; --12
        when "01000100" => datar <= "0111111101100001";datai <= "1111001101110100"; --16
        when "01000101" => datar <= "0111111100001001";datai <= "1111000001010101"; --20
        when "01000110" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "01000111" => datar <= "0111111000011101";datai <= "1110101000011110"; --28
        when "01001000" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "01001001" => datar <= "0111110011100011";datai <= "1110001111110101"; --36
        when "01001010" => datar <= "0111110000101001";datai <= "1110000011100110"; --40
        when "01001011" => datar <= "0111101101011100";datai <= "1101110111011101"; --44
        when "01001100" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "01001101" => datar <= "0111100110001001";datai <= "1101011111011010"; --52
        when "01001110" => datar <= "0111100010000100";datai <= "1101010011100001"; --56
        when "01001111" => datar <= "0111011101101011";datai <= "1101000111101111"; --60
        when "01010000" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "01010001" => datar <= "0111010100000100";datai <= "1100110000100001"; --68
        when "01010010" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "01010011" => datar <= "0111001001010100";datai <= "1100011001110100"; --76
        when "01010100" => datar <= "0111000011100010";datai <= "1100001110101010"; --80
        when "01010101" => datar <= "0110111101011110";datai <= "1100000011101001"; --84
        when "01010110" => datar <= "0110110111001001";datai <= "1011111000110010"; --88
        when "01010111" => datar <= "0110110000100011";datai <= "1011101110000110"; --92
        when "01011000" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "01011001" => datar <= "0110100010100110";datai <= "1011011001001100"; --100
        when "01011010" => datar <= "0110011011001111";datai <= "1011001111000001"; --104
        when "01011011" => datar <= "0110010011101000";datai <= "1011000101000001"; --108
        when "01011100" => datar <= "0110001011110001";datai <= "1010111011001101"; --112
        when "01011101" => datar <= "0110000011101011";datai <= "1010110001100101"; --116
        when "01011110" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "01011111" => datar <= "0101110010110011";datai <= "1010011110111110"; --124
        when "01100000" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "01100001" => datar <= "0101100001000010";datai <= "1010001101001101"; --132
        when "01100010" => datar <= "0101010111110101";datai <= "1010000100101001"; --136
        when "01100011" => datar <= "0101001110011011";datai <= "1001111100010101"; --140
        when "01100100" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "01100101" => datar <= "0100111010111111";datai <= "1001101100011000"; --148
        when "01100110" => datar <= "0100110000111111";datai <= "1001100100110001"; --152
        when "01100111" => datar <= "0100100110110100";datai <= "1001011101011010"; --156
        when "01101000" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "01101001" => datar <= "0100010001111010";datai <= "1001001111011101"; --164
        when "01101010" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "01101011" => datar <= "0011111100010111";datai <= "1001000010100010"; --172
        when "01101100" => datar <= "0011110001010110";datai <= "1000111100011110"; --176
        when "01101101" => datar <= "0011100110001100";datai <= "1000110110101100"; --180
        when "01101110" => datar <= "0011011010111010";datai <= "1000110001001011"; --184
        when "01101111" => datar <= "0011001111011111";datai <= "1000101011111100"; --188
        when "01110000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "01110001" => datar <= "0010111000010001";datai <= "1000100010010101"; --196
        when "01110010" => datar <= "0010101100011111";datai <= "1000011101111100"; --200
        when "01110011" => datar <= "0010100000100110";datai <= "1000011001110111"; --204
        when "01110100" => datar <= "0010010100101000";datai <= "1000010110000100"; --208
        when "01110101" => datar <= "0010001000100011";datai <= "1000010010100100"; --212
        when "01110110" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "01110111" => datar <= "0001110000001011";datai <= "1000001100011101"; --220
        when "01111000" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "01111001" => datar <= "0001010111100010";datai <= "1000000111100011"; --228
        when "01111010" => datar <= "0001001011001000";datai <= "1000000101100100"; --232
        when "01111011" => datar <= "0000111110101011";datai <= "1000000011110111"; --236
        when "01111100" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "01111101" => datar <= "0000100101101010";datai <= "1000000001011010"; --244
        when "01111110" => datar <= "0000011001001000";datai <= "1000000000101000"; --248
        when "01111111" => datar <= "0000001100100100";datai <= "1000000000001011"; --252
        when "10000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "10000001" => datar <= "0111111110100110";datai <= "1111011010010110"; --12
        when "10000010" => datar <= "0111111010011100";datai <= "1110110100111000"; --24
        when "10000011" => datar <= "0111110011100011";datai <= "1110001111110101"; --36
        when "10000100" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "10000101" => datar <= "0111011101101011";datai <= "1101000111101111"; --60
        when "10000110" => datar <= "0111001110110101";datai <= "1100100101000110"; --72
        when "10000111" => datar <= "0110111101011110";datai <= "1100000011101001"; --84
        when "10001000" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "10001001" => datar <= "0110010011101000";datai <= "1011000101000001"; --108
        when "10001010" => datar <= "0101111011010111";datai <= "1010101000001011"; --120
        when "10001011" => datar <= "0101100001000010";datai <= "1010001101001101"; --132
        when "10001100" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "10001101" => datar <= "0100100110110100";datai <= "1001011101011010"; --156
        when "10001110" => datar <= "0100000111001110";datai <= "1001001000110111"; --168
        when "10001111" => datar <= "0011100110001100";datai <= "1000110110101100"; --180
        when "10010000" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "10010001" => datar <= "0010100000100110";datai <= "1000011001110111"; --204
        when "10010010" => datar <= "0001111100011010";datai <= "1000001111010111"; --216
        when "10010011" => datar <= "0001010111100010";datai <= "1000000111100011"; --228
        when "10010100" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "10010101" => datar <= "0000001100100100";datai <= "1000000000001011"; --252
        when "10010110" => datar <= "1111100110111000";datai <= "1000000000101000"; --264
        when "10010111" => datar <= "1111000001010101";datai <= "1000000011110111"; --276
        when "10011000" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "10011001" => datar <= "1101110111011101";datai <= "1000010010100100"; --300
        when "10011010" => datar <= "1101010011100001";datai <= "1000011101111100"; --312
        when "10011011" => datar <= "1100110000100001";datai <= "1000101011111100"; --324
        when "10011100" => datar <= "1100001110101010";datai <= "1000111100011110"; --336
        when "10011101" => datar <= "1011101110000110";datai <= "1001001111011101"; --348
        when "10011110" => datar <= "1011001111000001";datai <= "1001100100110001"; --360
        when "10011111" => datar <= "1010110001100101";datai <= "1001111100010101"; --372
        when "10100000" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "10100001" => datar <= "1001111100010101";datai <= "1010110001100101"; --396
        when "10100010" => datar <= "1001100100110001";datai <= "1011001111000001"; --408
        when "10100011" => datar <= "1001001111011101";datai <= "1011101110000110"; --420
        when "10100100" => datar <= "1000111100011110";datai <= "1100001110101010"; --432
        when "10100101" => datar <= "1000101011111100";datai <= "1100110000100001"; --444
        when "10100110" => datar <= "1000011101111100";datai <= "1101010011100001"; --456
        when "10100111" => datar <= "1000010010100100";datai <= "1101110111011101"; --468
        when "10101000" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "10101001" => datar <= "1000000011110111";datai <= "1111000001010101"; --492
        when "10101010" => datar <= "1000000000101000";datai <= "1111100110111000"; --504
        when "10101011" => datar <= "1000000000001011";datai <= "0000001100100100"; --516
        when "10101100" => datar <= "1000000010011111";datai <= "0000110010001100"; --528
        when "10101101" => datar <= "1000000111100011";datai <= "0001010111100010"; --540
        when "10101110" => datar <= "1000001111010111";datai <= "0001111100011010"; --552
        when "10101111" => datar <= "1000011001110111";datai <= "0010100000100110"; --564
        when "10110000" => datar <= "1000100110111111";datai <= "0011000011111011"; --576
        when "10110001" => datar <= "1000110110101100";datai <= "0011100110001100"; --588
        when "10110010" => datar <= "1001001000110111";datai <= "0100000111001110"; --600
        when "10110011" => datar <= "1001011101011010";datai <= "0100100110110100"; --612
        when "10110100" => datar <= "1001110100001111";datai <= "0101000100110011"; --624
        when "10110101" => datar <= "1010001101001101";datai <= "0101100001000010"; --636
        when "10110110" => datar <= "1010101000001011";datai <= "0101111011010111"; --648
        when "10110111" => datar <= "1011000101000001";datai <= "0110010011101000"; --660
        when "10111000" => datar <= "1011100011100100";datai <= "0110101001101101"; --672
        when "10111001" => datar <= "1100000011101001";datai <= "0110111101011110"; --684
        when "10111010" => datar <= "1100100101000110";datai <= "0111001110110101"; --696
        when "10111011" => datar <= "1101000111101111";datai <= "0111011101101011"; --708
        when "10111100" => datar <= "1101101011011000";datai <= "0111101001111100"; --720
        when "10111101" => datar <= "1110001111110101";datai <= "0111110011100011"; --732
        when "10111110" => datar <= "1110110100111000";datai <= "0111111010011100"; --744
        when "10111111" => datar <= "1111011010010110";datai <= "0111111110100110"; --756
           when "11000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11000111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11001111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11010111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11011111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11100111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11101111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "11111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when others => for i in data_width-1 downto 0 loop
            datar(i)<='0';datai(i)<='0';end loop;
    end case;

    end if;

end process;
END behavior;
