/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`timescale 1ns / 1ps
`define P 20

`define M     503         // M is the degree of the irreducible polynomial
`define WIDTH (2*`M-1)    // width for a GF(3^M) element
`define WIDTH_D0 (1008-1)

module test_pe;

	// Inputs
	reg clk;
	reg reset;
	reg [10:0] ctrl;
	reg [`WIDTH_D0:0] d0;
	reg [`WIDTH:0] d1;
	reg [`WIDTH:0] d2;
    reg [`WIDTH:0] wish;

	// Outputs
	wire [`WIDTH:0] out;

	// Instantiate the Unit Under Test (UUT)
	PE uut (
		.clk(clk), 
		.reset(reset), 
		.ctrl(ctrl), 
		.d0(d0), 
		.d1(d1), 
        .d2(d2),
		.out(out)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		ctrl = 0;
		d0 = 0;
		d1 = 0;
        d2 = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
        // test mult
        d0 = 1006'h1119248464094a51549514585519508512555548915458194454a95a5a6550224816556284a5412965419544014a511556aa55955144aa5699655618601a19691a6691682455451456154a4585906a8615595595560656a15511545a9029959510158140619554a45a96a199aa69010216541569025125a4999591561495;
        d1 = 1006'h1a55960985561659551851556895049209954912568a591559455151a6a96614a415025691809658645a12a415a665241565a565896195925a558154045551590a9610255981a119295065a605955445a165985126506828941554156694564a29585611655965010115198aa64986559214641456656425290954464964;
        d2 = d1;
        wish = 1006'h296690698528561902a89185a6682428590645221996249986180602212996548298118549a161545666651980291a9806a99a9911a2044444908214800aaa04402a2209496440aa11991aa5949a0152899416598196510996a5a50629996aa68a4a9150058552196045aa42209094906684805604282410248094120a61;
        
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b00000_111111; #(168*`P);
        check;
        
        // test cubic
        d0 = {6'b10101, 1002'd0};
        d1 = 1006'h1119248464094a51549514585519508512555548915458194454a95a5a6550224816556284a5412965419544014a511556aa55955144aa5699655618601a19691a6691682455451456154a4585906a8615595595560656a15511545a9029959510158140619554a45a96a199aa69010216541569025125a4999591561495;
        d2 = d1;
        wish = 1006'h25025a210a560a450298548062454110aa9458192245809a45964889a65a258440598a41411492199a15615080a4159911826049059a691598688804a991996924864959490519956855484104849a08904919aa59886a56859269504516a0aa604a49215a25a129458a6944aa5495981061589105441842001a50899565;
        
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=1; #(`P);
        check;
        
        // test add
        d0 = {6'b000101, 1002'd0};
        d1 = 1006'h1119248464094a51549514585519508512555548915458194454a95a5a6550224816556284a5412965419544014a511556aa55955144aa5699655618601a19691a6691682455451456154a4585906a8615595595560656a15511545a9029959510158140619554a45a96a199aa69010216541569025125a4999591561495;
        d2 = 1006'h1a55960985561659551851556895049209954912568a591559455151a6a96614a415025691809658645a12a415a665241565a565896195925a558154045551590a9610255981a119295065a605955445a165985126506828941554156694564a29585611655965010115198aa64986559214641456656425290954464964;
        wish = 1006'h28628a81295051aaa9a165a181a25454182a925a2412a52291990aa80112860620285485556514459998a4281621860968100a0a1aa54025248a146064606a861509a151411626214065a0288a65820886822126495682992926a8600681281009611451962289a558a88a5451a68454a568494155865999869225995109;
        
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b10001; #(`P);
        check;

        // test sub
        d0 = {6'b001001, 1002'd0};
        d1 = 1006'h1119248464094a51549514585519508512555548915458194454a95a5a6550224816556284a5412965419544014a511556aa55955144aa5699655618601a19691a6691682455451456154a4585906a8615595595560656a15511545a9029959510158140619554a45a96a199aa69010216541569025125a4999591561495;
        d2 = 1006'h1a55960985561659551851556895049209954912568a591559455151a6a96614a415025691809658645a12a415a665241565a565896195925a558154045551590a9610255981a119295065a605955445a165985126506828941554156694564a29585611655965010115198aa64986559214641456656425290954464964;
        wish = 1006'h0684518aa2a664040289860629445826158018694a9902042a125809a488291a940156182625aa9101268690289428214145a060941615844210958468858810109081469a94940a69851592800a16416424894460a62a85810800456955425a26896a62084822a65981941204204aa94440a155a8288182a09849109a61;
        
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b10001; #(`P);
        check;

        $display("Good!");
        $finish;
	end

    initial #100 forever #(`P/2) clk = ~clk;

    task check;
        begin
          if (out !== wish)
            begin $display("E %h %h", out, wish); $finish; end
        end
    endtask
endmodule

