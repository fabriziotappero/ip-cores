----------------------------------------------------------------------
----                                                              ----
----  delayer_synth.vhd                                           ----
----                                                              ----
----  This file is part of the turbo decoder IP core project      ----
----  http://www.opencores.org/projects/turbocodes/               ----
----                                                              ----
----  Author(s):                                                  ----
----      - David Brochart(dbrochart@opencores.org)               ----
----                                                              ----
----  All additional information is available in the README.txt   ----
----  file.                                                       ----
----                                                              ----
----------------------------------------------------------------------
----                                                              ----
---- Copyright (C) 2005 Authors                                   ----
----                                                              ----
---- This source file may be used and distributed without         ----
---- restriction provided that this copyright statement is not    ----
---- removed from the file and that any derivative work contains  ----
---- the original copyright notice and the associated disclaimer. ----
----                                                              ----
---- This source file is free software; you can redistribute it   ----
---- and/or modify it under the terms of the GNU Lesser General   ----
---- Public License as published by the Free Software Foundation; ----
---- either version 2.1 of the License, or (at your option) any   ----
---- later version.                                               ----
----                                                              ----
---- This source is distributed in the hope that it will be       ----
---- useful, but WITHOUT ANY WARRANTY; without even the implied   ----
---- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ----
---- PURPOSE. See the GNU Lesser General Public License for more  ----
---- details.                                                     ----
----                                                              ----
---- You should have received a copy of the GNU Lesser General    ----
---- Public License along with this source; if not, download it   ----
---- from http://www.opencores.org/lgpl.shtml                     ----
----                                                              ----
----------------------------------------------------------------------



architecture synth of delayer is
    type ARRAYdelay is array (0 to delay - 1) of std_logic_vector(d'length - 1 downto 0);
    signal r    : ARRAYdelay;
begin
    process (clk, rst)
    begin
        if rst = '0' then
            q <= std_logic_vector(conv_unsigned(0, d'length));
            for i in 0 to delay - 1 loop
                r(i) <= (others => '0');
            end loop;
        elsif clk = '1' and clk'event then
            r(0)    <= d;
            q       <= r(delay - 1);
            for i in 0 to delay - 2 loop
                r(i + 1) <= r(i);
            end loop;
        end if;
    end process;
end;
