library verilog;
use verilog.vl_types.all;
entity testcase_1 is
end testcase_1;
