
///
/// created by oc8051 rom maker
/// author: Simon Teran (simont@opencores.org)
///
/// source file: D:\verilog\oc8051\test\testall.hex
/// date: 17.6.02
/// time: 10:53:03
///

module oc8051_rom (rst, clk, addr, ea_int, data1, data2, data3);

parameter INT_ROM_WID= 12;

input rst, clk;
input [15:0] addr;
output ea_int;
output [7:0] data1, data2, data3;
reg [7:0] data1, data2, data3;
reg [7:0] buff [65535:0];
integer i;

wire ea;

assign ea = | addr[15:INT_ROM_WID];
assign ea_int = ! ea;

initial
begin
    for (i=0; i<65536; i=i+1)
      buff [i] = 8'h00;
#2

    buff [16'h00_00] = 8'h78;
    buff [16'h00_01] = 8'h80;
    buff [16'h00_02] = 8'h18;
    buff [16'h00_03] = 8'h76;
    buff [16'h00_04] = 8'h00;
    buff [16'h00_05] = 8'hE8;
    buff [16'h00_06] = 8'h70;
    buff [16'h00_07] = 8'hFA;
    buff [16'h00_08] = 8'h75;
    buff [16'h00_09] = 8'hD0;
    buff [16'h00_0a] = 8'h00;
    buff [16'h00_0b] = 8'h74;
    buff [16'h00_0c] = 8'h0A;
    buff [16'h00_0d] = 8'h78;
    buff [16'h00_0e] = 8'h0A;
    buff [16'h00_0f] = 8'h28;
    buff [16'h00_10] = 8'h94;
    buff [16'h00_11] = 8'h14;
    buff [16'h00_12] = 8'h60;
    buff [16'h00_13] = 8'h06;
    buff [16'h00_14] = 8'h75;
    buff [16'h00_15] = 8'h90;
    buff [16'h00_16] = 8'h02;
    buff [16'h00_17] = 8'h02;
    buff [16'h00_18] = 8'h0A;
    buff [16'h00_19] = 8'hF0;
    buff [16'h00_1a] = 8'h78;
    buff [16'h00_1b] = 8'h80;
    buff [16'h00_1c] = 8'h18;
    buff [16'h00_1d] = 8'h76;
    buff [16'h00_1e] = 8'h00;
    buff [16'h00_1f] = 8'hE8;
    buff [16'h00_20] = 8'h70;
    buff [16'h00_21] = 8'hFA;
    buff [16'h00_22] = 8'h75;
    buff [16'h00_23] = 8'hD0;
    buff [16'h00_24] = 8'h00;
    buff [16'h00_25] = 8'h74;
    buff [16'h00_26] = 8'h0A;
    buff [16'h00_27] = 8'h75;
    buff [16'h00_28] = 8'h64;
    buff [16'h00_29] = 8'h0A;
    buff [16'h00_2a] = 8'h25;
    buff [16'h00_2b] = 8'h64;
    buff [16'h00_2c] = 8'h94;
    buff [16'h00_2d] = 8'h14;
    buff [16'h00_2e] = 8'h60;
    buff [16'h00_2f] = 8'h06;
    buff [16'h00_30] = 8'h75;
    buff [16'h00_31] = 8'h90;
    buff [16'h00_32] = 8'h03;
    buff [16'h00_33] = 8'h02;
    buff [16'h00_34] = 8'h0A;
    buff [16'h00_35] = 8'hF0;
    buff [16'h00_36] = 8'h78;
    buff [16'h00_37] = 8'h80;
    buff [16'h00_38] = 8'h18;
    buff [16'h00_39] = 8'h76;
    buff [16'h00_3a] = 8'h00;
    buff [16'h00_3b] = 8'hE8;
    buff [16'h00_3c] = 8'h70;
    buff [16'h00_3d] = 8'hFA;
    buff [16'h00_3e] = 8'h75;
    buff [16'h00_3f] = 8'hD0;
    buff [16'h00_40] = 8'h00;
    buff [16'h00_41] = 8'h74;
    buff [16'h00_42] = 8'h0A;
    buff [16'h00_43] = 8'h78;
    buff [16'h00_44] = 8'h64;
    buff [16'h00_45] = 8'h75;
    buff [16'h00_46] = 8'h64;
    buff [16'h00_47] = 8'h0A;
    buff [16'h00_48] = 8'h26;
    buff [16'h00_49] = 8'h94;
    buff [16'h00_4a] = 8'h14;
    buff [16'h00_4b] = 8'h60;
    buff [16'h00_4c] = 8'h06;
    buff [16'h00_4d] = 8'h75;
    buff [16'h00_4e] = 8'h90;
    buff [16'h00_4f] = 8'h04;
    buff [16'h00_50] = 8'h02;
    buff [16'h00_51] = 8'h0A;
    buff [16'h00_52] = 8'hF0;
    buff [16'h00_53] = 8'h78;
    buff [16'h00_54] = 8'h80;
    buff [16'h00_55] = 8'h18;
    buff [16'h00_56] = 8'h76;
    buff [16'h00_57] = 8'h00;
    buff [16'h00_58] = 8'hE8;
    buff [16'h00_59] = 8'h70;
    buff [16'h00_5a] = 8'hFA;
    buff [16'h00_5b] = 8'h75;
    buff [16'h00_5c] = 8'hD0;
    buff [16'h00_5d] = 8'h00;
    buff [16'h00_5e] = 8'h74;
    buff [16'h00_5f] = 8'h0A;
    buff [16'h00_60] = 8'h24;
    buff [16'h00_61] = 8'h05;
    buff [16'h00_62] = 8'h94;
    buff [16'h00_63] = 8'h0F;
    buff [16'h00_64] = 8'h60;
    buff [16'h00_65] = 8'h06;
    buff [16'h00_66] = 8'h75;
    buff [16'h00_67] = 8'h90;
    buff [16'h00_68] = 8'h05;
    buff [16'h00_69] = 8'h02;
    buff [16'h00_6a] = 8'h0A;
    buff [16'h00_6b] = 8'hF0;
    buff [16'h00_6c] = 8'h78;
    buff [16'h00_6d] = 8'h80;
    buff [16'h00_6e] = 8'h18;
    buff [16'h00_6f] = 8'h76;
    buff [16'h00_70] = 8'h00;
    buff [16'h00_71] = 8'hE8;
    buff [16'h00_72] = 8'h70;
    buff [16'h00_73] = 8'hFA;
    buff [16'h00_74] = 8'h75;
    buff [16'h00_75] = 8'hD0;
    buff [16'h00_76] = 8'h00;
    buff [16'h00_77] = 8'h74;
    buff [16'h00_78] = 8'h0A;
    buff [16'h00_79] = 8'h78;
    buff [16'h00_7a] = 8'h0A;
    buff [16'h00_7b] = 8'hB3;
    buff [16'h00_7c] = 8'h38;
    buff [16'h00_7d] = 8'h94;
    buff [16'h00_7e] = 8'h15;
    buff [16'h00_7f] = 8'h60;
    buff [16'h00_80] = 8'h06;
    buff [16'h00_81] = 8'h75;
    buff [16'h00_82] = 8'h90;
    buff [16'h00_83] = 8'h06;
    buff [16'h00_84] = 8'h02;
    buff [16'h00_85] = 8'h0A;
    buff [16'h00_86] = 8'hF0;
    buff [16'h00_87] = 8'h78;
    buff [16'h00_88] = 8'h80;
    buff [16'h00_89] = 8'h18;
    buff [16'h00_8a] = 8'h76;
    buff [16'h00_8b] = 8'h00;
    buff [16'h00_8c] = 8'hE8;
    buff [16'h00_8d] = 8'h70;
    buff [16'h00_8e] = 8'hFA;
    buff [16'h00_8f] = 8'h75;
    buff [16'h00_90] = 8'hD0;
    buff [16'h00_91] = 8'h00;
    buff [16'h00_92] = 8'h74;
    buff [16'h00_93] = 8'h0A;
    buff [16'h00_94] = 8'h75;
    buff [16'h00_95] = 8'h64;
    buff [16'h00_96] = 8'h0A;
    buff [16'h00_97] = 8'hB3;
    buff [16'h00_98] = 8'h35;
    buff [16'h00_99] = 8'h64;
    buff [16'h00_9a] = 8'h94;
    buff [16'h00_9b] = 8'h15;
    buff [16'h00_9c] = 8'h60;
    buff [16'h00_9d] = 8'h06;
    buff [16'h00_9e] = 8'h75;
    buff [16'h00_9f] = 8'h90;
    buff [16'h00_a0] = 8'h07;
    buff [16'h00_a1] = 8'h02;
    buff [16'h00_a2] = 8'h0A;
    buff [16'h00_a3] = 8'hF0;
    buff [16'h00_a4] = 8'h78;
    buff [16'h00_a5] = 8'h80;
    buff [16'h00_a6] = 8'h18;
    buff [16'h00_a7] = 8'h76;
    buff [16'h00_a8] = 8'h00;
    buff [16'h00_a9] = 8'hE8;
    buff [16'h00_aa] = 8'h70;
    buff [16'h00_ab] = 8'hFA;
    buff [16'h00_ac] = 8'h75;
    buff [16'h00_ad] = 8'hD0;
    buff [16'h00_ae] = 8'h00;
    buff [16'h00_af] = 8'h74;
    buff [16'h00_b0] = 8'h0A;
    buff [16'h00_b1] = 8'h78;
    buff [16'h00_b2] = 8'h64;
    buff [16'h00_b3] = 8'h75;
    buff [16'h00_b4] = 8'h64;
    buff [16'h00_b5] = 8'h0A;
    buff [16'h00_b6] = 8'hB3;
    buff [16'h00_b7] = 8'h36;
    buff [16'h00_b8] = 8'h94;
    buff [16'h00_b9] = 8'h15;
    buff [16'h00_ba] = 8'h60;
    buff [16'h00_bb] = 8'h06;
    buff [16'h00_bc] = 8'h75;
    buff [16'h00_bd] = 8'h90;
    buff [16'h00_be] = 8'h08;
    buff [16'h00_bf] = 8'h02;
    buff [16'h00_c0] = 8'h0A;
    buff [16'h00_c1] = 8'hF0;
    buff [16'h00_c2] = 8'h78;
    buff [16'h00_c3] = 8'h80;
    buff [16'h00_c4] = 8'h18;
    buff [16'h00_c5] = 8'h76;
    buff [16'h00_c6] = 8'h00;
    buff [16'h00_c7] = 8'hE8;
    buff [16'h00_c8] = 8'h70;
    buff [16'h00_c9] = 8'hFA;
    buff [16'h00_ca] = 8'h75;
    buff [16'h00_cb] = 8'hD0;
    buff [16'h00_cc] = 8'h00;
    buff [16'h00_cd] = 8'h74;
    buff [16'h00_ce] = 8'h0A;
    buff [16'h00_cf] = 8'hB3;
    buff [16'h00_d0] = 8'h34;
    buff [16'h00_d1] = 8'h05;
    buff [16'h00_d2] = 8'h94;
    buff [16'h00_d3] = 8'h10;
    buff [16'h00_d4] = 8'h60;
    buff [16'h00_d5] = 8'h06;
    buff [16'h00_d6] = 8'h75;
    buff [16'h00_d7] = 8'h90;
    buff [16'h00_d8] = 8'h09;
    buff [16'h00_d9] = 8'h02;
    buff [16'h00_da] = 8'h0A;
    buff [16'h00_db] = 8'hF0;
    buff [16'h00_dc] = 8'h78;
    buff [16'h00_dd] = 8'h80;
    buff [16'h00_de] = 8'h18;
    buff [16'h00_df] = 8'h76;
    buff [16'h00_e0] = 8'h00;
    buff [16'h00_e1] = 8'hE8;
    buff [16'h00_e2] = 8'h70;
    buff [16'h00_e3] = 8'hFA;
    buff [16'h00_e4] = 8'h75;
    buff [16'h00_e5] = 8'hD0;
    buff [16'h00_e6] = 8'h00;
    buff [16'h00_e7] = 8'h01;
    buff [16'h00_e8] = 8'hEF;
    buff [16'h00_e9] = 8'h75;
    buff [16'h00_ea] = 8'h90;
    buff [16'h00_eb] = 8'h0A;
    buff [16'h00_ec] = 8'h02;
    buff [16'h00_ed] = 8'h0A;
    buff [16'h00_ee] = 8'hF0;
    buff [16'h00_ef] = 8'h78;
    buff [16'h00_f0] = 8'h80;
    buff [16'h00_f1] = 8'h18;
    buff [16'h00_f2] = 8'h76;
    buff [16'h00_f3] = 8'h00;
    buff [16'h00_f4] = 8'hE8;
    buff [16'h00_f5] = 8'h70;
    buff [16'h00_f6] = 8'hFA;
    buff [16'h00_f7] = 8'h75;
    buff [16'h00_f8] = 8'hD0;
    buff [16'h00_f9] = 8'h00;
    buff [16'h00_fa] = 8'h78;
    buff [16'h00_fb] = 8'hFF;
    buff [16'h00_fc] = 8'h74;
    buff [16'h00_fd] = 8'hAA;
    buff [16'h00_fe] = 8'h58;
    buff [16'h00_ff] = 8'h94;
    buff [16'h01_00] = 8'hAA;
    buff [16'h01_01] = 8'h60;
    buff [16'h01_02] = 8'h06;
    buff [16'h01_03] = 8'h75;
    buff [16'h01_04] = 8'h90;
    buff [16'h01_05] = 8'h0B;
    buff [16'h01_06] = 8'h02;
    buff [16'h01_07] = 8'h0A;
    buff [16'h01_08] = 8'hF0;
    buff [16'h01_09] = 8'h78;
    buff [16'h01_0a] = 8'h80;
    buff [16'h01_0b] = 8'h18;
    buff [16'h01_0c] = 8'h76;
    buff [16'h01_0d] = 8'h00;
    buff [16'h01_0e] = 8'hE8;
    buff [16'h01_0f] = 8'h70;
    buff [16'h01_10] = 8'hFA;
    buff [16'h01_11] = 8'h75;
    buff [16'h01_12] = 8'hD0;
    buff [16'h01_13] = 8'h00;
    buff [16'h01_14] = 8'h75;
    buff [16'h01_15] = 8'h7F;
    buff [16'h01_16] = 8'h00;
    buff [16'h01_17] = 8'h74;
    buff [16'h01_18] = 8'hFF;
    buff [16'h01_19] = 8'h55;
    buff [16'h01_1a] = 8'h7F;
    buff [16'h01_1b] = 8'h60;
    buff [16'h01_1c] = 8'h06;
    buff [16'h01_1d] = 8'h75;
    buff [16'h01_1e] = 8'h90;
    buff [16'h01_1f] = 8'h0C;
    buff [16'h01_20] = 8'h02;
    buff [16'h01_21] = 8'h0A;
    buff [16'h01_22] = 8'hF0;
    buff [16'h01_23] = 8'h78;
    buff [16'h01_24] = 8'h80;
    buff [16'h01_25] = 8'h18;
    buff [16'h01_26] = 8'h76;
    buff [16'h01_27] = 8'h00;
    buff [16'h01_28] = 8'hE8;
    buff [16'h01_29] = 8'h70;
    buff [16'h01_2a] = 8'hFA;
    buff [16'h01_2b] = 8'h75;
    buff [16'h01_2c] = 8'hD0;
    buff [16'h01_2d] = 8'h00;
    buff [16'h01_2e] = 8'h78;
    buff [16'h01_2f] = 8'h7F;
    buff [16'h01_30] = 8'h75;
    buff [16'h01_31] = 8'h7F;
    buff [16'h01_32] = 8'h01;
    buff [16'h01_33] = 8'h74;
    buff [16'h01_34] = 8'hFE;
    buff [16'h01_35] = 8'h56;
    buff [16'h01_36] = 8'h60;
    buff [16'h01_37] = 8'h06;
    buff [16'h01_38] = 8'h75;
    buff [16'h01_39] = 8'h90;
    buff [16'h01_3a] = 8'h0D;
    buff [16'h01_3b] = 8'h02;
    buff [16'h01_3c] = 8'h0A;
    buff [16'h01_3d] = 8'hF0;
    buff [16'h01_3e] = 8'h78;
    buff [16'h01_3f] = 8'h80;
    buff [16'h01_40] = 8'h18;
    buff [16'h01_41] = 8'h76;
    buff [16'h01_42] = 8'h00;
    buff [16'h01_43] = 8'hE8;
    buff [16'h01_44] = 8'h70;
    buff [16'h01_45] = 8'hFA;
    buff [16'h01_46] = 8'h75;
    buff [16'h01_47] = 8'hD0;
    buff [16'h01_48] = 8'h00;
    buff [16'h01_49] = 8'h74;
    buff [16'h01_4a] = 8'hFF;
    buff [16'h01_4b] = 8'h54;
    buff [16'h01_4c] = 8'hFF;
    buff [16'h01_4d] = 8'h94;
    buff [16'h01_4e] = 8'hFF;
    buff [16'h01_4f] = 8'h60;
    buff [16'h01_50] = 8'h06;
    buff [16'h01_51] = 8'h75;
    buff [16'h01_52] = 8'h90;
    buff [16'h01_53] = 8'h0E;
    buff [16'h01_54] = 8'h02;
    buff [16'h01_55] = 8'h0A;
    buff [16'h01_56] = 8'hF0;
    buff [16'h01_57] = 8'h78;
    buff [16'h01_58] = 8'h80;
    buff [16'h01_59] = 8'h18;
    buff [16'h01_5a] = 8'h76;
    buff [16'h01_5b] = 8'h00;
    buff [16'h01_5c] = 8'hE8;
    buff [16'h01_5d] = 8'h70;
    buff [16'h01_5e] = 8'hFA;
    buff [16'h01_5f] = 8'h75;
    buff [16'h01_60] = 8'hD0;
    buff [16'h01_61] = 8'h00;
    buff [16'h01_62] = 8'h75;
    buff [16'h01_63] = 8'h32;
    buff [16'h01_64] = 8'hFF;
    buff [16'h01_65] = 8'h74;
    buff [16'h01_66] = 8'h00;
    buff [16'h01_67] = 8'h52;
    buff [16'h01_68] = 8'h32;
    buff [16'h01_69] = 8'hE5;
    buff [16'h01_6a] = 8'h32;
    buff [16'h01_6b] = 8'h60;
    buff [16'h01_6c] = 8'h06;
    buff [16'h01_6d] = 8'h75;
    buff [16'h01_6e] = 8'h90;
    buff [16'h01_6f] = 8'h0F;
    buff [16'h01_70] = 8'h02;
    buff [16'h01_71] = 8'h0A;
    buff [16'h01_72] = 8'hF0;
    buff [16'h01_73] = 8'h78;
    buff [16'h01_74] = 8'h80;
    buff [16'h01_75] = 8'h18;
    buff [16'h01_76] = 8'h76;
    buff [16'h01_77] = 8'h00;
    buff [16'h01_78] = 8'hE8;
    buff [16'h01_79] = 8'h70;
    buff [16'h01_7a] = 8'hFA;
    buff [16'h01_7b] = 8'h75;
    buff [16'h01_7c] = 8'hD0;
    buff [16'h01_7d] = 8'h00;
    buff [16'h01_7e] = 8'h75;
    buff [16'h01_7f] = 8'h19;
    buff [16'h01_80] = 8'h80;
    buff [16'h01_81] = 8'h53;
    buff [16'h01_82] = 8'h19;
    buff [16'h01_83] = 8'hFF;
    buff [16'h01_84] = 8'hE5;
    buff [16'h01_85] = 8'h19;
    buff [16'h01_86] = 8'h94;
    buff [16'h01_87] = 8'h80;
    buff [16'h01_88] = 8'h60;
    buff [16'h01_89] = 8'h06;
    buff [16'h01_8a] = 8'h75;
    buff [16'h01_8b] = 8'h90;
    buff [16'h01_8c] = 8'h10;
    buff [16'h01_8d] = 8'h02;
    buff [16'h01_8e] = 8'h0A;
    buff [16'h01_8f] = 8'hF0;
    buff [16'h01_90] = 8'h78;
    buff [16'h01_91] = 8'h80;
    buff [16'h01_92] = 8'h18;
    buff [16'h01_93] = 8'h76;
    buff [16'h01_94] = 8'h00;
    buff [16'h01_95] = 8'hE8;
    buff [16'h01_96] = 8'h70;
    buff [16'h01_97] = 8'hFA;
    buff [16'h01_98] = 8'h75;
    buff [16'h01_99] = 8'hD0;
    buff [16'h01_9a] = 8'h00;
    buff [16'h01_9b] = 8'h74;
    buff [16'h01_9c] = 8'h80;
    buff [16'h01_9d] = 8'hB3;
    buff [16'h01_9e] = 8'h82;
    buff [16'h01_9f] = 8'hE7;
    buff [16'h01_a0] = 8'h94;
    buff [16'h01_a1] = 8'h7F;
    buff [16'h01_a2] = 8'h60;
    buff [16'h01_a3] = 8'h06;
    buff [16'h01_a4] = 8'h75;
    buff [16'h01_a5] = 8'h90;
    buff [16'h01_a6] = 8'h11;
    buff [16'h01_a7] = 8'h02;
    buff [16'h01_a8] = 8'h0A;
    buff [16'h01_a9] = 8'hF0;
    buff [16'h01_aa] = 8'h78;
    buff [16'h01_ab] = 8'h80;
    buff [16'h01_ac] = 8'h18;
    buff [16'h01_ad] = 8'h76;
    buff [16'h01_ae] = 8'h00;
    buff [16'h01_af] = 8'hE8;
    buff [16'h01_b0] = 8'h70;
    buff [16'h01_b1] = 8'hFA;
    buff [16'h01_b2] = 8'h75;
    buff [16'h01_b3] = 8'hD0;
    buff [16'h01_b4] = 8'h00;
    buff [16'h01_b5] = 8'h74;
    buff [16'h01_b6] = 8'h80;
    buff [16'h01_b7] = 8'hB3;
    buff [16'h01_b8] = 8'hB0;
    buff [16'h01_b9] = 8'hE7;
    buff [16'h01_ba] = 8'h94;
    buff [16'h01_bb] = 8'h80;
    buff [16'h01_bc] = 8'h60;
    buff [16'h01_bd] = 8'h06;
    buff [16'h01_be] = 8'h75;
    buff [16'h01_bf] = 8'h90;
    buff [16'h01_c0] = 8'h12;
    buff [16'h01_c1] = 8'h02;
    buff [16'h01_c2] = 8'h0A;
    buff [16'h01_c3] = 8'hF0;
    buff [16'h01_c4] = 8'h78;
    buff [16'h01_c5] = 8'h80;
    buff [16'h01_c6] = 8'h18;
    buff [16'h01_c7] = 8'h76;
    buff [16'h01_c8] = 8'h00;
    buff [16'h01_c9] = 8'hE8;
    buff [16'h01_ca] = 8'h70;
    buff [16'h01_cb] = 8'hFA;
    buff [16'h01_cc] = 8'h75;
    buff [16'h01_cd] = 8'hD0;
    buff [16'h01_ce] = 8'h00;
    buff [16'h01_cf] = 8'h74;
    buff [16'h01_d0] = 8'h80;
    buff [16'h01_d1] = 8'h75;
    buff [16'h01_d2] = 8'h64;
    buff [16'h01_d3] = 8'h80;
    buff [16'h01_d4] = 8'hB5;
    buff [16'h01_d5] = 8'h64;
    buff [16'h01_d6] = 8'h05;
    buff [16'h01_d7] = 8'h74;
    buff [16'h01_d8] = 8'h7F;
    buff [16'h01_d9] = 8'hB5;
    buff [16'h01_da] = 8'h64;
    buff [16'h01_db] = 8'h06;
    buff [16'h01_dc] = 8'h75;
    buff [16'h01_dd] = 8'h90;
    buff [16'h01_de] = 8'h13;
    buff [16'h01_df] = 8'h02;
    buff [16'h01_e0] = 8'h0A;
    buff [16'h01_e1] = 8'hF0;
    buff [16'h01_e2] = 8'h40;
    buff [16'h01_e3] = 8'h06;
    buff [16'h01_e4] = 8'h75;
    buff [16'h01_e5] = 8'h90;
    buff [16'h01_e6] = 8'h13;
    buff [16'h01_e7] = 8'h02;
    buff [16'h01_e8] = 8'h0A;
    buff [16'h01_e9] = 8'hF0;
    buff [16'h01_ea] = 8'h78;
    buff [16'h01_eb] = 8'h80;
    buff [16'h01_ec] = 8'h18;
    buff [16'h01_ed] = 8'h76;
    buff [16'h01_ee] = 8'h00;
    buff [16'h01_ef] = 8'hE8;
    buff [16'h01_f0] = 8'h70;
    buff [16'h01_f1] = 8'hFA;
    buff [16'h01_f2] = 8'h75;
    buff [16'h01_f3] = 8'hD0;
    buff [16'h01_f4] = 8'h00;
    buff [16'h01_f5] = 8'h74;
    buff [16'h01_f6] = 8'h80;
    buff [16'h01_f7] = 8'hB4;
    buff [16'h01_f8] = 8'h80;
    buff [16'h01_f9] = 8'h05;
    buff [16'h01_fa] = 8'h74;
    buff [16'h01_fb] = 8'h7F;
    buff [16'h01_fc] = 8'hB4;
    buff [16'h01_fd] = 8'h80;
    buff [16'h01_fe] = 8'h06;
    buff [16'h01_ff] = 8'h75;
    buff [16'h02_00] = 8'h90;
    buff [16'h02_01] = 8'h14;
    buff [16'h02_02] = 8'h02;
    buff [16'h02_03] = 8'h0A;
    buff [16'h02_04] = 8'hF0;
    buff [16'h02_05] = 8'h40;
    buff [16'h02_06] = 8'h06;
    buff [16'h02_07] = 8'h75;
    buff [16'h02_08] = 8'h90;
    buff [16'h02_09] = 8'h14;
    buff [16'h02_0a] = 8'h02;
    buff [16'h02_0b] = 8'h0A;
    buff [16'h02_0c] = 8'hF0;
    buff [16'h02_0d] = 8'h78;
    buff [16'h02_0e] = 8'h80;
    buff [16'h02_0f] = 8'h18;
    buff [16'h02_10] = 8'h76;
    buff [16'h02_11] = 8'h00;
    buff [16'h02_12] = 8'hE8;
    buff [16'h02_13] = 8'h70;
    buff [16'h02_14] = 8'hFA;
    buff [16'h02_15] = 8'h75;
    buff [16'h02_16] = 8'hD0;
    buff [16'h02_17] = 8'h00;
    buff [16'h02_18] = 8'h79;
    buff [16'h02_19] = 8'h80;
    buff [16'h02_1a] = 8'hB9;
    buff [16'h02_1b] = 8'h80;
    buff [16'h02_1c] = 8'h05;
    buff [16'h02_1d] = 8'h79;
    buff [16'h02_1e] = 8'h7F;
    buff [16'h02_1f] = 8'hB9;
    buff [16'h02_20] = 8'h80;
    buff [16'h02_21] = 8'h06;
    buff [16'h02_22] = 8'h75;
    buff [16'h02_23] = 8'h90;
    buff [16'h02_24] = 8'h15;
    buff [16'h02_25] = 8'h02;
    buff [16'h02_26] = 8'h0A;
    buff [16'h02_27] = 8'hF0;
    buff [16'h02_28] = 8'h40;
    buff [16'h02_29] = 8'h06;
    buff [16'h02_2a] = 8'h75;
    buff [16'h02_2b] = 8'h90;
    buff [16'h02_2c] = 8'h15;
    buff [16'h02_2d] = 8'h02;
    buff [16'h02_2e] = 8'h0A;
    buff [16'h02_2f] = 8'hF0;
    buff [16'h02_30] = 8'h78;
    buff [16'h02_31] = 8'h80;
    buff [16'h02_32] = 8'h18;
    buff [16'h02_33] = 8'h76;
    buff [16'h02_34] = 8'h00;
    buff [16'h02_35] = 8'hE8;
    buff [16'h02_36] = 8'h70;
    buff [16'h02_37] = 8'hFA;
    buff [16'h02_38] = 8'h75;
    buff [16'h02_39] = 8'hD0;
    buff [16'h02_3a] = 8'h00;
    buff [16'h02_3b] = 8'h79;
    buff [16'h02_3c] = 8'h64;
    buff [16'h02_3d] = 8'h75;
    buff [16'h02_3e] = 8'h64;
    buff [16'h02_3f] = 8'h80;
    buff [16'h02_40] = 8'hB7;
    buff [16'h02_41] = 8'h80;
    buff [16'h02_42] = 8'h06;
    buff [16'h02_43] = 8'h75;
    buff [16'h02_44] = 8'h64;
    buff [16'h02_45] = 8'h7F;
    buff [16'h02_46] = 8'hB7;
    buff [16'h02_47] = 8'h80;
    buff [16'h02_48] = 8'h06;
    buff [16'h02_49] = 8'h75;
    buff [16'h02_4a] = 8'h90;
    buff [16'h02_4b] = 8'h16;
    buff [16'h02_4c] = 8'h02;
    buff [16'h02_4d] = 8'h0A;
    buff [16'h02_4e] = 8'hF0;
    buff [16'h02_4f] = 8'h40;
    buff [16'h02_50] = 8'h06;
    buff [16'h02_51] = 8'h75;
    buff [16'h02_52] = 8'h90;
    buff [16'h02_53] = 8'h16;
    buff [16'h02_54] = 8'h02;
    buff [16'h02_55] = 8'h0A;
    buff [16'h02_56] = 8'hF0;
    buff [16'h02_57] = 8'h78;
    buff [16'h02_58] = 8'h80;
    buff [16'h02_59] = 8'h18;
    buff [16'h02_5a] = 8'h76;
    buff [16'h02_5b] = 8'h00;
    buff [16'h02_5c] = 8'hE8;
    buff [16'h02_5d] = 8'h70;
    buff [16'h02_5e] = 8'hFA;
    buff [16'h02_5f] = 8'h75;
    buff [16'h02_60] = 8'hD0;
    buff [16'h02_61] = 8'h00;
    buff [16'h02_62] = 8'h74;
    buff [16'h02_63] = 8'h80;
    buff [16'h02_64] = 8'hE4;
    buff [16'h02_65] = 8'h60;
    buff [16'h02_66] = 8'h06;
    buff [16'h02_67] = 8'h75;
    buff [16'h02_68] = 8'h90;
    buff [16'h02_69] = 8'h17;
    buff [16'h02_6a] = 8'h02;
    buff [16'h02_6b] = 8'h0A;
    buff [16'h02_6c] = 8'hF0;
    buff [16'h02_6d] = 8'h78;
    buff [16'h02_6e] = 8'h80;
    buff [16'h02_6f] = 8'h18;
    buff [16'h02_70] = 8'h76;
    buff [16'h02_71] = 8'h00;
    buff [16'h02_72] = 8'hE8;
    buff [16'h02_73] = 8'h70;
    buff [16'h02_74] = 8'hFA;
    buff [16'h02_75] = 8'h75;
    buff [16'h02_76] = 8'hD0;
    buff [16'h02_77] = 8'h00;
    buff [16'h02_78] = 8'hB3;
    buff [16'h02_79] = 8'hC3;
    buff [16'h02_7a] = 8'h50;
    buff [16'h02_7b] = 8'h06;
    buff [16'h02_7c] = 8'h75;
    buff [16'h02_7d] = 8'h90;
    buff [16'h02_7e] = 8'h18;
    buff [16'h02_7f] = 8'h02;
    buff [16'h02_80] = 8'h0A;
    buff [16'h02_81] = 8'hF0;
    buff [16'h02_82] = 8'h78;
    buff [16'h02_83] = 8'h80;
    buff [16'h02_84] = 8'h18;
    buff [16'h02_85] = 8'h76;
    buff [16'h02_86] = 8'h00;
    buff [16'h02_87] = 8'hE8;
    buff [16'h02_88] = 8'h70;
    buff [16'h02_89] = 8'hFA;
    buff [16'h02_8a] = 8'h75;
    buff [16'h02_8b] = 8'hD0;
    buff [16'h02_8c] = 8'h00;
    buff [16'h02_8d] = 8'h74;
    buff [16'h02_8e] = 8'h40;
    buff [16'h02_8f] = 8'hC2;
    buff [16'h02_90] = 8'hE6;
    buff [16'h02_91] = 8'h60;
    buff [16'h02_92] = 8'h06;
    buff [16'h02_93] = 8'h75;
    buff [16'h02_94] = 8'h90;
    buff [16'h02_95] = 8'h19;
    buff [16'h02_96] = 8'h02;
    buff [16'h02_97] = 8'h0A;
    buff [16'h02_98] = 8'hF0;
    buff [16'h02_99] = 8'h78;
    buff [16'h02_9a] = 8'h80;
    buff [16'h02_9b] = 8'h18;
    buff [16'h02_9c] = 8'h76;
    buff [16'h02_9d] = 8'h00;
    buff [16'h02_9e] = 8'hE8;
    buff [16'h02_9f] = 8'h70;
    buff [16'h02_a0] = 8'hFA;
    buff [16'h02_a1] = 8'h75;
    buff [16'h02_a2] = 8'hD0;
    buff [16'h02_a3] = 8'h00;
    buff [16'h02_a4] = 8'h74;
    buff [16'h02_a5] = 8'hFF;
    buff [16'h02_a6] = 8'hF4;
    buff [16'h02_a7] = 8'h60;
    buff [16'h02_a8] = 8'h06;
    buff [16'h02_a9] = 8'h75;
    buff [16'h02_aa] = 8'h90;
    buff [16'h02_ab] = 8'h1A;
    buff [16'h02_ac] = 8'h02;
    buff [16'h02_ad] = 8'h0A;
    buff [16'h02_ae] = 8'hF0;
    buff [16'h02_af] = 8'h78;
    buff [16'h02_b0] = 8'h80;
    buff [16'h02_b1] = 8'h18;
    buff [16'h02_b2] = 8'h76;
    buff [16'h02_b3] = 8'h00;
    buff [16'h02_b4] = 8'hE8;
    buff [16'h02_b5] = 8'h70;
    buff [16'h02_b6] = 8'hFA;
    buff [16'h02_b7] = 8'h75;
    buff [16'h02_b8] = 8'hD0;
    buff [16'h02_b9] = 8'h00;
    buff [16'h02_ba] = 8'hB3;
    buff [16'h02_bb] = 8'h40;
    buff [16'h02_bc] = 8'h06;
    buff [16'h02_bd] = 8'h75;
    buff [16'h02_be] = 8'h90;
    buff [16'h02_bf] = 8'h1B;
    buff [16'h02_c0] = 8'h02;
    buff [16'h02_c1] = 8'h0A;
    buff [16'h02_c2] = 8'hF0;
    buff [16'h02_c3] = 8'h78;
    buff [16'h02_c4] = 8'h80;
    buff [16'h02_c5] = 8'h18;
    buff [16'h02_c6] = 8'h76;
    buff [16'h02_c7] = 8'h00;
    buff [16'h02_c8] = 8'hE8;
    buff [16'h02_c9] = 8'h70;
    buff [16'h02_ca] = 8'hFA;
    buff [16'h02_cb] = 8'h75;
    buff [16'h02_cc] = 8'hD0;
    buff [16'h02_cd] = 8'h00;
    buff [16'h02_ce] = 8'h74;
    buff [16'h02_cf] = 8'h20;
    buff [16'h02_d0] = 8'hB2;
    buff [16'h02_d1] = 8'hE5;
    buff [16'h02_d2] = 8'h60;
    buff [16'h02_d3] = 8'h06;
    buff [16'h02_d4] = 8'h75;
    buff [16'h02_d5] = 8'h90;
    buff [16'h02_d6] = 8'h1C;
    buff [16'h02_d7] = 8'h02;
    buff [16'h02_d8] = 8'h0A;
    buff [16'h02_d9] = 8'hF0;
    buff [16'h02_da] = 8'h78;
    buff [16'h02_db] = 8'h80;
    buff [16'h02_dc] = 8'h18;
    buff [16'h02_dd] = 8'h76;
    buff [16'h02_de] = 8'h00;
    buff [16'h02_df] = 8'hE8;
    buff [16'h02_e0] = 8'h70;
    buff [16'h02_e1] = 8'hFA;
    buff [16'h02_e2] = 8'h75;
    buff [16'h02_e3] = 8'hD0;
    buff [16'h02_e4] = 8'h00;
    buff [16'h02_e5] = 8'h74;
    buff [16'h02_e6] = 8'h80;
    buff [16'h02_e7] = 8'h24;
    buff [16'h02_e8] = 8'h99;
    buff [16'h02_e9] = 8'hD4;
    buff [16'h02_ea] = 8'h94;
    buff [16'h02_eb] = 8'h78;
    buff [16'h02_ec] = 8'h60;
    buff [16'h02_ed] = 8'h06;
    buff [16'h02_ee] = 8'h75;
    buff [16'h02_ef] = 8'h90;
    buff [16'h02_f0] = 8'h1D;
    buff [16'h02_f1] = 8'h02;
    buff [16'h02_f2] = 8'h0A;
    buff [16'h02_f3] = 8'hF0;
    buff [16'h02_f4] = 8'h78;
    buff [16'h02_f5] = 8'h80;
    buff [16'h02_f6] = 8'h18;
    buff [16'h02_f7] = 8'h76;
    buff [16'h02_f8] = 8'h00;
    buff [16'h02_f9] = 8'hE8;
    buff [16'h02_fa] = 8'h70;
    buff [16'h02_fb] = 8'hFA;
    buff [16'h02_fc] = 8'h75;
    buff [16'h02_fd] = 8'hD0;
    buff [16'h02_fe] = 8'h00;
    buff [16'h02_ff] = 8'h74;
    buff [16'h03_00] = 8'h0A;
    buff [16'h03_01] = 8'h14;
    buff [16'h03_02] = 8'h94;
    buff [16'h03_03] = 8'h09;
    buff [16'h03_04] = 8'h60;
    buff [16'h03_05] = 8'h06;
    buff [16'h03_06] = 8'h75;
    buff [16'h03_07] = 8'h90;
    buff [16'h03_08] = 8'h1E;
    buff [16'h03_09] = 8'h02;
    buff [16'h03_0a] = 8'h0A;
    buff [16'h03_0b] = 8'hF0;
    buff [16'h03_0c] = 8'h78;
    buff [16'h03_0d] = 8'h80;
    buff [16'h03_0e] = 8'h18;
    buff [16'h03_0f] = 8'h76;
    buff [16'h03_10] = 8'h00;
    buff [16'h03_11] = 8'hE8;
    buff [16'h03_12] = 8'h70;
    buff [16'h03_13] = 8'hFA;
    buff [16'h03_14] = 8'h75;
    buff [16'h03_15] = 8'hD0;
    buff [16'h03_16] = 8'h00;
    buff [16'h03_17] = 8'h78;
    buff [16'h03_18] = 8'h0A;
    buff [16'h03_19] = 8'h18;
    buff [16'h03_1a] = 8'hE8;
    buff [16'h03_1b] = 8'h94;
    buff [16'h03_1c] = 8'h09;
    buff [16'h03_1d] = 8'h60;
    buff [16'h03_1e] = 8'h06;
    buff [16'h03_1f] = 8'h75;
    buff [16'h03_20] = 8'h90;
    buff [16'h03_21] = 8'h1F;
    buff [16'h03_22] = 8'h02;
    buff [16'h03_23] = 8'h0A;
    buff [16'h03_24] = 8'hF0;
    buff [16'h03_25] = 8'h78;
    buff [16'h03_26] = 8'h80;
    buff [16'h03_27] = 8'h18;
    buff [16'h03_28] = 8'h76;
    buff [16'h03_29] = 8'h00;
    buff [16'h03_2a] = 8'hE8;
    buff [16'h03_2b] = 8'h70;
    buff [16'h03_2c] = 8'hFA;
    buff [16'h03_2d] = 8'h75;
    buff [16'h03_2e] = 8'hD0;
    buff [16'h03_2f] = 8'h00;
    buff [16'h03_30] = 8'h75;
    buff [16'h03_31] = 8'h7F;
    buff [16'h03_32] = 8'h0A;
    buff [16'h03_33] = 8'h15;
    buff [16'h03_34] = 8'h7F;
    buff [16'h03_35] = 8'hE5;
    buff [16'h03_36] = 8'h7F;
    buff [16'h03_37] = 8'h94;
    buff [16'h03_38] = 8'h09;
    buff [16'h03_39] = 8'h60;
    buff [16'h03_3a] = 8'h06;
    buff [16'h03_3b] = 8'h75;
    buff [16'h03_3c] = 8'h90;
    buff [16'h03_3d] = 8'h20;
    buff [16'h03_3e] = 8'h02;
    buff [16'h03_3f] = 8'h0A;
    buff [16'h03_40] = 8'hF0;
    buff [16'h03_41] = 8'h78;
    buff [16'h03_42] = 8'h80;
    buff [16'h03_43] = 8'h18;
    buff [16'h03_44] = 8'h76;
    buff [16'h03_45] = 8'h00;
    buff [16'h03_46] = 8'hE8;
    buff [16'h03_47] = 8'h70;
    buff [16'h03_48] = 8'hFA;
    buff [16'h03_49] = 8'h75;
    buff [16'h03_4a] = 8'hD0;
    buff [16'h03_4b] = 8'h00;
    buff [16'h03_4c] = 8'h78;
    buff [16'h03_4d] = 8'h7F;
    buff [16'h03_4e] = 8'h75;
    buff [16'h03_4f] = 8'h7F;
    buff [16'h03_50] = 8'h0A;
    buff [16'h03_51] = 8'h16;
    buff [16'h03_52] = 8'hE6;
    buff [16'h03_53] = 8'h94;
    buff [16'h03_54] = 8'h09;
    buff [16'h03_55] = 8'h60;
    buff [16'h03_56] = 8'h06;
    buff [16'h03_57] = 8'h75;
    buff [16'h03_58] = 8'h90;
    buff [16'h03_59] = 8'h21;
    buff [16'h03_5a] = 8'h02;
    buff [16'h03_5b] = 8'h0A;
    buff [16'h03_5c] = 8'hF0;
    buff [16'h03_5d] = 8'h78;
    buff [16'h03_5e] = 8'h80;
    buff [16'h03_5f] = 8'h18;
    buff [16'h03_60] = 8'h76;
    buff [16'h03_61] = 8'h00;
    buff [16'h03_62] = 8'hE8;
    buff [16'h03_63] = 8'h70;
    buff [16'h03_64] = 8'hFA;
    buff [16'h03_65] = 8'h75;
    buff [16'h03_66] = 8'hD0;
    buff [16'h03_67] = 8'h00;
    buff [16'h03_68] = 8'h74;
    buff [16'h03_69] = 8'hFB;
    buff [16'h03_6a] = 8'h75;
    buff [16'h03_6b] = 8'hF0;
    buff [16'h03_6c] = 8'h12;
    buff [16'h03_6d] = 8'h84;
    buff [16'h03_6e] = 8'h94;
    buff [16'h03_6f] = 8'h0D;
    buff [16'h03_70] = 8'h60;
    buff [16'h03_71] = 8'h03;
    buff [16'h03_72] = 8'h75;
    buff [16'h03_73] = 8'h90;
    buff [16'h03_74] = 8'h22;
    buff [16'h03_75] = 8'hE5;
    buff [16'h03_76] = 8'hF0;
    buff [16'h03_77] = 8'h94;
    buff [16'h03_78] = 8'h11;
    buff [16'h03_79] = 8'h60;
    buff [16'h03_7a] = 8'h06;
    buff [16'h03_7b] = 8'h75;
    buff [16'h03_7c] = 8'h90;
    buff [16'h03_7d] = 8'h22;
    buff [16'h03_7e] = 8'h02;
    buff [16'h03_7f] = 8'h0A;
    buff [16'h03_80] = 8'hF0;
    buff [16'h03_81] = 8'h78;
    buff [16'h03_82] = 8'h80;
    buff [16'h03_83] = 8'h18;
    buff [16'h03_84] = 8'h76;
    buff [16'h03_85] = 8'h00;
    buff [16'h03_86] = 8'hE8;
    buff [16'h03_87] = 8'h70;
    buff [16'h03_88] = 8'hFA;
    buff [16'h03_89] = 8'h75;
    buff [16'h03_8a] = 8'hD0;
    buff [16'h03_8b] = 8'h00;
    buff [16'h03_8c] = 8'h78;
    buff [16'h03_8d] = 8'h0A;
    buff [16'h03_8e] = 8'hD8;
    buff [16'h03_8f] = 8'h06;
    buff [16'h03_90] = 8'h75;
    buff [16'h03_91] = 8'h90;
    buff [16'h03_92] = 8'h23;
    buff [16'h03_93] = 8'h02;
    buff [16'h03_94] = 8'h0A;
    buff [16'h03_95] = 8'hF0;
    buff [16'h03_96] = 8'h78;
    buff [16'h03_97] = 8'h01;
    buff [16'h03_98] = 8'hD8;
    buff [16'h03_99] = 8'h02;
    buff [16'h03_9a] = 8'h61;
    buff [16'h03_9b] = 8'hA2;
    buff [16'h03_9c] = 8'h75;
    buff [16'h03_9d] = 8'h90;
    buff [16'h03_9e] = 8'h23;
    buff [16'h03_9f] = 8'h02;
    buff [16'h03_a0] = 8'h0A;
    buff [16'h03_a1] = 8'hF0;
    buff [16'h03_a2] = 8'h78;
    buff [16'h03_a3] = 8'h80;
    buff [16'h03_a4] = 8'h18;
    buff [16'h03_a5] = 8'h76;
    buff [16'h03_a6] = 8'h00;
    buff [16'h03_a7] = 8'hE8;
    buff [16'h03_a8] = 8'h70;
    buff [16'h03_a9] = 8'hFA;
    buff [16'h03_aa] = 8'h75;
    buff [16'h03_ab] = 8'hD0;
    buff [16'h03_ac] = 8'h00;
    buff [16'h03_ad] = 8'h75;
    buff [16'h03_ae] = 8'h7F;
    buff [16'h03_af] = 8'h0A;
    buff [16'h03_b0] = 8'hD5;
    buff [16'h03_b1] = 8'h7F;
    buff [16'h03_b2] = 8'h06;
    buff [16'h03_b3] = 8'h75;
    buff [16'h03_b4] = 8'h90;
    buff [16'h03_b5] = 8'h24;
    buff [16'h03_b6] = 8'h02;
    buff [16'h03_b7] = 8'h0A;
    buff [16'h03_b8] = 8'hF0;
    buff [16'h03_b9] = 8'h75;
    buff [16'h03_ba] = 8'h7F;
    buff [16'h03_bb] = 8'h01;
    buff [16'h03_bc] = 8'hD5;
    buff [16'h03_bd] = 8'h7F;
    buff [16'h03_be] = 8'h02;
    buff [16'h03_bf] = 8'h61;
    buff [16'h03_c0] = 8'hC7;
    buff [16'h03_c1] = 8'h75;
    buff [16'h03_c2] = 8'h90;
    buff [16'h03_c3] = 8'h24;
    buff [16'h03_c4] = 8'h02;
    buff [16'h03_c5] = 8'h0A;
    buff [16'h03_c6] = 8'hF0;
    buff [16'h03_c7] = 8'h78;
    buff [16'h03_c8] = 8'h80;
    buff [16'h03_c9] = 8'h18;
    buff [16'h03_ca] = 8'h76;
    buff [16'h03_cb] = 8'h00;
    buff [16'h03_cc] = 8'hE8;
    buff [16'h03_cd] = 8'h70;
    buff [16'h03_ce] = 8'hFA;
    buff [16'h03_cf] = 8'h75;
    buff [16'h03_d0] = 8'hD0;
    buff [16'h03_d1] = 8'h00;
    buff [16'h03_d2] = 8'h74;
    buff [16'h03_d3] = 8'h0A;
    buff [16'h03_d4] = 8'h04;
    buff [16'h03_d5] = 8'h94;
    buff [16'h03_d6] = 8'h0B;
    buff [16'h03_d7] = 8'h60;
    buff [16'h03_d8] = 8'h06;
    buff [16'h03_d9] = 8'h75;
    buff [16'h03_da] = 8'h90;
    buff [16'h03_db] = 8'h25;
    buff [16'h03_dc] = 8'h02;
    buff [16'h03_dd] = 8'h0A;
    buff [16'h03_de] = 8'hF0;
    buff [16'h03_df] = 8'h78;
    buff [16'h03_e0] = 8'h80;
    buff [16'h03_e1] = 8'h18;
    buff [16'h03_e2] = 8'h76;
    buff [16'h03_e3] = 8'h00;
    buff [16'h03_e4] = 8'hE8;
    buff [16'h03_e5] = 8'h70;
    buff [16'h03_e6] = 8'hFA;
    buff [16'h03_e7] = 8'h75;
    buff [16'h03_e8] = 8'hD0;
    buff [16'h03_e9] = 8'h00;
    buff [16'h03_ea] = 8'h78;
    buff [16'h03_eb] = 8'h0A;
    buff [16'h03_ec] = 8'h08;
    buff [16'h03_ed] = 8'hE8;
    buff [16'h03_ee] = 8'h94;
    buff [16'h03_ef] = 8'h0B;
    buff [16'h03_f0] = 8'h60;
    buff [16'h03_f1] = 8'h06;
    buff [16'h03_f2] = 8'h75;
    buff [16'h03_f3] = 8'h90;
    buff [16'h03_f4] = 8'h26;
    buff [16'h03_f5] = 8'h02;
    buff [16'h03_f6] = 8'h0A;
    buff [16'h03_f7] = 8'hF0;
    buff [16'h03_f8] = 8'h78;
    buff [16'h03_f9] = 8'h80;
    buff [16'h03_fa] = 8'h18;
    buff [16'h03_fb] = 8'h76;
    buff [16'h03_fc] = 8'h00;
    buff [16'h03_fd] = 8'hE8;
    buff [16'h03_fe] = 8'h70;
    buff [16'h03_ff] = 8'hFA;
    buff [16'h04_00] = 8'h75;
    buff [16'h04_01] = 8'hD0;
    buff [16'h04_02] = 8'h00;
    buff [16'h04_03] = 8'h75;
    buff [16'h04_04] = 8'h7F;
    buff [16'h04_05] = 8'h0A;
    buff [16'h04_06] = 8'h05;
    buff [16'h04_07] = 8'h7F;
    buff [16'h04_08] = 8'hE5;
    buff [16'h04_09] = 8'h7F;
    buff [16'h04_0a] = 8'h94;
    buff [16'h04_0b] = 8'h0B;
    buff [16'h04_0c] = 8'h60;
    buff [16'h04_0d] = 8'h06;
    buff [16'h04_0e] = 8'h75;
    buff [16'h04_0f] = 8'h90;
    buff [16'h04_10] = 8'h27;
    buff [16'h04_11] = 8'h02;
    buff [16'h04_12] = 8'h0A;
    buff [16'h04_13] = 8'hF0;
    buff [16'h04_14] = 8'h78;
    buff [16'h04_15] = 8'h80;
    buff [16'h04_16] = 8'h18;
    buff [16'h04_17] = 8'h76;
    buff [16'h04_18] = 8'h00;
    buff [16'h04_19] = 8'hE8;
    buff [16'h04_1a] = 8'h70;
    buff [16'h04_1b] = 8'hFA;
    buff [16'h04_1c] = 8'h75;
    buff [16'h04_1d] = 8'hD0;
    buff [16'h04_1e] = 8'h00;
    buff [16'h04_1f] = 8'h75;
    buff [16'h04_20] = 8'h7F;
    buff [16'h04_21] = 8'h0A;
    buff [16'h04_22] = 8'h78;
    buff [16'h04_23] = 8'h7F;
    buff [16'h04_24] = 8'h06;
    buff [16'h04_25] = 8'hE6;
    buff [16'h04_26] = 8'h94;
    buff [16'h04_27] = 8'h0B;
    buff [16'h04_28] = 8'h60;
    buff [16'h04_29] = 8'h06;
    buff [16'h04_2a] = 8'h75;
    buff [16'h04_2b] = 8'h90;
    buff [16'h04_2c] = 8'h28;
    buff [16'h04_2d] = 8'h02;
    buff [16'h04_2e] = 8'h0A;
    buff [16'h04_2f] = 8'hF0;
    buff [16'h04_30] = 8'h78;
    buff [16'h04_31] = 8'h80;
    buff [16'h04_32] = 8'h18;
    buff [16'h04_33] = 8'h76;
    buff [16'h04_34] = 8'h00;
    buff [16'h04_35] = 8'hE8;
    buff [16'h04_36] = 8'h70;
    buff [16'h04_37] = 8'hFA;
    buff [16'h04_38] = 8'h75;
    buff [16'h04_39] = 8'hD0;
    buff [16'h04_3a] = 8'h00;
    buff [16'h04_3b] = 8'h90;
    buff [16'h04_3c] = 8'h12;
    buff [16'h04_3d] = 8'hFF;
    buff [16'h04_3e] = 8'hA3;
    buff [16'h04_3f] = 8'hE5;
    buff [16'h04_40] = 8'h83;
    buff [16'h04_41] = 8'h94;
    buff [16'h04_42] = 8'h13;
    buff [16'h04_43] = 8'h60;
    buff [16'h04_44] = 8'h06;
    buff [16'h04_45] = 8'h75;
    buff [16'h04_46] = 8'h90;
    buff [16'h04_47] = 8'h29;
    buff [16'h04_48] = 8'h02;
    buff [16'h04_49] = 8'h0A;
    buff [16'h04_4a] = 8'hF0;
    buff [16'h04_4b] = 8'hE5;
    buff [16'h04_4c] = 8'h82;
    buff [16'h04_4d] = 8'h60;
    buff [16'h04_4e] = 8'h06;
    buff [16'h04_4f] = 8'h75;
    buff [16'h04_50] = 8'h90;
    buff [16'h04_51] = 8'h29;
    buff [16'h04_52] = 8'h02;
    buff [16'h04_53] = 8'h0A;
    buff [16'h04_54] = 8'hF0;
    buff [16'h04_55] = 8'h78;
    buff [16'h04_56] = 8'h80;
    buff [16'h04_57] = 8'h18;
    buff [16'h04_58] = 8'h76;
    buff [16'h04_59] = 8'h00;
    buff [16'h04_5a] = 8'hE8;
    buff [16'h04_5b] = 8'h70;
    buff [16'h04_5c] = 8'hFA;
    buff [16'h04_5d] = 8'h75;
    buff [16'h04_5e] = 8'hD0;
    buff [16'h04_5f] = 8'h00;
    buff [16'h04_60] = 8'h74;
    buff [16'h04_61] = 8'h10;
    buff [16'h04_62] = 8'h20;
    buff [16'h04_63] = 8'hE4;
    buff [16'h04_64] = 8'h06;
    buff [16'h04_65] = 8'h75;
    buff [16'h04_66] = 8'h90;
    buff [16'h04_67] = 8'h2A;
    buff [16'h04_68] = 8'h02;
    buff [16'h04_69] = 8'h0A;
    buff [16'h04_6a] = 8'hF0;
    buff [16'h04_6b] = 8'h78;
    buff [16'h04_6c] = 8'h80;
    buff [16'h04_6d] = 8'h18;
    buff [16'h04_6e] = 8'h76;
    buff [16'h04_6f] = 8'h00;
    buff [16'h04_70] = 8'hE8;
    buff [16'h04_71] = 8'h70;
    buff [16'h04_72] = 8'hFA;
    buff [16'h04_73] = 8'h75;
    buff [16'h04_74] = 8'hD0;
    buff [16'h04_75] = 8'h00;
    buff [16'h04_76] = 8'h74;
    buff [16'h04_77] = 8'h08;
    buff [16'h04_78] = 8'h10;
    buff [16'h04_79] = 8'hE3;
    buff [16'h04_7a] = 8'h06;
    buff [16'h04_7b] = 8'h75;
    buff [16'h04_7c] = 8'h90;
    buff [16'h04_7d] = 8'h2B;
    buff [16'h04_7e] = 8'h02;
    buff [16'h04_7f] = 8'h0A;
    buff [16'h04_80] = 8'hF0;
    buff [16'h04_81] = 8'h60;
    buff [16'h04_82] = 8'h06;
    buff [16'h04_83] = 8'h75;
    buff [16'h04_84] = 8'h90;
    buff [16'h04_85] = 8'h2B;
    buff [16'h04_86] = 8'h02;
    buff [16'h04_87] = 8'h0A;
    buff [16'h04_88] = 8'hF0;
    buff [16'h04_89] = 8'h78;
    buff [16'h04_8a] = 8'h80;
    buff [16'h04_8b] = 8'h18;
    buff [16'h04_8c] = 8'h76;
    buff [16'h04_8d] = 8'h00;
    buff [16'h04_8e] = 8'hE8;
    buff [16'h04_8f] = 8'h70;
    buff [16'h04_90] = 8'hFA;
    buff [16'h04_91] = 8'h75;
    buff [16'h04_92] = 8'hD0;
    buff [16'h04_93] = 8'h00;
    buff [16'h04_94] = 8'h40;
    buff [16'h04_95] = 8'h03;
    buff [16'h04_96] = 8'hB3;
    buff [16'h04_97] = 8'h40;
    buff [16'h04_98] = 8'h06;
    buff [16'h04_99] = 8'h75;
    buff [16'h04_9a] = 8'h90;
    buff [16'h04_9b] = 8'h2C;
    buff [16'h04_9c] = 8'h02;
    buff [16'h04_9d] = 8'h0A;
    buff [16'h04_9e] = 8'hF0;
    buff [16'h04_9f] = 8'h78;
    buff [16'h04_a0] = 8'h80;
    buff [16'h04_a1] = 8'h18;
    buff [16'h04_a2] = 8'h76;
    buff [16'h04_a3] = 8'h00;
    buff [16'h04_a4] = 8'hE8;
    buff [16'h04_a5] = 8'h70;
    buff [16'h04_a6] = 8'hFA;
    buff [16'h04_a7] = 8'h75;
    buff [16'h04_a8] = 8'hD0;
    buff [16'h04_a9] = 8'h00;
    buff [16'h04_aa] = 8'h74;
    buff [16'h04_ab] = 8'h04;
    buff [16'h04_ac] = 8'h90;
    buff [16'h04_ad] = 8'h04;
    buff [16'h04_ae] = 8'hB0;
    buff [16'h04_af] = 8'h73;
    buff [16'h04_b0] = 8'h81;
    buff [16'h04_b1] = 8'hB8;
    buff [16'h04_b2] = 8'h81;
    buff [16'h04_b3] = 8'hB8;
    buff [16'h04_b4] = 8'h81;
    buff [16'h04_b5] = 8'hBE;
    buff [16'h04_b6] = 8'h81;
    buff [16'h04_b7] = 8'hB8;
    buff [16'h04_b8] = 8'h75;
    buff [16'h04_b9] = 8'h90;
    buff [16'h04_ba] = 8'h2B;
    buff [16'h04_bb] = 8'h02;
    buff [16'h04_bc] = 8'h0A;
    buff [16'h04_bd] = 8'hF0;
    buff [16'h04_be] = 8'h78;
    buff [16'h04_bf] = 8'h80;
    buff [16'h04_c0] = 8'h18;
    buff [16'h04_c1] = 8'h76;
    buff [16'h04_c2] = 8'h00;
    buff [16'h04_c3] = 8'hE8;
    buff [16'h04_c4] = 8'h70;
    buff [16'h04_c5] = 8'hFA;
    buff [16'h04_c6] = 8'h75;
    buff [16'h04_c7] = 8'hD0;
    buff [16'h04_c8] = 8'h00;
    buff [16'h04_c9] = 8'h74;
    buff [16'h04_ca] = 8'h04;
    buff [16'h04_cb] = 8'h30;
    buff [16'h04_cc] = 8'hE2;
    buff [16'h04_cd] = 8'h03;
    buff [16'h04_ce] = 8'h30;
    buff [16'h04_cf] = 8'hE1;
    buff [16'h04_d0] = 8'h06;
    buff [16'h04_d1] = 8'h75;
    buff [16'h04_d2] = 8'h90;
    buff [16'h04_d3] = 8'h2E;
    buff [16'h04_d4] = 8'h02;
    buff [16'h04_d5] = 8'h0A;
    buff [16'h04_d6] = 8'hF0;
    buff [16'h04_d7] = 8'h78;
    buff [16'h04_d8] = 8'h80;
    buff [16'h04_d9] = 8'h18;
    buff [16'h04_da] = 8'h76;
    buff [16'h04_db] = 8'h00;
    buff [16'h04_dc] = 8'hE8;
    buff [16'h04_dd] = 8'h70;
    buff [16'h04_de] = 8'hFA;
    buff [16'h04_df] = 8'h75;
    buff [16'h04_e0] = 8'hD0;
    buff [16'h04_e1] = 8'h00;
    buff [16'h04_e2] = 8'hB3;
    buff [16'h04_e3] = 8'h50;
    buff [16'h04_e4] = 8'h03;
    buff [16'h04_e5] = 8'hB3;
    buff [16'h04_e6] = 8'h50;
    buff [16'h04_e7] = 8'h06;
    buff [16'h04_e8] = 8'h75;
    buff [16'h04_e9] = 8'h90;
    buff [16'h04_ea] = 8'h2F;
    buff [16'h04_eb] = 8'h02;
    buff [16'h04_ec] = 8'h0A;
    buff [16'h04_ed] = 8'hF0;
    buff [16'h04_ee] = 8'h78;
    buff [16'h04_ef] = 8'h80;
    buff [16'h04_f0] = 8'h18;
    buff [16'h04_f1] = 8'h76;
    buff [16'h04_f2] = 8'h00;
    buff [16'h04_f3] = 8'hE8;
    buff [16'h04_f4] = 8'h70;
    buff [16'h04_f5] = 8'hFA;
    buff [16'h04_f6] = 8'h75;
    buff [16'h04_f7] = 8'hD0;
    buff [16'h04_f8] = 8'h00;
    buff [16'h04_f9] = 8'h70;
    buff [16'h04_fa] = 8'h04;
    buff [16'h04_fb] = 8'h74;
    buff [16'h04_fc] = 8'h01;
    buff [16'h04_fd] = 8'h70;
    buff [16'h04_fe] = 8'h06;
    buff [16'h04_ff] = 8'h75;
    buff [16'h05_00] = 8'h90;
    buff [16'h05_01] = 8'h30;
    buff [16'h05_02] = 8'h02;
    buff [16'h05_03] = 8'h0A;
    buff [16'h05_04] = 8'hF0;
    buff [16'h05_05] = 8'h78;
    buff [16'h05_06] = 8'h80;
    buff [16'h05_07] = 8'h18;
    buff [16'h05_08] = 8'h76;
    buff [16'h05_09] = 8'h00;
    buff [16'h05_0a] = 8'hE8;
    buff [16'h05_0b] = 8'h70;
    buff [16'h05_0c] = 8'hFA;
    buff [16'h05_0d] = 8'h75;
    buff [16'h05_0e] = 8'hD0;
    buff [16'h05_0f] = 8'h00;
    buff [16'h05_10] = 8'h74;
    buff [16'h05_11] = 8'h02;
    buff [16'h05_12] = 8'h60;
    buff [16'h05_13] = 8'h04;
    buff [16'h05_14] = 8'h74;
    buff [16'h05_15] = 8'h00;
    buff [16'h05_16] = 8'h60;
    buff [16'h05_17] = 8'h06;
    buff [16'h05_18] = 8'h75;
    buff [16'h05_19] = 8'h90;
    buff [16'h05_1a] = 8'h31;
    buff [16'h05_1b] = 8'h02;
    buff [16'h05_1c] = 8'h0A;
    buff [16'h05_1d] = 8'hF0;
    buff [16'h05_1e] = 8'h78;
    buff [16'h05_1f] = 8'h80;
    buff [16'h05_20] = 8'h18;
    buff [16'h05_21] = 8'h76;
    buff [16'h05_22] = 8'h00;
    buff [16'h05_23] = 8'hE8;
    buff [16'h05_24] = 8'h70;
    buff [16'h05_25] = 8'hFA;
    buff [16'h05_26] = 8'h75;
    buff [16'h05_27] = 8'hD0;
    buff [16'h05_28] = 8'h00;
    buff [16'h05_29] = 8'h02;
    buff [16'h05_2a] = 8'h05;
    buff [16'h05_2b] = 8'h32;
    buff [16'h05_2c] = 8'h75;
    buff [16'h05_2d] = 8'h90;
    buff [16'h05_2e] = 8'h33;
    buff [16'h05_2f] = 8'h02;
    buff [16'h05_30] = 8'h0A;
    buff [16'h05_31] = 8'hF0;
    buff [16'h05_32] = 8'h78;
    buff [16'h05_33] = 8'h80;
    buff [16'h05_34] = 8'h18;
    buff [16'h05_35] = 8'h76;
    buff [16'h05_36] = 8'h00;
    buff [16'h05_37] = 8'hE8;
    buff [16'h05_38] = 8'h70;
    buff [16'h05_39] = 8'hFA;
    buff [16'h05_3a] = 8'h75;
    buff [16'h05_3b] = 8'hD0;
    buff [16'h05_3c] = 8'h00;
    buff [16'h05_3d] = 8'h78;
    buff [16'h05_3e] = 8'h0A;
    buff [16'h05_3f] = 8'hE8;
    buff [16'h05_40] = 8'h94;
    buff [16'h05_41] = 8'h0A;
    buff [16'h05_42] = 8'h60;
    buff [16'h05_43] = 8'h06;
    buff [16'h05_44] = 8'h75;
    buff [16'h05_45] = 8'h90;
    buff [16'h05_46] = 8'h34;
    buff [16'h05_47] = 8'h02;
    buff [16'h05_48] = 8'h0A;
    buff [16'h05_49] = 8'hF0;
    buff [16'h05_4a] = 8'h78;
    buff [16'h05_4b] = 8'h80;
    buff [16'h05_4c] = 8'h18;
    buff [16'h05_4d] = 8'h76;
    buff [16'h05_4e] = 8'h00;
    buff [16'h05_4f] = 8'hE8;
    buff [16'h05_50] = 8'h70;
    buff [16'h05_51] = 8'hFA;
    buff [16'h05_52] = 8'h75;
    buff [16'h05_53] = 8'hD0;
    buff [16'h05_54] = 8'h00;
    buff [16'h05_55] = 8'h75;
    buff [16'h05_56] = 8'h7F;
    buff [16'h05_57] = 8'h0A;
    buff [16'h05_58] = 8'hE5;
    buff [16'h05_59] = 8'h7F;
    buff [16'h05_5a] = 8'h94;
    buff [16'h05_5b] = 8'h0A;
    buff [16'h05_5c] = 8'h60;
    buff [16'h05_5d] = 8'h06;
    buff [16'h05_5e] = 8'h75;
    buff [16'h05_5f] = 8'h90;
    buff [16'h05_60] = 8'h35;
    buff [16'h05_61] = 8'h02;
    buff [16'h05_62] = 8'h0A;
    buff [16'h05_63] = 8'hF0;
    buff [16'h05_64] = 8'h78;
    buff [16'h05_65] = 8'h80;
    buff [16'h05_66] = 8'h18;
    buff [16'h05_67] = 8'h76;
    buff [16'h05_68] = 8'h00;
    buff [16'h05_69] = 8'hE8;
    buff [16'h05_6a] = 8'h70;
    buff [16'h05_6b] = 8'hFA;
    buff [16'h05_6c] = 8'h75;
    buff [16'h05_6d] = 8'hD0;
    buff [16'h05_6e] = 8'h00;
    buff [16'h05_6f] = 8'h78;
    buff [16'h05_70] = 8'h7F;
    buff [16'h05_71] = 8'h75;
    buff [16'h05_72] = 8'h7F;
    buff [16'h05_73] = 8'h0A;
    buff [16'h05_74] = 8'hE6;
    buff [16'h05_75] = 8'h94;
    buff [16'h05_76] = 8'h0A;
    buff [16'h05_77] = 8'h60;
    buff [16'h05_78] = 8'h06;
    buff [16'h05_79] = 8'h75;
    buff [16'h05_7a] = 8'h90;
    buff [16'h05_7b] = 8'h36;
    buff [16'h05_7c] = 8'h02;
    buff [16'h05_7d] = 8'h0A;
    buff [16'h05_7e] = 8'hF0;
    buff [16'h05_7f] = 8'h78;
    buff [16'h05_80] = 8'h80;
    buff [16'h05_81] = 8'h18;
    buff [16'h05_82] = 8'h76;
    buff [16'h05_83] = 8'h00;
    buff [16'h05_84] = 8'hE8;
    buff [16'h05_85] = 8'h70;
    buff [16'h05_86] = 8'hFA;
    buff [16'h05_87] = 8'h75;
    buff [16'h05_88] = 8'hD0;
    buff [16'h05_89] = 8'h00;
    buff [16'h05_8a] = 8'h74;
    buff [16'h05_8b] = 8'h0A;
    buff [16'h05_8c] = 8'h94;
    buff [16'h05_8d] = 8'h0A;
    buff [16'h05_8e] = 8'h60;
    buff [16'h05_8f] = 8'h06;
    buff [16'h05_90] = 8'h75;
    buff [16'h05_91] = 8'h90;
    buff [16'h05_92] = 8'h37;
    buff [16'h05_93] = 8'h02;
    buff [16'h05_94] = 8'h0A;
    buff [16'h05_95] = 8'hF0;
    buff [16'h05_96] = 8'h78;
    buff [16'h05_97] = 8'h80;
    buff [16'h05_98] = 8'h18;
    buff [16'h05_99] = 8'h76;
    buff [16'h05_9a] = 8'h00;
    buff [16'h05_9b] = 8'hE8;
    buff [16'h05_9c] = 8'h70;
    buff [16'h05_9d] = 8'hFA;
    buff [16'h05_9e] = 8'h75;
    buff [16'h05_9f] = 8'hD0;
    buff [16'h05_a0] = 8'h00;
    buff [16'h05_a1] = 8'h74;
    buff [16'h05_a2] = 8'h0A;
    buff [16'h05_a3] = 8'hF8;
    buff [16'h05_a4] = 8'hE4;
    buff [16'h05_a5] = 8'hE8;
    buff [16'h05_a6] = 8'h94;
    buff [16'h05_a7] = 8'h0A;
    buff [16'h05_a8] = 8'h60;
    buff [16'h05_a9] = 8'h06;
    buff [16'h05_aa] = 8'h75;
    buff [16'h05_ab] = 8'h90;
    buff [16'h05_ac] = 8'h38;
    buff [16'h05_ad] = 8'h02;
    buff [16'h05_ae] = 8'h0A;
    buff [16'h05_af] = 8'hF0;
    buff [16'h05_b0] = 8'h78;
    buff [16'h05_b1] = 8'h80;
    buff [16'h05_b2] = 8'h18;
    buff [16'h05_b3] = 8'h76;
    buff [16'h05_b4] = 8'h00;
    buff [16'h05_b5] = 8'hE8;
    buff [16'h05_b6] = 8'h70;
    buff [16'h05_b7] = 8'hFA;
    buff [16'h05_b8] = 8'h75;
    buff [16'h05_b9] = 8'hD0;
    buff [16'h05_ba] = 8'h00;
    buff [16'h05_bb] = 8'h75;
    buff [16'h05_bc] = 8'h7F;
    buff [16'h05_bd] = 8'h0A;
    buff [16'h05_be] = 8'hA8;
    buff [16'h05_bf] = 8'h7F;
    buff [16'h05_c0] = 8'hE8;
    buff [16'h05_c1] = 8'h94;
    buff [16'h05_c2] = 8'h0A;
    buff [16'h05_c3] = 8'h60;
    buff [16'h05_c4] = 8'h06;
    buff [16'h05_c5] = 8'h75;
    buff [16'h05_c6] = 8'h90;
    buff [16'h05_c7] = 8'h39;
    buff [16'h05_c8] = 8'h02;
    buff [16'h05_c9] = 8'h0A;
    buff [16'h05_ca] = 8'hF0;
    buff [16'h05_cb] = 8'h78;
    buff [16'h05_cc] = 8'h80;
    buff [16'h05_cd] = 8'h18;
    buff [16'h05_ce] = 8'h76;
    buff [16'h05_cf] = 8'h00;
    buff [16'h05_d0] = 8'hE8;
    buff [16'h05_d1] = 8'h70;
    buff [16'h05_d2] = 8'hFA;
    buff [16'h05_d3] = 8'h75;
    buff [16'h05_d4] = 8'hD0;
    buff [16'h05_d5] = 8'h00;
    buff [16'h05_d6] = 8'h78;
    buff [16'h05_d7] = 8'h0A;
    buff [16'h05_d8] = 8'hE8;
    buff [16'h05_d9] = 8'h94;
    buff [16'h05_da] = 8'h0A;
    buff [16'h05_db] = 8'h60;
    buff [16'h05_dc] = 8'h06;
    buff [16'h05_dd] = 8'h75;
    buff [16'h05_de] = 8'h90;
    buff [16'h05_df] = 8'h3A;
    buff [16'h05_e0] = 8'h02;
    buff [16'h05_e1] = 8'h0A;
    buff [16'h05_e2] = 8'hF0;
    buff [16'h05_e3] = 8'h78;
    buff [16'h05_e4] = 8'h80;
    buff [16'h05_e5] = 8'h18;
    buff [16'h05_e6] = 8'h76;
    buff [16'h05_e7] = 8'h00;
    buff [16'h05_e8] = 8'hE8;
    buff [16'h05_e9] = 8'h70;
    buff [16'h05_ea] = 8'hFA;
    buff [16'h05_eb] = 8'h75;
    buff [16'h05_ec] = 8'hD0;
    buff [16'h05_ed] = 8'h00;
    buff [16'h05_ee] = 8'h74;
    buff [16'h05_ef] = 8'h0A;
    buff [16'h05_f0] = 8'hF5;
    buff [16'h05_f1] = 8'h7F;
    buff [16'h05_f2] = 8'hE4;
    buff [16'h05_f3] = 8'hE5;
    buff [16'h05_f4] = 8'h7F;
    buff [16'h05_f5] = 8'h94;
    buff [16'h05_f6] = 8'h0A;
    buff [16'h05_f7] = 8'h60;
    buff [16'h05_f8] = 8'h06;
    buff [16'h05_f9] = 8'h75;
    buff [16'h05_fa] = 8'h90;
    buff [16'h05_fb] = 8'h3B;
    buff [16'h05_fc] = 8'h02;
    buff [16'h05_fd] = 8'h0A;
    buff [16'h05_fe] = 8'hF0;
    buff [16'h05_ff] = 8'h78;
    buff [16'h06_00] = 8'h80;
    buff [16'h06_01] = 8'h18;
    buff [16'h06_02] = 8'h76;
    buff [16'h06_03] = 8'h00;
    buff [16'h06_04] = 8'hE8;
    buff [16'h06_05] = 8'h70;
    buff [16'h06_06] = 8'hFA;
    buff [16'h06_07] = 8'h75;
    buff [16'h06_08] = 8'hD0;
    buff [16'h06_09] = 8'h00;
    buff [16'h06_0a] = 8'h78;
    buff [16'h06_0b] = 8'h0A;
    buff [16'h06_0c] = 8'h88;
    buff [16'h06_0d] = 8'h7F;
    buff [16'h06_0e] = 8'hE5;
    buff [16'h06_0f] = 8'h7F;
    buff [16'h06_10] = 8'h94;
    buff [16'h06_11] = 8'h0A;
    buff [16'h06_12] = 8'h60;
    buff [16'h06_13] = 8'h06;
    buff [16'h06_14] = 8'h75;
    buff [16'h06_15] = 8'h90;
    buff [16'h06_16] = 8'h3C;
    buff [16'h06_17] = 8'h02;
    buff [16'h06_18] = 8'h0A;
    buff [16'h06_19] = 8'hF0;
    buff [16'h06_1a] = 8'h78;
    buff [16'h06_1b] = 8'h80;
    buff [16'h06_1c] = 8'h18;
    buff [16'h06_1d] = 8'h76;
    buff [16'h06_1e] = 8'h00;
    buff [16'h06_1f] = 8'hE8;
    buff [16'h06_20] = 8'h70;
    buff [16'h06_21] = 8'hFA;
    buff [16'h06_22] = 8'h75;
    buff [16'h06_23] = 8'hD0;
    buff [16'h06_24] = 8'h00;
    buff [16'h06_25] = 8'h75;
    buff [16'h06_26] = 8'h7F;
    buff [16'h06_27] = 8'h0A;
    buff [16'h06_28] = 8'h85;
    buff [16'h06_29] = 8'h7F;
    buff [16'h06_2a] = 8'h7E;
    buff [16'h06_2b] = 8'hE5;
    buff [16'h06_2c] = 8'h7E;
    buff [16'h06_2d] = 8'h94;
    buff [16'h06_2e] = 8'h0A;
    buff [16'h06_2f] = 8'h60;
    buff [16'h06_30] = 8'h06;
    buff [16'h06_31] = 8'h75;
    buff [16'h06_32] = 8'h90;
    buff [16'h06_33] = 8'h3D;
    buff [16'h06_34] = 8'h02;
    buff [16'h06_35] = 8'h0A;
    buff [16'h06_36] = 8'hF0;
    buff [16'h06_37] = 8'h78;
    buff [16'h06_38] = 8'h80;
    buff [16'h06_39] = 8'h18;
    buff [16'h06_3a] = 8'h76;
    buff [16'h06_3b] = 8'h00;
    buff [16'h06_3c] = 8'hE8;
    buff [16'h06_3d] = 8'h70;
    buff [16'h06_3e] = 8'hFA;
    buff [16'h06_3f] = 8'h75;
    buff [16'h06_40] = 8'hD0;
    buff [16'h06_41] = 8'h00;
    buff [16'h06_42] = 8'h75;
    buff [16'h06_43] = 8'h7F;
    buff [16'h06_44] = 8'h0A;
    buff [16'h06_45] = 8'h78;
    buff [16'h06_46] = 8'h7F;
    buff [16'h06_47] = 8'h86;
    buff [16'h06_48] = 8'h7E;
    buff [16'h06_49] = 8'hE5;
    buff [16'h06_4a] = 8'h7E;
    buff [16'h06_4b] = 8'h94;
    buff [16'h06_4c] = 8'h0A;
    buff [16'h06_4d] = 8'h60;
    buff [16'h06_4e] = 8'h06;
    buff [16'h06_4f] = 8'h75;
    buff [16'h06_50] = 8'h90;
    buff [16'h06_51] = 8'h3E;
    buff [16'h06_52] = 8'h02;
    buff [16'h06_53] = 8'h0A;
    buff [16'h06_54] = 8'hF0;
    buff [16'h06_55] = 8'h78;
    buff [16'h06_56] = 8'h80;
    buff [16'h06_57] = 8'h18;
    buff [16'h06_58] = 8'h76;
    buff [16'h06_59] = 8'h00;
    buff [16'h06_5a] = 8'hE8;
    buff [16'h06_5b] = 8'h70;
    buff [16'h06_5c] = 8'hFA;
    buff [16'h06_5d] = 8'h75;
    buff [16'h06_5e] = 8'hD0;
    buff [16'h06_5f] = 8'h00;
    buff [16'h06_60] = 8'h75;
    buff [16'h06_61] = 8'h7F;
    buff [16'h06_62] = 8'h0A;
    buff [16'h06_63] = 8'hE5;
    buff [16'h06_64] = 8'h7F;
    buff [16'h06_65] = 8'h94;
    buff [16'h06_66] = 8'h0A;
    buff [16'h06_67] = 8'h60;
    buff [16'h06_68] = 8'h06;
    buff [16'h06_69] = 8'h75;
    buff [16'h06_6a] = 8'h90;
    buff [16'h06_6b] = 8'h3F;
    buff [16'h06_6c] = 8'h02;
    buff [16'h06_6d] = 8'h0A;
    buff [16'h06_6e] = 8'hF0;
    buff [16'h06_6f] = 8'h78;
    buff [16'h06_70] = 8'h80;
    buff [16'h06_71] = 8'h18;
    buff [16'h06_72] = 8'h76;
    buff [16'h06_73] = 8'h00;
    buff [16'h06_74] = 8'hE8;
    buff [16'h06_75] = 8'h70;
    buff [16'h06_76] = 8'hFA;
    buff [16'h06_77] = 8'h75;
    buff [16'h06_78] = 8'hD0;
    buff [16'h06_79] = 8'h00;
    buff [16'h06_7a] = 8'h74;
    buff [16'h06_7b] = 8'h0A;
    buff [16'h06_7c] = 8'h78;
    buff [16'h06_7d] = 8'h7F;
    buff [16'h06_7e] = 8'hF6;
    buff [16'h06_7f] = 8'hE4;
    buff [16'h06_80] = 8'hE5;
    buff [16'h06_81] = 8'h7F;
    buff [16'h06_82] = 8'h94;
    buff [16'h06_83] = 8'h0A;
    buff [16'h06_84] = 8'h60;
    buff [16'h06_85] = 8'h06;
    buff [16'h06_86] = 8'h75;
    buff [16'h06_87] = 8'h90;
    buff [16'h06_88] = 8'h40;
    buff [16'h06_89] = 8'h02;
    buff [16'h06_8a] = 8'h0A;
    buff [16'h06_8b] = 8'hF0;
    buff [16'h06_8c] = 8'h78;
    buff [16'h06_8d] = 8'h80;
    buff [16'h06_8e] = 8'h18;
    buff [16'h06_8f] = 8'h76;
    buff [16'h06_90] = 8'h00;
    buff [16'h06_91] = 8'hE8;
    buff [16'h06_92] = 8'h70;
    buff [16'h06_93] = 8'hFA;
    buff [16'h06_94] = 8'h75;
    buff [16'h06_95] = 8'hD0;
    buff [16'h06_96] = 8'h00;
    buff [16'h06_97] = 8'h75;
    buff [16'h06_98] = 8'h7F;
    buff [16'h06_99] = 8'h0A;
    buff [16'h06_9a] = 8'h78;
    buff [16'h06_9b] = 8'h7E;
    buff [16'h06_9c] = 8'hA6;
    buff [16'h06_9d] = 8'h7F;
    buff [16'h06_9e] = 8'hE5;
    buff [16'h06_9f] = 8'h7E;
    buff [16'h06_a0] = 8'h94;
    buff [16'h06_a1] = 8'h0A;
    buff [16'h06_a2] = 8'h60;
    buff [16'h06_a3] = 8'h06;
    buff [16'h06_a4] = 8'h75;
    buff [16'h06_a5] = 8'h90;
    buff [16'h06_a6] = 8'h41;
    buff [16'h06_a7] = 8'h02;
    buff [16'h06_a8] = 8'h0A;
    buff [16'h06_a9] = 8'hF0;
    buff [16'h06_aa] = 8'h78;
    buff [16'h06_ab] = 8'h80;
    buff [16'h06_ac] = 8'h18;
    buff [16'h06_ad] = 8'h76;
    buff [16'h06_ae] = 8'h00;
    buff [16'h06_af] = 8'hE8;
    buff [16'h06_b0] = 8'h70;
    buff [16'h06_b1] = 8'hFA;
    buff [16'h06_b2] = 8'h75;
    buff [16'h06_b3] = 8'hD0;
    buff [16'h06_b4] = 8'h00;
    buff [16'h06_b5] = 8'h78;
    buff [16'h06_b6] = 8'h7F;
    buff [16'h06_b7] = 8'h76;
    buff [16'h06_b8] = 8'h0A;
    buff [16'h06_b9] = 8'hE5;
    buff [16'h06_ba] = 8'h7F;
    buff [16'h06_bb] = 8'h94;
    buff [16'h06_bc] = 8'h0A;
    buff [16'h06_bd] = 8'h60;
    buff [16'h06_be] = 8'h06;
    buff [16'h06_bf] = 8'h75;
    buff [16'h06_c0] = 8'h90;
    buff [16'h06_c1] = 8'h42;
    buff [16'h06_c2] = 8'h02;
    buff [16'h06_c3] = 8'h0A;
    buff [16'h06_c4] = 8'hF0;
    buff [16'h06_c5] = 8'h78;
    buff [16'h06_c6] = 8'h80;
    buff [16'h06_c7] = 8'h18;
    buff [16'h06_c8] = 8'h76;
    buff [16'h06_c9] = 8'h00;
    buff [16'h06_ca] = 8'hE8;
    buff [16'h06_cb] = 8'h70;
    buff [16'h06_cc] = 8'hFA;
    buff [16'h06_cd] = 8'h75;
    buff [16'h06_ce] = 8'hD0;
    buff [16'h06_cf] = 8'h00;
    buff [16'h06_d0] = 8'h74;
    buff [16'h06_d1] = 8'h01;
    buff [16'h06_d2] = 8'hA2;
    buff [16'h06_d3] = 8'hE0;
    buff [16'h06_d4] = 8'h40;
    buff [16'h06_d5] = 8'h06;
    buff [16'h06_d6] = 8'h75;
    buff [16'h06_d7] = 8'h90;
    buff [16'h06_d8] = 8'h43;
    buff [16'h06_d9] = 8'h02;
    buff [16'h06_da] = 8'h0A;
    buff [16'h06_db] = 8'hF0;
    buff [16'h06_dc] = 8'h78;
    buff [16'h06_dd] = 8'h80;
    buff [16'h06_de] = 8'h18;
    buff [16'h06_df] = 8'h76;
    buff [16'h06_e0] = 8'h00;
    buff [16'h06_e1] = 8'hE8;
    buff [16'h06_e2] = 8'h70;
    buff [16'h06_e3] = 8'hFA;
    buff [16'h06_e4] = 8'h75;
    buff [16'h06_e5] = 8'hD0;
    buff [16'h06_e6] = 8'h00;
    buff [16'h06_e7] = 8'hB3;
    buff [16'h06_e8] = 8'h92;
    buff [16'h06_e9] = 8'hE0;
    buff [16'h06_ea] = 8'hB3;
    buff [16'h06_eb] = 8'h94;
    buff [16'h06_ec] = 8'h01;
    buff [16'h06_ed] = 8'h60;
    buff [16'h06_ee] = 8'h06;
    buff [16'h06_ef] = 8'h75;
    buff [16'h06_f0] = 8'h90;
    buff [16'h06_f1] = 8'h44;
    buff [16'h06_f2] = 8'h02;
    buff [16'h06_f3] = 8'h0A;
    buff [16'h06_f4] = 8'hF0;
    buff [16'h06_f5] = 8'h78;
    buff [16'h06_f6] = 8'h80;
    buff [16'h06_f7] = 8'h18;
    buff [16'h06_f8] = 8'h76;
    buff [16'h06_f9] = 8'h00;
    buff [16'h06_fa] = 8'hE8;
    buff [16'h06_fb] = 8'h70;
    buff [16'h06_fc] = 8'hFA;
    buff [16'h06_fd] = 8'h75;
    buff [16'h06_fe] = 8'hD0;
    buff [16'h06_ff] = 8'h00;
    buff [16'h07_00] = 8'h90;
    buff [16'h07_01] = 8'h12;
    buff [16'h07_02] = 8'h34;
    buff [16'h07_03] = 8'hE5;
    buff [16'h07_04] = 8'h83;
    buff [16'h07_05] = 8'h94;
    buff [16'h07_06] = 8'h12;
    buff [16'h07_07] = 8'h70;
    buff [16'h07_08] = 8'h06;
    buff [16'h07_09] = 8'hE5;
    buff [16'h07_0a] = 8'h82;
    buff [16'h07_0b] = 8'h94;
    buff [16'h07_0c] = 8'h34;
    buff [16'h07_0d] = 8'h60;
    buff [16'h07_0e] = 8'h06;
    buff [16'h07_0f] = 8'h75;
    buff [16'h07_10] = 8'h90;
    buff [16'h07_11] = 8'h45;
    buff [16'h07_12] = 8'h02;
    buff [16'h07_13] = 8'h0A;
    buff [16'h07_14] = 8'hF0;
    buff [16'h07_15] = 8'h78;
    buff [16'h07_16] = 8'h80;
    buff [16'h07_17] = 8'h18;
    buff [16'h07_18] = 8'h76;
    buff [16'h07_19] = 8'h00;
    buff [16'h07_1a] = 8'hE8;
    buff [16'h07_1b] = 8'h70;
    buff [16'h07_1c] = 8'hFA;
    buff [16'h07_1d] = 8'h75;
    buff [16'h07_1e] = 8'hD0;
    buff [16'h07_1f] = 8'h00;
    buff [16'h07_20] = 8'h90;
    buff [16'h07_21] = 8'h07;
    buff [16'h07_22] = 8'h31;
    buff [16'h07_23] = 8'h93;
    buff [16'h07_24] = 8'h94;
    buff [16'h07_25] = 8'h66;
    buff [16'h07_26] = 8'h70;
    buff [16'h07_27] = 8'h0B;
    buff [16'h07_28] = 8'h74;
    buff [16'h07_29] = 8'h01;
    buff [16'h07_2a] = 8'h93;
    buff [16'h07_2b] = 8'h94;
    buff [16'h07_2c] = 8'h77;
    buff [16'h07_2d] = 8'h60;
    buff [16'h07_2e] = 8'h0A;
    buff [16'h07_2f] = 8'h70;
    buff [16'h07_30] = 8'h02;
    buff [16'h07_31] = 8'h66;
    buff [16'h07_32] = 8'h77;
    buff [16'h07_33] = 8'h75;
    buff [16'h07_34] = 8'h90;
    buff [16'h07_35] = 8'h46;
    buff [16'h07_36] = 8'h02;
    buff [16'h07_37] = 8'h0A;
    buff [16'h07_38] = 8'hF0;
    buff [16'h07_39] = 8'h78;
    buff [16'h07_3a] = 8'h80;
    buff [16'h07_3b] = 8'h18;
    buff [16'h07_3c] = 8'h76;
    buff [16'h07_3d] = 8'h00;
    buff [16'h07_3e] = 8'hE8;
    buff [16'h07_3f] = 8'h70;
    buff [16'h07_40] = 8'hFA;
    buff [16'h07_41] = 8'h75;
    buff [16'h07_42] = 8'hD0;
    buff [16'h07_43] = 8'h00;
    buff [16'h07_44] = 8'h74;
    buff [16'h07_45] = 8'h0D;
    buff [16'h07_46] = 8'h83;
    buff [16'h07_47] = 8'h94;
    buff [16'h07_48] = 8'h66;
    buff [16'h07_49] = 8'h70;
    buff [16'h07_4a] = 8'h0B;
    buff [16'h07_4b] = 8'h74;
    buff [16'h07_4c] = 8'h07;
    buff [16'h07_4d] = 8'h83;
    buff [16'h07_4e] = 8'h94;
    buff [16'h07_4f] = 8'h77;
    buff [16'h07_50] = 8'h60;
    buff [16'h07_51] = 8'h0A;
    buff [16'h07_52] = 8'h70;
    buff [16'h07_53] = 8'h02;
    buff [16'h07_54] = 8'h66;
    buff [16'h07_55] = 8'h77;
    buff [16'h07_56] = 8'h75;
    buff [16'h07_57] = 8'h90;
    buff [16'h07_58] = 8'h47;
    buff [16'h07_59] = 8'h02;
    buff [16'h07_5a] = 8'h0A;
    buff [16'h07_5b] = 8'hF0;
    buff [16'h07_5c] = 8'h78;
    buff [16'h07_5d] = 8'h80;
    buff [16'h07_5e] = 8'h18;
    buff [16'h07_5f] = 8'h76;
    buff [16'h07_60] = 8'h00;
    buff [16'h07_61] = 8'hE8;
    buff [16'h07_62] = 8'h70;
    buff [16'h07_63] = 8'hFA;
    buff [16'h07_64] = 8'h75;
    buff [16'h07_65] = 8'hD0;
    buff [16'h07_66] = 8'h00;
    buff [16'h07_67] = 8'h74;
    buff [16'h07_68] = 8'h50;
    buff [16'h07_69] = 8'h75;
    buff [16'h07_6a] = 8'hF0;
    buff [16'h07_6b] = 8'hA0;
    buff [16'h07_6c] = 8'hA4;
    buff [16'h07_6d] = 8'h70;
    buff [16'h07_6e] = 8'h06;
    buff [16'h07_6f] = 8'hE5;
    buff [16'h07_70] = 8'hF0;
    buff [16'h07_71] = 8'h94;
    buff [16'h07_72] = 8'h32;
    buff [16'h07_73] = 8'h60;
    buff [16'h07_74] = 8'h06;
    buff [16'h07_75] = 8'h75;
    buff [16'h07_76] = 8'h90;
    buff [16'h07_77] = 8'h4C;
    buff [16'h07_78] = 8'h02;
    buff [16'h07_79] = 8'h0A;
    buff [16'h07_7a] = 8'hF0;
    buff [16'h07_7b] = 8'h78;
    buff [16'h07_7c] = 8'h80;
    buff [16'h07_7d] = 8'h18;
    buff [16'h07_7e] = 8'h76;
    buff [16'h07_7f] = 8'h00;
    buff [16'h07_80] = 8'hE8;
    buff [16'h07_81] = 8'h70;
    buff [16'h07_82] = 8'hFA;
    buff [16'h07_83] = 8'h75;
    buff [16'h07_84] = 8'hD0;
    buff [16'h07_85] = 8'h00;
    buff [16'h07_86] = 8'h74;
    buff [16'h07_87] = 8'h90;
    buff [16'h07_88] = 8'h78;
    buff [16'h07_89] = 8'h09;
    buff [16'h07_8a] = 8'h48;
    buff [16'h07_8b] = 8'h94;
    buff [16'h07_8c] = 8'h99;
    buff [16'h07_8d] = 8'h60;
    buff [16'h07_8e] = 8'h06;
    buff [16'h07_8f] = 8'h75;
    buff [16'h07_90] = 8'h90;
    buff [16'h07_91] = 8'h4E;
    buff [16'h07_92] = 8'h02;
    buff [16'h07_93] = 8'h0A;
    buff [16'h07_94] = 8'hF0;
    buff [16'h07_95] = 8'h78;
    buff [16'h07_96] = 8'h80;
    buff [16'h07_97] = 8'h18;
    buff [16'h07_98] = 8'h76;
    buff [16'h07_99] = 8'h00;
    buff [16'h07_9a] = 8'hE8;
    buff [16'h07_9b] = 8'h70;
    buff [16'h07_9c] = 8'hFA;
    buff [16'h07_9d] = 8'h75;
    buff [16'h07_9e] = 8'hD0;
    buff [16'h07_9f] = 8'h00;
    buff [16'h07_a0] = 8'h74;
    buff [16'h07_a1] = 8'h09;
    buff [16'h07_a2] = 8'h75;
    buff [16'h07_a3] = 8'h7F;
    buff [16'h07_a4] = 8'h90;
    buff [16'h07_a5] = 8'h45;
    buff [16'h07_a6] = 8'h7F;
    buff [16'h07_a7] = 8'h94;
    buff [16'h07_a8] = 8'h99;
    buff [16'h07_a9] = 8'h60;
    buff [16'h07_aa] = 8'h06;
    buff [16'h07_ab] = 8'h75;
    buff [16'h07_ac] = 8'h90;
    buff [16'h07_ad] = 8'h4F;
    buff [16'h07_ae] = 8'h02;
    buff [16'h07_af] = 8'h0A;
    buff [16'h07_b0] = 8'hF0;
    buff [16'h07_b1] = 8'h78;
    buff [16'h07_b2] = 8'h80;
    buff [16'h07_b3] = 8'h18;
    buff [16'h07_b4] = 8'h76;
    buff [16'h07_b5] = 8'h00;
    buff [16'h07_b6] = 8'hE8;
    buff [16'h07_b7] = 8'h70;
    buff [16'h07_b8] = 8'hFA;
    buff [16'h07_b9] = 8'h75;
    buff [16'h07_ba] = 8'hD0;
    buff [16'h07_bb] = 8'h00;
    buff [16'h07_bc] = 8'h74;
    buff [16'h07_bd] = 8'h90;
    buff [16'h07_be] = 8'h78;
    buff [16'h07_bf] = 8'h7F;
    buff [16'h07_c0] = 8'h75;
    buff [16'h07_c1] = 8'h7F;
    buff [16'h07_c2] = 8'h06;
    buff [16'h07_c3] = 8'h46;
    buff [16'h07_c4] = 8'h94;
    buff [16'h07_c5] = 8'h96;
    buff [16'h07_c6] = 8'h60;
    buff [16'h07_c7] = 8'h06;
    buff [16'h07_c8] = 8'h75;
    buff [16'h07_c9] = 8'h90;
    buff [16'h07_ca] = 8'h50;
    buff [16'h07_cb] = 8'h02;
    buff [16'h07_cc] = 8'h0A;
    buff [16'h07_cd] = 8'hF0;
    buff [16'h07_ce] = 8'h78;
    buff [16'h07_cf] = 8'h80;
    buff [16'h07_d0] = 8'h18;
    buff [16'h07_d1] = 8'h76;
    buff [16'h07_d2] = 8'h00;
    buff [16'h07_d3] = 8'hE8;
    buff [16'h07_d4] = 8'h70;
    buff [16'h07_d5] = 8'hFA;
    buff [16'h07_d6] = 8'h75;
    buff [16'h07_d7] = 8'hD0;
    buff [16'h07_d8] = 8'h00;
    buff [16'h07_d9] = 8'h74;
    buff [16'h07_da] = 8'h11;
    buff [16'h07_db] = 8'h44;
    buff [16'h07_dc] = 8'h22;
    buff [16'h07_dd] = 8'h94;
    buff [16'h07_de] = 8'h33;
    buff [16'h07_df] = 8'h60;
    buff [16'h07_e0] = 8'h06;
    buff [16'h07_e1] = 8'h75;
    buff [16'h07_e2] = 8'h90;
    buff [16'h07_e3] = 8'h51;
    buff [16'h07_e4] = 8'h02;
    buff [16'h07_e5] = 8'h0A;
    buff [16'h07_e6] = 8'hF0;
    buff [16'h07_e7] = 8'h78;
    buff [16'h07_e8] = 8'h80;
    buff [16'h07_e9] = 8'h18;
    buff [16'h07_ea] = 8'h76;
    buff [16'h07_eb] = 8'h00;
    buff [16'h07_ec] = 8'hE8;
    buff [16'h07_ed] = 8'h70;
    buff [16'h07_ee] = 8'hFA;
    buff [16'h07_ef] = 8'h75;
    buff [16'h07_f0] = 8'hD0;
    buff [16'h07_f1] = 8'h00;
    buff [16'h07_f2] = 8'h74;
    buff [16'h07_f3] = 8'h90;
    buff [16'h07_f4] = 8'h75;
    buff [16'h07_f5] = 8'h7F;
    buff [16'h07_f6] = 8'h09;
    buff [16'h07_f7] = 8'h42;
    buff [16'h07_f8] = 8'h7F;
    buff [16'h07_f9] = 8'hE4;
    buff [16'h07_fa] = 8'hE5;
    buff [16'h07_fb] = 8'h7F;
    buff [16'h07_fc] = 8'h94;
    buff [16'h07_fd] = 8'h99;
    buff [16'h07_fe] = 8'h60;
    buff [16'h07_ff] = 8'h06;
    buff [16'h08_00] = 8'h75;
    buff [16'h08_01] = 8'h90;
    buff [16'h08_02] = 8'h52;
    buff [16'h08_03] = 8'h02;
    buff [16'h08_04] = 8'h0A;
    buff [16'h08_05] = 8'hF0;
    buff [16'h08_06] = 8'h78;
    buff [16'h08_07] = 8'h80;
    buff [16'h08_08] = 8'h18;
    buff [16'h08_09] = 8'h76;
    buff [16'h08_0a] = 8'h00;
    buff [16'h08_0b] = 8'hE8;
    buff [16'h08_0c] = 8'h70;
    buff [16'h08_0d] = 8'hFA;
    buff [16'h08_0e] = 8'h75;
    buff [16'h08_0f] = 8'hD0;
    buff [16'h08_10] = 8'h00;
    buff [16'h08_11] = 8'h75;
    buff [16'h08_12] = 8'h7F;
    buff [16'h08_13] = 8'h90;
    buff [16'h08_14] = 8'h43;
    buff [16'h08_15] = 8'h7F;
    buff [16'h08_16] = 8'h09;
    buff [16'h08_17] = 8'hE5;
    buff [16'h08_18] = 8'h7F;
    buff [16'h08_19] = 8'h94;
    buff [16'h08_1a] = 8'h99;
    buff [16'h08_1b] = 8'h60;
    buff [16'h08_1c] = 8'h06;
    buff [16'h08_1d] = 8'h75;
    buff [16'h08_1e] = 8'h90;
    buff [16'h08_1f] = 8'h53;
    buff [16'h08_20] = 8'h02;
    buff [16'h08_21] = 8'h0A;
    buff [16'h08_22] = 8'hF0;
    buff [16'h08_23] = 8'h78;
    buff [16'h08_24] = 8'h80;
    buff [16'h08_25] = 8'h18;
    buff [16'h08_26] = 8'h76;
    buff [16'h08_27] = 8'h00;
    buff [16'h08_28] = 8'hE8;
    buff [16'h08_29] = 8'h70;
    buff [16'h08_2a] = 8'hFA;
    buff [16'h08_2b] = 8'h75;
    buff [16'h08_2c] = 8'hD0;
    buff [16'h08_2d] = 8'h00;
    buff [16'h08_2e] = 8'h72;
    buff [16'h08_2f] = 8'hE0;
    buff [16'h08_30] = 8'h40;
    buff [16'h08_31] = 8'h0A;
    buff [16'h08_32] = 8'h74;
    buff [16'h08_33] = 8'h01;
    buff [16'h08_34] = 8'h72;
    buff [16'h08_35] = 8'hE0;
    buff [16'h08_36] = 8'h50;
    buff [16'h08_37] = 8'h04;
    buff [16'h08_38] = 8'h72;
    buff [16'h08_39] = 8'hE1;
    buff [16'h08_3a] = 8'h40;
    buff [16'h08_3b] = 8'h06;
    buff [16'h08_3c] = 8'h75;
    buff [16'h08_3d] = 8'h90;
    buff [16'h08_3e] = 8'h54;
    buff [16'h08_3f] = 8'h02;
    buff [16'h08_40] = 8'h0A;
    buff [16'h08_41] = 8'hF0;
    buff [16'h08_42] = 8'h78;
    buff [16'h08_43] = 8'h80;
    buff [16'h08_44] = 8'h18;
    buff [16'h08_45] = 8'h76;
    buff [16'h08_46] = 8'h00;
    buff [16'h08_47] = 8'hE8;
    buff [16'h08_48] = 8'h70;
    buff [16'h08_49] = 8'hFA;
    buff [16'h08_4a] = 8'h75;
    buff [16'h08_4b] = 8'hD0;
    buff [16'h08_4c] = 8'h00;
    buff [16'h08_4d] = 8'h74;
    buff [16'h08_4e] = 8'h01;
    buff [16'h08_4f] = 8'hA0;
    buff [16'h08_50] = 8'hE0;
    buff [16'h08_51] = 8'h40;
    buff [16'h08_52] = 8'h08;
    buff [16'h08_53] = 8'hA0;
    buff [16'h08_54] = 8'hE1;
    buff [16'h08_55] = 8'h50;
    buff [16'h08_56] = 8'h04;
    buff [16'h08_57] = 8'hA0;
    buff [16'h08_58] = 8'hE0;
    buff [16'h08_59] = 8'h40;
    buff [16'h08_5a] = 8'h06;
    buff [16'h08_5b] = 8'h75;
    buff [16'h08_5c] = 8'h90;
    buff [16'h08_5d] = 8'h55;
    buff [16'h08_5e] = 8'h02;
    buff [16'h08_5f] = 8'h0A;
    buff [16'h08_60] = 8'hF0;
    buff [16'h08_61] = 8'h78;
    buff [16'h08_62] = 8'h80;
    buff [16'h08_63] = 8'h18;
    buff [16'h08_64] = 8'h76;
    buff [16'h08_65] = 8'h00;
    buff [16'h08_66] = 8'hE8;
    buff [16'h08_67] = 8'h70;
    buff [16'h08_68] = 8'hFA;
    buff [16'h08_69] = 8'h75;
    buff [16'h08_6a] = 8'hD0;
    buff [16'h08_6b] = 8'h00;
    buff [16'h08_6c] = 8'h90;
    buff [16'h08_6d] = 8'h01;
    buff [16'h08_6e] = 8'h23;
    buff [16'h08_6f] = 8'h75;
    buff [16'h08_70] = 8'h7F;
    buff [16'h08_71] = 8'h08;
    buff [16'h08_72] = 8'hC0;
    buff [16'h08_73] = 8'h82;
    buff [16'h08_74] = 8'hC0;
    buff [16'h08_75] = 8'h83;
    buff [16'h08_76] = 8'hC0;
    buff [16'h08_77] = 8'h7F;
    buff [16'h08_78] = 8'hE5;
    buff [16'h08_79] = 8'h08;
    buff [16'h08_7a] = 8'h94;
    buff [16'h08_7b] = 8'h23;
    buff [16'h08_7c] = 8'h70;
    buff [16'h08_7d] = 8'h0C;
    buff [16'h08_7e] = 8'hE5;
    buff [16'h08_7f] = 8'h09;
    buff [16'h08_80] = 8'h94;
    buff [16'h08_81] = 8'h01;
    buff [16'h08_82] = 8'h70;
    buff [16'h08_83] = 8'h06;
    buff [16'h08_84] = 8'hE5;
    buff [16'h08_85] = 8'h0A;
    buff [16'h08_86] = 8'h94;
    buff [16'h08_87] = 8'h08;
    buff [16'h08_88] = 8'h60;
    buff [16'h08_89] = 8'h06;
    buff [16'h08_8a] = 8'h75;
    buff [16'h08_8b] = 8'h90;
    buff [16'h08_8c] = 8'h57;
    buff [16'h08_8d] = 8'h02;
    buff [16'h08_8e] = 8'h0A;
    buff [16'h08_8f] = 8'hF0;
    buff [16'h08_90] = 8'hD0;
    buff [16'h08_91] = 8'h81;
    buff [16'h08_92] = 8'hD0;
    buff [16'h08_93] = 8'h64;
    buff [16'h08_94] = 8'hE5;
    buff [16'h08_95] = 8'h64;
    buff [16'h08_96] = 8'h94;
    buff [16'h08_97] = 8'h23;
    buff [16'h08_98] = 8'h60;
    buff [16'h08_99] = 8'h06;
    buff [16'h08_9a] = 8'h75;
    buff [16'h08_9b] = 8'h90;
    buff [16'h08_9c] = 8'h56;
    buff [16'h08_9d] = 8'h02;
    buff [16'h08_9e] = 8'h0A;
    buff [16'h08_9f] = 8'hF0;
    buff [16'h08_a0] = 8'h78;
    buff [16'h08_a1] = 8'h80;
    buff [16'h08_a2] = 8'h18;
    buff [16'h08_a3] = 8'h76;
    buff [16'h08_a4] = 8'h00;
    buff [16'h08_a5] = 8'hE8;
    buff [16'h08_a6] = 8'h70;
    buff [16'h08_a7] = 8'hFA;
    buff [16'h08_a8] = 8'h75;
    buff [16'h08_a9] = 8'hD0;
    buff [16'h08_aa] = 8'h00;
    buff [16'h08_ab] = 8'h74;
    buff [16'h08_ac] = 8'h81;
    buff [16'h08_ad] = 8'h23;
    buff [16'h08_ae] = 8'h94;
    buff [16'h08_af] = 8'h03;
    buff [16'h08_b0] = 8'h60;
    buff [16'h08_b1] = 8'h06;
    buff [16'h08_b2] = 8'h75;
    buff [16'h08_b3] = 8'h90;
    buff [16'h08_b4] = 8'h5A;
    buff [16'h08_b5] = 8'h02;
    buff [16'h08_b6] = 8'h0A;
    buff [16'h08_b7] = 8'hF0;
    buff [16'h08_b8] = 8'h78;
    buff [16'h08_b9] = 8'h80;
    buff [16'h08_ba] = 8'h18;
    buff [16'h08_bb] = 8'h76;
    buff [16'h08_bc] = 8'h00;
    buff [16'h08_bd] = 8'hE8;
    buff [16'h08_be] = 8'h70;
    buff [16'h08_bf] = 8'hFA;
    buff [16'h08_c0] = 8'h75;
    buff [16'h08_c1] = 8'hD0;
    buff [16'h08_c2] = 8'h00;
    buff [16'h08_c3] = 8'h74;
    buff [16'h08_c4] = 8'h81;
    buff [16'h08_c5] = 8'h33;
    buff [16'h08_c6] = 8'h94;
    buff [16'h08_c7] = 8'h01;
    buff [16'h08_c8] = 8'h60;
    buff [16'h08_c9] = 8'h06;
    buff [16'h08_ca] = 8'h75;
    buff [16'h08_cb] = 8'h90;
    buff [16'h08_cc] = 8'h5B;
    buff [16'h08_cd] = 8'h02;
    buff [16'h08_ce] = 8'h0A;
    buff [16'h08_cf] = 8'hF0;
    buff [16'h08_d0] = 8'h78;
    buff [16'h08_d1] = 8'h80;
    buff [16'h08_d2] = 8'h18;
    buff [16'h08_d3] = 8'h76;
    buff [16'h08_d4] = 8'h00;
    buff [16'h08_d5] = 8'hE8;
    buff [16'h08_d6] = 8'h70;
    buff [16'h08_d7] = 8'hFA;
    buff [16'h08_d8] = 8'h75;
    buff [16'h08_d9] = 8'hD0;
    buff [16'h08_da] = 8'h00;
    buff [16'h08_db] = 8'h74;
    buff [16'h08_dc] = 8'h81;
    buff [16'h08_dd] = 8'h03;
    buff [16'h08_de] = 8'h94;
    buff [16'h08_df] = 8'hC0;
    buff [16'h08_e0] = 8'h60;
    buff [16'h08_e1] = 8'h06;
    buff [16'h08_e2] = 8'h75;
    buff [16'h08_e3] = 8'h90;
    buff [16'h08_e4] = 8'h5C;
    buff [16'h08_e5] = 8'h02;
    buff [16'h08_e6] = 8'h0A;
    buff [16'h08_e7] = 8'hF0;
    buff [16'h08_e8] = 8'h78;
    buff [16'h08_e9] = 8'h80;
    buff [16'h08_ea] = 8'h18;
    buff [16'h08_eb] = 8'h76;
    buff [16'h08_ec] = 8'h00;
    buff [16'h08_ed] = 8'hE8;
    buff [16'h08_ee] = 8'h70;
    buff [16'h08_ef] = 8'hFA;
    buff [16'h08_f0] = 8'h75;
    buff [16'h08_f1] = 8'hD0;
    buff [16'h08_f2] = 8'h00;
    buff [16'h08_f3] = 8'h74;
    buff [16'h08_f4] = 8'h03;
    buff [16'h08_f5] = 8'h13;
    buff [16'h08_f6] = 8'h94;
    buff [16'h08_f7] = 8'h00;
    buff [16'h08_f8] = 8'h60;
    buff [16'h08_f9] = 8'h06;
    buff [16'h08_fa] = 8'h75;
    buff [16'h08_fb] = 8'h90;
    buff [16'h08_fc] = 8'h5D;
    buff [16'h08_fd] = 8'h02;
    buff [16'h08_fe] = 8'h0A;
    buff [16'h08_ff] = 8'hF0;
    buff [16'h09_00] = 8'h78;
    buff [16'h09_01] = 8'h80;
    buff [16'h09_02] = 8'h18;
    buff [16'h09_03] = 8'h76;
    buff [16'h09_04] = 8'h00;
    buff [16'h09_05] = 8'hE8;
    buff [16'h09_06] = 8'h70;
    buff [16'h09_07] = 8'hFA;
    buff [16'h09_08] = 8'h75;
    buff [16'h09_09] = 8'hD0;
    buff [16'h09_0a] = 8'h00;
    buff [16'h09_0b] = 8'hD3;
    buff [16'h09_0c] = 8'h74;
    buff [16'h09_0d] = 8'h01;
    buff [16'h09_0e] = 8'h94;
    buff [16'h09_0f] = 8'h00;
    buff [16'h09_10] = 8'h60;
    buff [16'h09_11] = 8'h06;
    buff [16'h09_12] = 8'h75;
    buff [16'h09_13] = 8'h90;
    buff [16'h09_14] = 8'h5E;
    buff [16'h09_15] = 8'h02;
    buff [16'h09_16] = 8'h0A;
    buff [16'h09_17] = 8'hF0;
    buff [16'h09_18] = 8'h78;
    buff [16'h09_19] = 8'h80;
    buff [16'h09_1a] = 8'h18;
    buff [16'h09_1b] = 8'h76;
    buff [16'h09_1c] = 8'h00;
    buff [16'h09_1d] = 8'hE8;
    buff [16'h09_1e] = 8'h70;
    buff [16'h09_1f] = 8'hFA;
    buff [16'h09_20] = 8'h75;
    buff [16'h09_21] = 8'hD0;
    buff [16'h09_22] = 8'h00;
    buff [16'h09_23] = 8'hD2;
    buff [16'h09_24] = 8'hE7;
    buff [16'h09_25] = 8'h94;
    buff [16'h09_26] = 8'h80;
    buff [16'h09_27] = 8'h60;
    buff [16'h09_28] = 8'h06;
    buff [16'h09_29] = 8'h75;
    buff [16'h09_2a] = 8'h90;
    buff [16'h09_2b] = 8'h5F;
    buff [16'h09_2c] = 8'h02;
    buff [16'h09_2d] = 8'h0A;
    buff [16'h09_2e] = 8'hF0;
    buff [16'h09_2f] = 8'h78;
    buff [16'h09_30] = 8'h80;
    buff [16'h09_31] = 8'h18;
    buff [16'h09_32] = 8'h76;
    buff [16'h09_33] = 8'h00;
    buff [16'h09_34] = 8'hE8;
    buff [16'h09_35] = 8'h70;
    buff [16'h09_36] = 8'hFA;
    buff [16'h09_37] = 8'h75;
    buff [16'h09_38] = 8'hD0;
    buff [16'h09_39] = 8'h00;
    buff [16'h09_3a] = 8'h80;
    buff [16'h09_3b] = 8'h06;
    buff [16'h09_3c] = 8'h75;
    buff [16'h09_3d] = 8'h90;
    buff [16'h09_3e] = 8'h60;
    buff [16'h09_3f] = 8'h02;
    buff [16'h09_40] = 8'h0A;
    buff [16'h09_41] = 8'hF0;
    buff [16'h09_42] = 8'h78;
    buff [16'h09_43] = 8'h80;
    buff [16'h09_44] = 8'h18;
    buff [16'h09_45] = 8'h76;
    buff [16'h09_46] = 8'h00;
    buff [16'h09_47] = 8'hE8;
    buff [16'h09_48] = 8'h70;
    buff [16'h09_49] = 8'hFA;
    buff [16'h09_4a] = 8'h75;
    buff [16'h09_4b] = 8'hD0;
    buff [16'h09_4c] = 8'h00;
    buff [16'h09_4d] = 8'h74;
    buff [16'h09_4e] = 8'h0A;
    buff [16'h09_4f] = 8'h78;
    buff [16'h09_50] = 8'h0A;
    buff [16'h09_51] = 8'h98;
    buff [16'h09_52] = 8'h60;
    buff [16'h09_53] = 8'h06;
    buff [16'h09_54] = 8'h75;
    buff [16'h09_55] = 8'h90;
    buff [16'h09_56] = 8'h61;
    buff [16'h09_57] = 8'h02;
    buff [16'h09_58] = 8'h0A;
    buff [16'h09_59] = 8'hF0;
    buff [16'h09_5a] = 8'h78;
    buff [16'h09_5b] = 8'h80;
    buff [16'h09_5c] = 8'h18;
    buff [16'h09_5d] = 8'h76;
    buff [16'h09_5e] = 8'h00;
    buff [16'h09_5f] = 8'hE8;
    buff [16'h09_60] = 8'h70;
    buff [16'h09_61] = 8'hFA;
    buff [16'h09_62] = 8'h75;
    buff [16'h09_63] = 8'hD0;
    buff [16'h09_64] = 8'h00;
    buff [16'h09_65] = 8'h74;
    buff [16'h09_66] = 8'h0A;
    buff [16'h09_67] = 8'h75;
    buff [16'h09_68] = 8'h7F;
    buff [16'h09_69] = 8'h0A;
    buff [16'h09_6a] = 8'h95;
    buff [16'h09_6b] = 8'h7F;
    buff [16'h09_6c] = 8'h60;
    buff [16'h09_6d] = 8'h06;
    buff [16'h09_6e] = 8'h75;
    buff [16'h09_6f] = 8'h90;
    buff [16'h09_70] = 8'h62;
    buff [16'h09_71] = 8'h02;
    buff [16'h09_72] = 8'h0A;
    buff [16'h09_73] = 8'hF0;
    buff [16'h09_74] = 8'h78;
    buff [16'h09_75] = 8'h80;
    buff [16'h09_76] = 8'h18;
    buff [16'h09_77] = 8'h76;
    buff [16'h09_78] = 8'h00;
    buff [16'h09_79] = 8'hE8;
    buff [16'h09_7a] = 8'h70;
    buff [16'h09_7b] = 8'hFA;
    buff [16'h09_7c] = 8'h75;
    buff [16'h09_7d] = 8'hD0;
    buff [16'h09_7e] = 8'h00;
    buff [16'h09_7f] = 8'h74;
    buff [16'h09_80] = 8'h0A;
    buff [16'h09_81] = 8'h78;
    buff [16'h09_82] = 8'h7F;
    buff [16'h09_83] = 8'h75;
    buff [16'h09_84] = 8'h7F;
    buff [16'h09_85] = 8'h0A;
    buff [16'h09_86] = 8'h96;
    buff [16'h09_87] = 8'h60;
    buff [16'h09_88] = 8'h06;
    buff [16'h09_89] = 8'h75;
    buff [16'h09_8a] = 8'h90;
    buff [16'h09_8b] = 8'h63;
    buff [16'h09_8c] = 8'h02;
    buff [16'h09_8d] = 8'h0A;
    buff [16'h09_8e] = 8'hF0;
    buff [16'h09_8f] = 8'h78;
    buff [16'h09_90] = 8'h80;
    buff [16'h09_91] = 8'h18;
    buff [16'h09_92] = 8'h76;
    buff [16'h09_93] = 8'h00;
    buff [16'h09_94] = 8'hE8;
    buff [16'h09_95] = 8'h70;
    buff [16'h09_96] = 8'hFA;
    buff [16'h09_97] = 8'h75;
    buff [16'h09_98] = 8'hD0;
    buff [16'h09_99] = 8'h00;
    buff [16'h09_9a] = 8'h74;
    buff [16'h09_9b] = 8'h0A;
    buff [16'h09_9c] = 8'h94;
    buff [16'h09_9d] = 8'h0A;
    buff [16'h09_9e] = 8'h60;
    buff [16'h09_9f] = 8'h06;
    buff [16'h09_a0] = 8'h75;
    buff [16'h09_a1] = 8'h90;
    buff [16'h09_a2] = 8'h64;
    buff [16'h09_a3] = 8'h02;
    buff [16'h09_a4] = 8'h0A;
    buff [16'h09_a5] = 8'hF0;
    buff [16'h09_a6] = 8'h78;
    buff [16'h09_a7] = 8'h80;
    buff [16'h09_a8] = 8'h18;
    buff [16'h09_a9] = 8'h76;
    buff [16'h09_aa] = 8'h00;
    buff [16'h09_ab] = 8'hE8;
    buff [16'h09_ac] = 8'h70;
    buff [16'h09_ad] = 8'hFA;
    buff [16'h09_ae] = 8'h75;
    buff [16'h09_af] = 8'hD0;
    buff [16'h09_b0] = 8'h00;
    buff [16'h09_b1] = 8'h74;
    buff [16'h09_b2] = 8'h23;
    buff [16'h09_b3] = 8'hC4;
    buff [16'h09_b4] = 8'h94;
    buff [16'h09_b5] = 8'h32;
    buff [16'h09_b6] = 8'h60;
    buff [16'h09_b7] = 8'h06;
    buff [16'h09_b8] = 8'h75;
    buff [16'h09_b9] = 8'h90;
    buff [16'h09_ba] = 8'h65;
    buff [16'h09_bb] = 8'h02;
    buff [16'h09_bc] = 8'h0A;
    buff [16'h09_bd] = 8'hF0;
    buff [16'h09_be] = 8'h78;
    buff [16'h09_bf] = 8'h80;
    buff [16'h09_c0] = 8'h18;
    buff [16'h09_c1] = 8'h76;
    buff [16'h09_c2] = 8'h00;
    buff [16'h09_c3] = 8'hE8;
    buff [16'h09_c4] = 8'h70;
    buff [16'h09_c5] = 8'hFA;
    buff [16'h09_c6] = 8'h75;
    buff [16'h09_c7] = 8'hD0;
    buff [16'h09_c8] = 8'h00;
    buff [16'h09_c9] = 8'h74;
    buff [16'h09_ca] = 8'h0A;
    buff [16'h09_cb] = 8'h78;
    buff [16'h09_cc] = 8'h63;
    buff [16'h09_cd] = 8'hC8;
    buff [16'h09_ce] = 8'h94;
    buff [16'h09_cf] = 8'h63;
    buff [16'h09_d0] = 8'h70;
    buff [16'h09_d1] = 8'h05;
    buff [16'h09_d2] = 8'hE8;
    buff [16'h09_d3] = 8'h94;
    buff [16'h09_d4] = 8'h0A;
    buff [16'h09_d5] = 8'h60;
    buff [16'h09_d6] = 8'h06;
    buff [16'h09_d7] = 8'h75;
    buff [16'h09_d8] = 8'h90;
    buff [16'h09_d9] = 8'h66;
    buff [16'h09_da] = 8'h02;
    buff [16'h09_db] = 8'h0A;
    buff [16'h09_dc] = 8'hF0;
    buff [16'h09_dd] = 8'h78;
    buff [16'h09_de] = 8'h80;
    buff [16'h09_df] = 8'h18;
    buff [16'h09_e0] = 8'h76;
    buff [16'h09_e1] = 8'h00;
    buff [16'h09_e2] = 8'hE8;
    buff [16'h09_e3] = 8'h70;
    buff [16'h09_e4] = 8'hFA;
    buff [16'h09_e5] = 8'h75;
    buff [16'h09_e6] = 8'hD0;
    buff [16'h09_e7] = 8'h00;
    buff [16'h09_e8] = 8'h74;
    buff [16'h09_e9] = 8'h0A;
    buff [16'h09_ea] = 8'h75;
    buff [16'h09_eb] = 8'h7F;
    buff [16'h09_ec] = 8'h63;
    buff [16'h09_ed] = 8'hC5;
    buff [16'h09_ee] = 8'h7F;
    buff [16'h09_ef] = 8'h94;
    buff [16'h09_f0] = 8'h63;
    buff [16'h09_f1] = 8'h70;
    buff [16'h09_f2] = 8'h06;
    buff [16'h09_f3] = 8'hE5;
    buff [16'h09_f4] = 8'h7F;
    buff [16'h09_f5] = 8'h94;
    buff [16'h09_f6] = 8'h0A;
    buff [16'h09_f7] = 8'h60;
    buff [16'h09_f8] = 8'h06;
    buff [16'h09_f9] = 8'h75;
    buff [16'h09_fa] = 8'h90;
    buff [16'h09_fb] = 8'h67;
    buff [16'h09_fc] = 8'h02;
    buff [16'h09_fd] = 8'h0A;
    buff [16'h09_fe] = 8'hF0;
    buff [16'h09_ff] = 8'h78;
    buff [16'h0a_00] = 8'h80;
    buff [16'h0a_01] = 8'h18;
    buff [16'h0a_02] = 8'h76;
    buff [16'h0a_03] = 8'h00;
    buff [16'h0a_04] = 8'hE8;
    buff [16'h0a_05] = 8'h70;
    buff [16'h0a_06] = 8'hFA;
    buff [16'h0a_07] = 8'h75;
    buff [16'h0a_08] = 8'hD0;
    buff [16'h0a_09] = 8'h00;
    buff [16'h0a_0a] = 8'h74;
    buff [16'h0a_0b] = 8'h0A;
    buff [16'h0a_0c] = 8'h78;
    buff [16'h0a_0d] = 8'h7F;
    buff [16'h0a_0e] = 8'h75;
    buff [16'h0a_0f] = 8'h7F;
    buff [16'h0a_10] = 8'h63;
    buff [16'h0a_11] = 8'hC6;
    buff [16'h0a_12] = 8'h94;
    buff [16'h0a_13] = 8'h63;
    buff [16'h0a_14] = 8'h70;
    buff [16'h0a_15] = 8'h06;
    buff [16'h0a_16] = 8'hE5;
    buff [16'h0a_17] = 8'h7F;
    buff [16'h0a_18] = 8'h94;
    buff [16'h0a_19] = 8'h0A;
    buff [16'h0a_1a] = 8'h60;
    buff [16'h0a_1b] = 8'h06;
    buff [16'h0a_1c] = 8'h75;
    buff [16'h0a_1d] = 8'h90;
    buff [16'h0a_1e] = 8'h68;
    buff [16'h0a_1f] = 8'h02;
    buff [16'h0a_20] = 8'h0A;
    buff [16'h0a_21] = 8'hF0;
    buff [16'h0a_22] = 8'h78;
    buff [16'h0a_23] = 8'h80;
    buff [16'h0a_24] = 8'h18;
    buff [16'h0a_25] = 8'h76;
    buff [16'h0a_26] = 8'h00;
    buff [16'h0a_27] = 8'hE8;
    buff [16'h0a_28] = 8'h70;
    buff [16'h0a_29] = 8'hFA;
    buff [16'h0a_2a] = 8'h75;
    buff [16'h0a_2b] = 8'hD0;
    buff [16'h0a_2c] = 8'h00;
    buff [16'h0a_2d] = 8'h74;
    buff [16'h0a_2e] = 8'h44;
    buff [16'h0a_2f] = 8'h78;
    buff [16'h0a_30] = 8'h7F;
    buff [16'h0a_31] = 8'h75;
    buff [16'h0a_32] = 8'h7F;
    buff [16'h0a_33] = 8'h55;
    buff [16'h0a_34] = 8'hD6;
    buff [16'h0a_35] = 8'h94;
    buff [16'h0a_36] = 8'h45;
    buff [16'h0a_37] = 8'h70;
    buff [16'h0a_38] = 8'h06;
    buff [16'h0a_39] = 8'hE5;
    buff [16'h0a_3a] = 8'h7F;
    buff [16'h0a_3b] = 8'h94;
    buff [16'h0a_3c] = 8'h54;
    buff [16'h0a_3d] = 8'h60;
    buff [16'h0a_3e] = 8'h06;
    buff [16'h0a_3f] = 8'h75;
    buff [16'h0a_40] = 8'h90;
    buff [16'h0a_41] = 8'h69;
    buff [16'h0a_42] = 8'h02;
    buff [16'h0a_43] = 8'h0A;
    buff [16'h0a_44] = 8'hF0;
    buff [16'h0a_45] = 8'h78;
    buff [16'h0a_46] = 8'h80;
    buff [16'h0a_47] = 8'h18;
    buff [16'h0a_48] = 8'h76;
    buff [16'h0a_49] = 8'h00;
    buff [16'h0a_4a] = 8'hE8;
    buff [16'h0a_4b] = 8'h70;
    buff [16'h0a_4c] = 8'hFA;
    buff [16'h0a_4d] = 8'h75;
    buff [16'h0a_4e] = 8'hD0;
    buff [16'h0a_4f] = 8'h00;
    buff [16'h0a_50] = 8'h74;
    buff [16'h0a_51] = 8'h35;
    buff [16'h0a_52] = 8'h78;
    buff [16'h0a_53] = 8'h53;
    buff [16'h0a_54] = 8'h68;
    buff [16'h0a_55] = 8'h94;
    buff [16'h0a_56] = 8'h66;
    buff [16'h0a_57] = 8'h60;
    buff [16'h0a_58] = 8'h06;
    buff [16'h0a_59] = 8'h75;
    buff [16'h0a_5a] = 8'h90;
    buff [16'h0a_5b] = 8'h6A;
    buff [16'h0a_5c] = 8'h02;
    buff [16'h0a_5d] = 8'h0A;
    buff [16'h0a_5e] = 8'hF0;
    buff [16'h0a_5f] = 8'h78;
    buff [16'h0a_60] = 8'h80;
    buff [16'h0a_61] = 8'h18;
    buff [16'h0a_62] = 8'h76;
    buff [16'h0a_63] = 8'h00;
    buff [16'h0a_64] = 8'hE8;
    buff [16'h0a_65] = 8'h70;
    buff [16'h0a_66] = 8'hFA;
    buff [16'h0a_67] = 8'h75;
    buff [16'h0a_68] = 8'hD0;
    buff [16'h0a_69] = 8'h00;
    buff [16'h0a_6a] = 8'h74;
    buff [16'h0a_6b] = 8'h53;
    buff [16'h0a_6c] = 8'h75;
    buff [16'h0a_6d] = 8'h7F;
    buff [16'h0a_6e] = 8'h35;
    buff [16'h0a_6f] = 8'h65;
    buff [16'h0a_70] = 8'h7F;
    buff [16'h0a_71] = 8'h94;
    buff [16'h0a_72] = 8'h66;
    buff [16'h0a_73] = 8'h60;
    buff [16'h0a_74] = 8'h06;
    buff [16'h0a_75] = 8'h75;
    buff [16'h0a_76] = 8'h90;
    buff [16'h0a_77] = 8'h6B;
    buff [16'h0a_78] = 8'h02;
    buff [16'h0a_79] = 8'h0A;
    buff [16'h0a_7a] = 8'hF0;
    buff [16'h0a_7b] = 8'h78;
    buff [16'h0a_7c] = 8'h80;
    buff [16'h0a_7d] = 8'h18;
    buff [16'h0a_7e] = 8'h76;
    buff [16'h0a_7f] = 8'h00;
    buff [16'h0a_80] = 8'hE8;
    buff [16'h0a_81] = 8'h70;
    buff [16'h0a_82] = 8'hFA;
    buff [16'h0a_83] = 8'h75;
    buff [16'h0a_84] = 8'hD0;
    buff [16'h0a_85] = 8'h00;
    buff [16'h0a_86] = 8'h74;
    buff [16'h0a_87] = 8'h35;
    buff [16'h0a_88] = 8'h78;
    buff [16'h0a_89] = 8'h7F;
    buff [16'h0a_8a] = 8'h75;
    buff [16'h0a_8b] = 8'h7F;
    buff [16'h0a_8c] = 8'h53;
    buff [16'h0a_8d] = 8'h66;
    buff [16'h0a_8e] = 8'h94;
    buff [16'h0a_8f] = 8'h66;
    buff [16'h0a_90] = 8'h60;
    buff [16'h0a_91] = 8'h06;
    buff [16'h0a_92] = 8'h75;
    buff [16'h0a_93] = 8'h90;
    buff [16'h0a_94] = 8'h6C;
    buff [16'h0a_95] = 8'h02;
    buff [16'h0a_96] = 8'h0A;
    buff [16'h0a_97] = 8'hF0;
    buff [16'h0a_98] = 8'h78;
    buff [16'h0a_99] = 8'h80;
    buff [16'h0a_9a] = 8'h18;
    buff [16'h0a_9b] = 8'h76;
    buff [16'h0a_9c] = 8'h00;
    buff [16'h0a_9d] = 8'hE8;
    buff [16'h0a_9e] = 8'h70;
    buff [16'h0a_9f] = 8'hFA;
    buff [16'h0a_a0] = 8'h75;
    buff [16'h0a_a1] = 8'hD0;
    buff [16'h0a_a2] = 8'h00;
    buff [16'h0a_a3] = 8'h74;
    buff [16'h0a_a4] = 8'h35;
    buff [16'h0a_a5] = 8'h64;
    buff [16'h0a_a6] = 8'h53;
    buff [16'h0a_a7] = 8'h94;
    buff [16'h0a_a8] = 8'h66;
    buff [16'h0a_a9] = 8'h60;
    buff [16'h0a_aa] = 8'h06;
    buff [16'h0a_ab] = 8'h75;
    buff [16'h0a_ac] = 8'h90;
    buff [16'h0a_ad] = 8'h6D;
    buff [16'h0a_ae] = 8'h02;
    buff [16'h0a_af] = 8'h0A;
    buff [16'h0a_b0] = 8'hF0;
    buff [16'h0a_b1] = 8'h78;
    buff [16'h0a_b2] = 8'h80;
    buff [16'h0a_b3] = 8'h18;
    buff [16'h0a_b4] = 8'h76;
    buff [16'h0a_b5] = 8'h00;
    buff [16'h0a_b6] = 8'hE8;
    buff [16'h0a_b7] = 8'h70;
    buff [16'h0a_b8] = 8'hFA;
    buff [16'h0a_b9] = 8'h75;
    buff [16'h0a_ba] = 8'hD0;
    buff [16'h0a_bb] = 8'h00;
    buff [16'h0a_bc] = 8'h74;
    buff [16'h0a_bd] = 8'h35;
    buff [16'h0a_be] = 8'h75;
    buff [16'h0a_bf] = 8'h7F;
    buff [16'h0a_c0] = 8'h53;
    buff [16'h0a_c1] = 8'h62;
    buff [16'h0a_c2] = 8'h7F;
    buff [16'h0a_c3] = 8'hE4;
    buff [16'h0a_c4] = 8'hE5;
    buff [16'h0a_c5] = 8'h7F;
    buff [16'h0a_c6] = 8'h94;
    buff [16'h0a_c7] = 8'h66;
    buff [16'h0a_c8] = 8'h60;
    buff [16'h0a_c9] = 8'h06;
    buff [16'h0a_ca] = 8'h75;
    buff [16'h0a_cb] = 8'h90;
    buff [16'h0a_cc] = 8'h6E;
    buff [16'h0a_cd] = 8'h02;
    buff [16'h0a_ce] = 8'h0A;
    buff [16'h0a_cf] = 8'hF0;
    buff [16'h0a_d0] = 8'h78;
    buff [16'h0a_d1] = 8'h80;
    buff [16'h0a_d2] = 8'h18;
    buff [16'h0a_d3] = 8'h76;
    buff [16'h0a_d4] = 8'h00;
    buff [16'h0a_d5] = 8'hE8;
    buff [16'h0a_d6] = 8'h70;
    buff [16'h0a_d7] = 8'hFA;
    buff [16'h0a_d8] = 8'h75;
    buff [16'h0a_d9] = 8'hD0;
    buff [16'h0a_da] = 8'h00;
    buff [16'h0a_db] = 8'h75;
    buff [16'h0a_dc] = 8'h7F;
    buff [16'h0a_dd] = 8'h35;
    buff [16'h0a_de] = 8'h63;
    buff [16'h0a_df] = 8'h7F;
    buff [16'h0a_e0] = 8'h53;
    buff [16'h0a_e1] = 8'hE5;
    buff [16'h0a_e2] = 8'h7F;
    buff [16'h0a_e3] = 8'h94;
    buff [16'h0a_e4] = 8'h66;
    buff [16'h0a_e5] = 8'h60;
    buff [16'h0a_e6] = 8'h06;
    buff [16'h0a_e7] = 8'h75;
    buff [16'h0a_e8] = 8'h90;
    buff [16'h0a_e9] = 8'h6F;
    buff [16'h0a_ea] = 8'h02;
    buff [16'h0a_eb] = 8'h0A;
    buff [16'h0a_ec] = 8'hF0;
    buff [16'h0a_ed] = 8'h75;
    buff [16'h0a_ee] = 8'h90;
    buff [16'h0a_ef] = 8'h7F;
    buff [16'h0a_f0] = 8'h80;
    buff [16'h0a_f1] = 8'hFE;
    buff [16'h0a_f2] = 8'h22;
end

always @(posedge clk)
begin
  data1 <= #1 buff [addr];
  data2 <= #1 buff [addr+1];
  data3 <= #1 buff [addr+2];
end

endmodule
