-- GR USB 2.0 Device Controller
  constant CFG_GRUSBDC        : integer := CONFIG_GRUSBDC_ENABLE;
  constant CFG_GRUSBDC_AIFACE : integer := CONFIG_GRUSBDC_AIFACE;
  constant CFG_GRUSBDC_UIFACE : integer := CONFIG_GRUSBDC_UIFACE;
  constant CFG_GRUSBDC_DW     : integer := CONFIG_GRUSBDC_DW;
  constant CFG_GRUSBDC_NEPI   : integer := CONFIG_GRUSBDC_NEPI;
  constant CFG_GRUSBDC_NEPO   : integer := CONFIG_GRUSBDC_NEPO;
  constant CFG_GRUSBDC_I0     : integer := CONFIG_GRUSBDC_I0;
  constant CFG_GRUSBDC_I1     : integer := CONFIG_GRUSBDC_I1;
  constant CFG_GRUSBDC_I2     : integer := CONFIG_GRUSBDC_I2;
  constant CFG_GRUSBDC_I3     : integer := CONFIG_GRUSBDC_I3;
  constant CFG_GRUSBDC_I4     : integer := CONFIG_GRUSBDC_I4;
  constant CFG_GRUSBDC_I5     : integer := CONFIG_GRUSBDC_I5;
  constant CFG_GRUSBDC_I6     : integer := CONFIG_GRUSBDC_I6;
  constant CFG_GRUSBDC_I7     : integer := CONFIG_GRUSBDC_I7;
  constant CFG_GRUSBDC_I8     : integer := CONFIG_GRUSBDC_I8;
  constant CFG_GRUSBDC_I9     : integer := CONFIG_GRUSBDC_I9;
  constant CFG_GRUSBDC_I10    : integer := CONFIG_GRUSBDC_I10;
  constant CFG_GRUSBDC_I11    : integer := CONFIG_GRUSBDC_I11;
  constant CFG_GRUSBDC_I12    : integer := CONFIG_GRUSBDC_I12;
  constant CFG_GRUSBDC_I13    : integer := CONFIG_GRUSBDC_I13;
  constant CFG_GRUSBDC_I14    : integer := CONFIG_GRUSBDC_I14;
  constant CFG_GRUSBDC_I15    : integer := CONFIG_GRUSBDC_I15;
  constant CFG_GRUSBDC_O0     : integer := CONFIG_GRUSBDC_O0;
  constant CFG_GRUSBDC_O1     : integer := CONFIG_GRUSBDC_O1;
  constant CFG_GRUSBDC_O2     : integer := CONFIG_GRUSBDC_O2;
  constant CFG_GRUSBDC_O3     : integer := CONFIG_GRUSBDC_O3;
  constant CFG_GRUSBDC_O4     : integer := CONFIG_GRUSBDC_O4;
  constant CFG_GRUSBDC_O5     : integer := CONFIG_GRUSBDC_O5;
  constant CFG_GRUSBDC_O6     : integer := CONFIG_GRUSBDC_O6;
  constant CFG_GRUSBDC_O7     : integer := CONFIG_GRUSBDC_O7;
  constant CFG_GRUSBDC_O8     : integer := CONFIG_GRUSBDC_O8;
  constant CFG_GRUSBDC_O9     : integer := CONFIG_GRUSBDC_O9;
  constant CFG_GRUSBDC_O10    : integer := CONFIG_GRUSBDC_O10;
  constant CFG_GRUSBDC_O11    : integer := CONFIG_GRUSBDC_O11;
  constant CFG_GRUSBDC_O12    : integer := CONFIG_GRUSBDC_O12;
  constant CFG_GRUSBDC_O13    : integer := CONFIG_GRUSBDC_O13;
  constant CFG_GRUSBDC_O14    : integer := CONFIG_GRUSBDC_O14;
  constant CFG_GRUSBDC_O15    : integer := CONFIG_GRUSBDC_O15;
