-- LCD SVGA controller
  constant CFG_LCD_ENABLE : integer := CONFIG_LCD_ENABLE;

-- LCD 3-wire serial interface
  constant CFG_LCD3T_ENABLE : integer := CONFIG_LCD3T_ENABLE;
  
