-- PROM/SRAM controller
  constant CFG_SRCTRL           : integer := CONFIG_SRCTRL;
  constant CFG_SRCTRL_PROMWS    : integer := CONFIG_SRCTRL_PROMWS;
  constant CFG_SRCTRL_RAMWS     : integer := CONFIG_SRCTRL_RAMWS;
  constant CFG_SRCTRL_IOWS      : integer := CONFIG_SRCTRL_IOWS;
  constant CFG_SRCTRL_RMW       : integer := CONFIG_SRCTRL_RMW;
  constant CFG_SRCTRL_8BIT      : integer := CONFIG_SRCTRL_8BIT;

  constant CFG_SRCTRL_SRBANKS   : integer := CFG_SR_CTRL_SRBANKS;
  constant CFG_SRCTRL_BANKSZ    : integer := CFG_SR_CTRL_BANKSZ;
  constant CFG_SRCTRL_ROMASEL   : integer := CONFIG_SRCTRL_ROMASEL;
