library verilog;
use verilog.vl_types.all;
entity testbench_top is
end testbench_top;
