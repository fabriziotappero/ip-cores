-- SPI controller
  constant CFG_SPICTRL_ENABLE : integer := CONFIG_SPICTRL_ENABLE;
  constant CFG_SPICTRL_SLVS   : integer := CONFIG_SPICTRL_SLVS;
  constant CFG_SPICTRL_FIFO   : integer := CONFIG_SPICTRL_FIFO;
  constant CFG_SPICTRL_SLVREG : integer := CONFIG_SPICTRL_SLVREG;

