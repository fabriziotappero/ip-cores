	//--------------------------------------------------------
	//
	// 128-bit decryption test vectors
	//
	//--------------------------------------------------------
	
	// FIPS-197 Sample Vector 128-bit
	`define FIPS197_128_VEC_SIZE 1
	logic	[0:127]	FIPS197_128_kt[`FIPS197_128_VEC_SIZE] = {128'h000102030405060708090a0b0c0d0e0f};
	logic	[0:127]	FIPS197_128_pt[`FIPS197_128_VEC_SIZE] = {128'h00112233445566778899aabbccddeeff};
	logic	[0:127]	FIPS197_128_ct[`FIPS197_128_VEC_SIZE] = {128'h69c4e0d86a7b0430d8cdb78070b4c55a};
	
	// ECB-AES128.Decrypt sample vector test
	// SP800-38a appendix F.1.2
	`define ECB_DECRYPT_128_VEC_SIZE 4
	int	ECBDecrypt_128_failed = 0;
	logic	[0:127]	ECBDecrypt_128_kt = 128'h2b7e151628aed2a6abf7158809cf4f3c;	
	logic	[0:127]	ECBDecrypt_128_ct [`ECB_DECRYPT_128_VEC_SIZE] = {
	128'h3ad77bb40d7a3660a89ecaf32466ef97,
	128'hf5d3d58503b9699de785895a96fdbaaf,
	128'h43b1cd7f598ece23881b00e3ed030688,
	128'h7b0c785e27e8ad3f8223207104725dd4
	};
	
	logic	[0:127]	ECBDecrypt_128_pt [`ECB_DECRYPT_128_VEC_SIZE] = {
	128'h6bc1bee22e409f96e93d7e117393172a,
	128'hae2d8a571e03ac9c9eb76fac45af8e51,
	128'h30c81c46a35ce411e5fbc1191a0a52ef,
	128'hf69f2445df4f9b17ad2b417be66c3710
	};
	
	// 128-bit GFSbox Known Answer Test vectors.
	// AESAVS appendix B.1
	`define GFSbox_128_VEC_SIZE 7
	int	GFSbox_128_failed=0;
	logic	[0:127]	GFSbox_128_kt = 'h0;
	logic	[0:127]	GFSbox_128_ct[`GFSbox_128_VEC_SIZE] = {
	128'h0336763e966d92595a567cc9ce537f5e,
    128'ha9a1631bf4996954ebc093957b234589,
    128'hff4f8391a6a40ca5b25d23bedd44a597,
    128'hdc43be40be0e53712f7e2bf5ca707209,
    128'h92beedab1895a94faa69b632e5cc47ce,
    128'h459264f4798f6a78bacb89c15ed3d601,
    128'h08a4e2efec8a8e3312ca7460b9040bbf
	};
										
	logic	[0:127]	GFSbox_128_pt[`GFSbox_128_VEC_SIZE] = {
	128'hf34481ec3cc627bacd5dc3fb08f273e6,
	128'h9798c4640bad75c7c3227db910174e72,
	128'h96ab5c2ff612d9dfaae8c31f30c42168,
	128'h6a118a874519e64e9963798a503f1d35,
	128'hcb9fceec81286ca3e989bd979b0cb284,
	128'hb26aeb1874e47ca8358ff22378f09144,
	128'h58c8e00b2631686d54eab84b91f0aca1
	};
	
	// 128-bit KeySBox Known Answer Test vectors
	// AESAVS appendix C.1
	`define KEYSBOX_128_VEC_SIZE 21
	int	KeySbox_128_failed = 0;
	logic	[0:127]	KeySbox_128_pt = 'h0;
	logic	[0:127]	KeySbox_128_ct[`KEYSBOX_128_VEC_SIZE] = {
	128'h6d251e6944b051e04eaa6fb4dbf78465,
    128'h6e29201190152df4ee058139def610bb,
    128'hc3b44b95d9d2f25670eee9a0de099fa3,
    128'h5d9b05578fc944b3cf1ccf0e746cd581,
    128'hf7efc89d5dba578104016ce5ad659c05,
    128'h0306194f666d183624aa230a8b264ae7,
    128'h858075d536d79ccee571f7d7204b1f67,
    128'h35870c6a57e9e92314bcb8087cde72ce,
    128'h6c68e9be5ec41e22c825b7c7affb4363,
    128'hf5df39990fc688f1b07224cc03e86cea,
    128'hbba071bcb470f8f6586e5d3add18bc66,
    128'h43c9f7e62f5d288bb27aa40ef8fe1ea8,
    128'h3580d19cff44f1014a7c966a69059de5,
	128'h806da864dd29d48deafbe764f8202aef,
	128'ha303d940ded8f0baff6f75414cac5243,
	128'hc2dabd117f8a3ecabfbb11d12194d9d0,
	128'hfff60a4740086b3b9c56195b98d91a7b,
	128'h8146a08e2357f0caa30ca8c94d1a0544,
	128'h4b98e06d356deb07ebb824e5713f7be3,
	128'h7a20a53d460fc9ce0423a7a0764c6cf2,
	128'hf4a70d8af877f9b02b4c40df57d45b17	
	};
									
	logic	[0:127]	KeySbox_128_kt[`KEYSBOX_128_VEC_SIZE] = {
	128'h10a58869d74be5a374cf867cfb473859,
    128'hcaea65cdbb75e9169ecd22ebe6e54675,
    128'ha2e2fa9baf7d20822ca9f0542f764a41,
    128'hb6364ac4e1de1e285eaf144a2415f7a0,
    128'h64cf9c7abc50b888af65f49d521944b2,
    128'h47d6742eefcc0465dc96355e851b64d9,
    128'h3eb39790678c56bee34bbcdeccf6cdb5,
    128'h64110a924f0743d500ccadae72c13427,
    128'h18d8126516f8a12ab1a36d9f04d68e51,
    128'hf530357968578480b398a3c251cd1093,
    128'hda84367f325d42d601b4326964802e8e,
    128'he37b1c6aa2846f6fdb413f238b089f23,
    128'h6c002b682483e0cabcc731c253be5674,
	128'h143ae8ed6555aba96110ab58893a8ae1,
	128'hb69418a85332240dc82492353956ae0c,
	128'h71b5c08a1993e1362e4d0ce9b22b78d5,
    128'he234cdca2606b81f29408d5f6da21206,
    128'h13237c49074a3da078dc1d828bb78c6f,
    128'h3071a2a48fe6cbd04f1a129098e308f8,
    128'h90f42ec0f68385f2ffc5dfc03a654dce,
    128'hfebd9a24d8b65c1c787d50a4ed3619a9
	};
	
	// 128-bit VarTxt Known Answer Test vectors
	// AESAVS appendix D.1
	`define VARTXT_128_VEC_SIZE 128
	int	VarTxt_128_failed = 0;
	logic	[0:127]	VarTxt_128_kt = 'h0;
	logic	[0:127]	VarTxt_128_pt[`VARTXT_128_VEC_SIZE] = {
	128'h80000000000000000000000000000000, 
	128'hc0000000000000000000000000000000, 
	128'he0000000000000000000000000000000, 
	128'hf0000000000000000000000000000000, 
	128'hf8000000000000000000000000000000, 
	128'hfc000000000000000000000000000000, 
	128'hfe000000000000000000000000000000, 
	128'hff000000000000000000000000000000, 
	128'hff800000000000000000000000000000, 
	128'hffc00000000000000000000000000000, 
	128'hffe00000000000000000000000000000, 
	128'hfff00000000000000000000000000000, 
	128'hfff80000000000000000000000000000, 
	128'hfffc0000000000000000000000000000, 
	128'hfffe0000000000000000000000000000, 
	128'hffff0000000000000000000000000000, 
	128'hffff8000000000000000000000000000, 
	128'hffffc000000000000000000000000000, 
	128'hffffe000000000000000000000000000, 
	128'hfffff000000000000000000000000000, 
	128'hfffff800000000000000000000000000, 
	128'hfffffc00000000000000000000000000, 
	128'hfffffe00000000000000000000000000, 
	128'hffffff00000000000000000000000000, 
	128'hffffff80000000000000000000000000, 
	128'hffffffc0000000000000000000000000, 
	128'hffffffe0000000000000000000000000, 
	128'hfffffff0000000000000000000000000, 
	128'hfffffff8000000000000000000000000, 
	128'hfffffffc000000000000000000000000, 
	128'hfffffffe000000000000000000000000, 
	128'hffffffff000000000000000000000000, 
	128'hffffffff800000000000000000000000, 
	128'hffffffffc00000000000000000000000, 
	128'hffffffffe00000000000000000000000, 
	128'hfffffffff00000000000000000000000, 
	128'hfffffffff80000000000000000000000, 
	128'hfffffffffc0000000000000000000000, 
	128'hfffffffffe0000000000000000000000, 
	128'hffffffffff0000000000000000000000, 
	128'hffffffffff8000000000000000000000, 
	128'hffffffffffc000000000000000000000, 
	128'hffffffffffe000000000000000000000, 
	128'hfffffffffff000000000000000000000, 
	128'hfffffffffff800000000000000000000, 
	128'hfffffffffffc00000000000000000000, 
	128'hfffffffffffe00000000000000000000, 
	128'hffffffffffff00000000000000000000, 
	128'hffffffffffff80000000000000000000, 
	128'hffffffffffffc0000000000000000000, 
	128'hffffffffffffe0000000000000000000, 
	128'hfffffffffffff0000000000000000000, 
	128'hfffffffffffff8000000000000000000, 
	128'hfffffffffffffc000000000000000000, 
	128'hfffffffffffffe000000000000000000, 
	128'hffffffffffffff000000000000000000, 
	128'hffffffffffffff800000000000000000, 
	128'hffffffffffffffc00000000000000000, 
	128'hffffffffffffffe00000000000000000, 
	128'hfffffffffffffff00000000000000000, 
	128'hfffffffffffffff80000000000000000, 
	128'hfffffffffffffffc0000000000000000, 
	128'hfffffffffffffffe0000000000000000, 
	128'hffffffffffffffff0000000000000000, 
	128'hffffffffffffffff8000000000000000, 
	128'hffffffffffffffffc000000000000000, 
	128'hffffffffffffffffe000000000000000, 
	128'hfffffffffffffffff000000000000000, 
	128'hfffffffffffffffff800000000000000, 
	128'hfffffffffffffffffc00000000000000, 
	128'hfffffffffffffffffe00000000000000, 
	128'hffffffffffffffffff00000000000000, 
	128'hffffffffffffffffff80000000000000, 
	128'hffffffffffffffffffc0000000000000, 
	128'hffffffffffffffffffe0000000000000, 
	128'hfffffffffffffffffff0000000000000, 
	128'hfffffffffffffffffff8000000000000, 
	128'hfffffffffffffffffffc000000000000, 
	128'hfffffffffffffffffffe000000000000, 
	128'hffffffffffffffffffff000000000000, 
	128'hffffffffffffffffffff800000000000, 
	128'hffffffffffffffffffffc00000000000, 
	128'hffffffffffffffffffffe00000000000, 
	128'hfffffffffffffffffffff00000000000, 
	128'hfffffffffffffffffffff80000000000, 
	128'hfffffffffffffffffffffc0000000000, 
	128'hfffffffffffffffffffffe0000000000, 
	128'hffffffffffffffffffffff0000000000, 
	128'hffffffffffffffffffffff8000000000, 
	128'hffffffffffffffffffffffc000000000, 
	128'hffffffffffffffffffffffe000000000, 
	128'hfffffffffffffffffffffff000000000, 
	128'hfffffffffffffffffffffff800000000, 
	128'hfffffffffffffffffffffffc00000000, 
	128'hfffffffffffffffffffffffe00000000, 
	128'hffffffffffffffffffffffff00000000, 
	128'hffffffffffffffffffffffff80000000, 
	128'hffffffffffffffffffffffffc0000000, 
	128'hffffffffffffffffffffffffe0000000, 
	128'hfffffffffffffffffffffffff0000000, 
	128'hfffffffffffffffffffffffff8000000, 
	128'hfffffffffffffffffffffffffc000000, 
	128'hfffffffffffffffffffffffffe000000, 
	128'hffffffffffffffffffffffffff000000, 
	128'hffffffffffffffffffffffffff800000, 
	128'hffffffffffffffffffffffffffc00000, 
	128'hffffffffffffffffffffffffffe00000, 
	128'hfffffffffffffffffffffffffff00000, 
	128'hfffffffffffffffffffffffffff80000, 
	128'hfffffffffffffffffffffffffffc0000, 
	128'hfffffffffffffffffffffffffffe0000, 
	128'hffffffffffffffffffffffffffff0000, 
	128'hffffffffffffffffffffffffffff8000, 
	128'hffffffffffffffffffffffffffffc000, 
	128'hffffffffffffffffffffffffffffe000, 
	128'hfffffffffffffffffffffffffffff000, 
	128'hfffffffffffffffffffffffffffff800, 
	128'hfffffffffffffffffffffffffffffc00, 
	128'hfffffffffffffffffffffffffffffe00, 
	128'hffffffffffffffffffffffffffffff00, 
	128'hffffffffffffffffffffffffffffff80, 
	128'hffffffffffffffffffffffffffffffc0, 
	128'hffffffffffffffffffffffffffffffe0, 
	128'hfffffffffffffffffffffffffffffff0, 
	128'hfffffffffffffffffffffffffffffff8, 
	128'hfffffffffffffffffffffffffffffffc, 
	128'hfffffffffffffffffffffffffffffffe, 
	128'hffffffffffffffffffffffffffffffff
	}; 
	
	logic	[0:127]	VarTxt_128_ct[`VARTXT_128_VEC_SIZE] = {
	128'h3ad78e726c1ec02b7ebfe92b23d9ec34,
	128'haae5939c8efdf2f04e60b9fe7117b2c2,
	128'hf031d4d74f5dcbf39daaf8ca3af6e527,
	128'h96d9fd5cc4f07441727df0f33e401a36,
	128'h30ccdb044646d7e1f3ccea3dca08b8c0,
	128'h16ae4ce5042a67ee8e177b7c587ecc82,
	128'hb6da0bb11a23855d9c5cb1b4c6412e0a,
	128'hdb4f1aa530967d6732ce4715eb0ee24b,
	128'ha81738252621dd180a34f3455b4baa2f,
	128'h77e2b508db7fd89234caf7939ee5621a,
	128'hb8499c251f8442ee13f0933b688fcd19,
	128'h965135f8a81f25c9d630b17502f68e53,
	128'h8b87145a01ad1c6cede995ea3670454f,
	128'h8eae3b10a0c8ca6d1d3b0fa61e56b0b2,
	128'h64b4d629810fda6bafdf08f3b0d8d2c5,
	128'hd7e5dbd3324595f8fdc7d7c571da6c2a,
	128'hf3f72375264e167fca9de2c1527d9606,
	128'h8ee79dd4f401ff9b7ea945d86666c13b,
	128'hdd35cea2799940b40db3f819cb94c08b,
	128'h6941cb6b3e08c2b7afa581ebdd607b87,
	128'h2c20f439f6bb097b29b8bd6d99aad799,
	128'h625d01f058e565f77ae86378bd2c49b3,
	128'hc0b5fd98190ef45fbb4301438d095950,
	128'h13001ff5d99806efd25da34f56be854b,
	128'h3b594c60f5c8277a5113677f94208d82,
	128'he9c0fc1818e4aa46bd2e39d638f89e05,
	128'hf8023ee9c3fdc45a019b4e985c7e1a54,
	128'h35f40182ab4662f3023baec1ee796b57,
	128'h3aebbad7303649b4194a6945c6cc3694,
	128'ha2124bea53ec2834279bed7f7eb0f938,
	128'hb9fb4399fa4facc7309e14ec98360b0a,
	128'hc26277437420c5d634f715aea81a9132,
	128'h171a0e1b2dd424f0e089af2c4c10f32f,
	128'h7cadbe402d1b208fe735edce00aee7ce,
	128'h43b02ff929a1485af6f5c6d6558baa0f,
	128'h092faacc9bf43508bf8fa8613ca75dea,
	128'hcb2bf8280f3f9742c7ed513fe802629c,
	128'h215a41ee442fa992a6e323986ded3f68,
	128'hf21e99cf4f0f77cea836e11a2fe75fb1,
	128'h95e3a0ca9079e646331df8b4e70d2cd6,
	128'h4afe7f120ce7613f74fc12a01a828073,
	128'h827f000e75e2c8b9d479beed913fe678,
	128'h35830c8e7aaefe2d30310ef381cbf691,
	128'h191aa0f2c8570144f38657ea4085ebe5,
	128'h85062c2c909f15d9269b6c18ce99c4f0,
	128'h678034dc9e41b5a560ed239eeab1bc78,
	128'hc2f93a4ce5ab6d5d56f1b93cf19911c1,
	128'h1c3112bcb0c1dcc749d799743691bf82,
	128'h00c55bd75c7f9c881989d3ec1911c0d4,
	128'hea2e6b5ef182b7dff3629abd6a12045f,
	128'h22322327e01780b17397f24087f8cc6f,
	128'hc9cacb5cd11692c373b2411768149ee7,
	128'ha18e3dbbca577860dab6b80da3139256,
	128'h79b61c37bf328ecca8d743265a3d425c,
	128'hd2d99c6bcc1f06fda8e27e8ae3f1ccc7,
	128'h1bfd4b91c701fd6b61b7f997829d663b,
	128'h11005d52f25f16bdc9545a876a63490a,
	128'h3a4d354f02bb5a5e47d39666867f246a,
	128'hd451b8d6e1e1a0ebb155fbbf6e7b7dc3,
	128'h6898d4f42fa7ba6a10ac05e87b9f2080,
	128'hb611295e739ca7d9b50f8e4c0e754a3f,
	128'h7d33fc7d8abe3ca1936759f8f5deaf20,
	128'h3b5e0f566dc96c298f0c12637539b25c,
	128'hf807c3e7985fe0f5a50e2cdb25c5109e,
	128'h41f992a856fb278b389a62f5d274d7e9,
	128'h10d3ed7a6fe15ab4d91acbc7d0767ab1,
	128'h21feecd45b2e675973ac33bf0c5424fc,
	128'h1480cb3955ba62d09eea668f7c708817,
	128'h66404033d6b72b609354d5496e7eb511,
	128'h1c317a220a7d700da2b1e075b00266e1,
	128'hab3b89542233f1271bf8fd0c0f403545,
	128'hd93eae966fac46dca927d6b114fa3f9e,
	128'h1bdec521316503d9d5ee65df3ea94ddf,
	128'heef456431dea8b4acf83bdae3717f75f,
	128'h06f2519a2fafaa596bfef5cfa15c21b9,
	128'h251a7eac7e2fe809e4aa8d0d7012531a,
	128'h3bffc16e4c49b268a20f8d96a60b4058,
	128'he886f9281999c5bb3b3e8862e2f7c988,
	128'h563bf90d61beef39f48dd625fcef1361,
	128'h4d37c850644563c69fd0acd9a049325b,
	128'hb87c921b91829ef3b13ca541ee1130a6,
	128'h2e65eb6b6ea383e109accce8326b0393,
	128'h9ca547f7439edc3e255c0f4d49aa8990,
	128'ha5e652614c9300f37816b1f9fd0c87f9,
	128'h14954f0b4697776f44494fe458d814ed,
	128'h7c8d9ab6c2761723fe42f8bb506cbcf7,
	128'hdb7e1932679fdd99742aab04aa0d5a80,
	128'h4c6a1c83e568cd10f27c2d73ded19c28,
	128'h90ecbe6177e674c98de412413f7ac915,
	128'h90684a2ac55fe1ec2b8ebd5622520b73,
	128'h7472f9a7988607ca79707795991035e6,
	128'h56aff089878bf3352f8df172a3ae47d8,
	128'h65c0526cbe40161b8019a2a3171abd23,
	128'h377be0be33b4e3e310b4aabda173f84f,
	128'h9402e9aa6f69de6504da8d20c4fcaa2f,
	128'h123c1f4af313ad8c2ce648b2e71fb6e1,
	128'h1ffc626d30203dcdb0019fb80f726cf4,
	128'h76da1fbe3a50728c50fd2e621b5ad885,
	128'h082eb8be35f442fb52668e16a591d1d6,
	128'he656f9ecf5fe27ec3e4a73d00c282fb3,
	128'h2ca8209d63274cd9a29bb74bcd77683a,
	128'h79bf5dce14bb7dd73a8e3611de7ce026,
	128'h3c849939a5d29399f344c4a0eca8a576,
	128'hed3c0a94d59bece98835da7aa4f07ca2,
	128'h63919ed4ce10196438b6ad09d99cd795,
	128'h7678f3a833f19fea95f3c6029e2bc610,
	128'h3aa426831067d36b92be7c5f81c13c56,
	128'h9272e2d2cdd11050998c845077a30ea0,
	128'h088c4b53f5ec0ff814c19adae7f6246c,
	128'h4010a5e401fdf0a0354ddbcc0d012b17,
	128'ha87a385736c0a6189bd6589bd8445a93,
	128'h545f2b83d9616dccf60fa9830e9cd287,
	128'h4b706f7f92406352394037a6d4f4688d,
	128'hb7972b3941c44b90afa7b264bfba7387,
	128'h6f45732cf10881546f0fd23896d2bb60,
	128'h2e3579ca15af27f64b3c955a5bfc30ba,
	128'h34a2c5a91ae2aec99b7d1b5fa6780447,
	128'ha4d6616bd04f87335b0e53351227a9ee,
	128'h7f692b03945867d16179a8cefc83ea3f,
	128'h3bd141ee84a0e6414a26e7a4f281f8a2,
	128'hd1788f572d98b2b16ec5d5f3922b99bc,
	128'h0833ff6f61d98a57b288e8c3586b85a6,
	128'h8568261797de176bf0b43becc6285afb,
	128'hf9b0fda0c4a898f5b9e6f661c4ce4d07,
	128'h8ade895913685c67c5269f8aae42983e,
	128'h39bde67d5c8ed8a8b1c37eb8fa9f5ac0,
	128'h5c005e72c1418c44f569f2ea33ba54f3,
	128'h3f5b8cc9ea855a0afa7347d23e8d664e
	};
	
	// 128-bit VarKey Known Answer Test
	// AESAVS appendix E.1
	`define VARKEY_128_VEC_SIZE 128
	int	VarKey_128_failed = 0;
	logic	[0:127]	VarKey_128_pt = 'h0;
	logic	[0:127]	VarKey_128_kt[`VARKEY_128_VEC_SIZE] = {
	128'h80000000000000000000000000000000,	
	128'hc0000000000000000000000000000000,	
	128'he0000000000000000000000000000000,	
	128'hf0000000000000000000000000000000,	
	128'hf8000000000000000000000000000000,	
	128'hfc000000000000000000000000000000,	
	128'hfe000000000000000000000000000000,	
	128'hff000000000000000000000000000000,	
	128'hff800000000000000000000000000000,	
	128'hffc00000000000000000000000000000,	
	128'hffe00000000000000000000000000000,	
	128'hfff00000000000000000000000000000,	
	128'hfff80000000000000000000000000000,	
	128'hfffc0000000000000000000000000000,	
	128'hfffe0000000000000000000000000000,	
	128'hffff0000000000000000000000000000,	
	128'hffff8000000000000000000000000000,	
	128'hffffc000000000000000000000000000,	
	128'hffffe000000000000000000000000000,	
	128'hfffff000000000000000000000000000,	
	128'hfffff800000000000000000000000000,	
	128'hfffffc00000000000000000000000000,	
	128'hfffffe00000000000000000000000000,	
	128'hffffff00000000000000000000000000,	
	128'hffffff80000000000000000000000000,	
	128'hffffffc0000000000000000000000000,	
	128'hffffffe0000000000000000000000000,	
	128'hfffffff0000000000000000000000000,	
	128'hfffffff8000000000000000000000000,	
	128'hfffffffc000000000000000000000000,	
	128'hfffffffe000000000000000000000000,	
	128'hffffffff000000000000000000000000,	
	128'hffffffff800000000000000000000000,	
	128'hffffffffc00000000000000000000000,	
	128'hffffffffe00000000000000000000000,	
	128'hfffffffff00000000000000000000000,	
	128'hfffffffff80000000000000000000000,	
	128'hfffffffffc0000000000000000000000,	
	128'hfffffffffe0000000000000000000000,	
	128'hffffffffff0000000000000000000000,	
	128'hffffffffff8000000000000000000000,	
	128'hffffffffffc000000000000000000000,	
	128'hffffffffffe000000000000000000000,	
	128'hfffffffffff000000000000000000000,	
	128'hfffffffffff800000000000000000000,	
	128'hfffffffffffc00000000000000000000,	
	128'hfffffffffffe00000000000000000000,	
	128'hffffffffffff00000000000000000000,	
	128'hffffffffffff80000000000000000000,	
	128'hffffffffffffc0000000000000000000,	
	128'hffffffffffffe0000000000000000000,	
	128'hfffffffffffff0000000000000000000,	
	128'hfffffffffffff8000000000000000000,	
	128'hfffffffffffffc000000000000000000,	
	128'hfffffffffffffe000000000000000000,	
	128'hffffffffffffff000000000000000000,	
	128'hffffffffffffff800000000000000000,	
	128'hffffffffffffffc00000000000000000,	
	128'hffffffffffffffe00000000000000000,	
	128'hfffffffffffffff00000000000000000,	
	128'hfffffffffffffff80000000000000000,	
	128'hfffffffffffffffc0000000000000000,	
	128'hfffffffffffffffe0000000000000000,	
	128'hffffffffffffffff0000000000000000,	
	128'hffffffffffffffff8000000000000000,	
	128'hffffffffffffffffc000000000000000,	
	128'hffffffffffffffffe000000000000000,	
	128'hfffffffffffffffff000000000000000,	
	128'hfffffffffffffffff800000000000000,	
	128'hfffffffffffffffffc00000000000000,	
	128'hfffffffffffffffffe00000000000000,	
	128'hffffffffffffffffff00000000000000,	
	128'hffffffffffffffffff80000000000000,	
	128'hffffffffffffffffffc0000000000000,	
	128'hffffffffffffffffffe0000000000000,	
	128'hfffffffffffffffffff0000000000000,	
	128'hfffffffffffffffffff8000000000000,	
	128'hfffffffffffffffffffc000000000000,	
	128'hfffffffffffffffffffe000000000000,	
	128'hffffffffffffffffffff000000000000,	
	128'hffffffffffffffffffff800000000000,	
	128'hffffffffffffffffffffc00000000000,	
	128'hffffffffffffffffffffe00000000000,	
	128'hfffffffffffffffffffff00000000000,	
	128'hfffffffffffffffffffff80000000000,	
	128'hfffffffffffffffffffffc0000000000,	
	128'hfffffffffffffffffffffe0000000000,	
	128'hffffffffffffffffffffff0000000000,	
	128'hffffffffffffffffffffff8000000000,	
	128'hffffffffffffffffffffffc000000000,	
	128'hffffffffffffffffffffffe000000000,	
	128'hfffffffffffffffffffffff000000000,	
	128'hfffffffffffffffffffffff800000000,	
	128'hfffffffffffffffffffffffc00000000,	
	128'hfffffffffffffffffffffffe00000000,	
	128'hffffffffffffffffffffffff00000000,	
	128'hffffffffffffffffffffffff80000000,	
	128'hffffffffffffffffffffffffc0000000,	
	128'hffffffffffffffffffffffffe0000000,	
	128'hfffffffffffffffffffffffff0000000,	
	128'hfffffffffffffffffffffffff8000000,	
	128'hfffffffffffffffffffffffffc000000,	
	128'hfffffffffffffffffffffffffe000000,	
	128'hffffffffffffffffffffffffff000000,	
	128'hffffffffffffffffffffffffff800000,	
	128'hffffffffffffffffffffffffffc00000,	
	128'hffffffffffffffffffffffffffe00000,	
	128'hfffffffffffffffffffffffffff00000,	
	128'hfffffffffffffffffffffffffff80000,	
	128'hfffffffffffffffffffffffffffc0000,	
	128'hfffffffffffffffffffffffffffe0000,	
	128'hffffffffffffffffffffffffffff0000,	
	128'hffffffffffffffffffffffffffff8000,	
	128'hffffffffffffffffffffffffffffc000,	
	128'hffffffffffffffffffffffffffffe000,	
	128'hfffffffffffffffffffffffffffff000,	
	128'hfffffffffffffffffffffffffffff800,	
	128'hfffffffffffffffffffffffffffffc00,	
	128'hfffffffffffffffffffffffffffffe00,	
	128'hffffffffffffffffffffffffffffff00,	
	128'hffffffffffffffffffffffffffffff80,	
	128'hffffffffffffffffffffffffffffffc0,	
	128'hffffffffffffffffffffffffffffffe0,	
	128'hfffffffffffffffffffffffffffffff0,	
	128'hfffffffffffffffffffffffffffffff8,	
	128'hfffffffffffffffffffffffffffffffc,	
	128'hfffffffffffffffffffffffffffffffe,	
	128'hffffffffffffffffffffffffffffffff
	};
	
	logic	[0:127]	VarKey_128_ct[`VARKEY_128_VEC_SIZE] = {
	128'h0edd33d3c621e546455bd8ba1418bec8,	
	128'h4bc3f883450c113c64ca42e1112a9e87,	
	128'h72a1da770f5d7ac4c9ef94d822affd97,	
	128'h970014d634e2b7650777e8e84d03ccd8,	
	128'hf17e79aed0db7e279e955b5f493875a7,	
	128'h9ed5a75136a940d0963da379db4af26a,	
	128'hc4295f83465c7755e8fa364bac6a7ea5,	
	128'hb1d758256b28fd850ad4944208cf1155,	
	128'h42ffb34c743de4d88ca38011c990890b,	
	128'h9958f0ecea8b2172c0c1995f9182c0f3,	
	128'h956d7798fac20f82a8823f984d06f7f5,	
	128'ha01bf44f2d16be928ca44aaf7b9b106b,	
	128'hb5f1a33e50d40d103764c76bd4c6b6f8,	
	128'h2637050c9fc0d4817e2d69de878aee8d,	
	128'h113ecbe4a453269a0dd26069467fb5b5,	
	128'h97d0754fe68f11b9e375d070a608c884,	
	128'hc6a0b3e998d05068a5399778405200b4,	
	128'hdf556a33438db87bc41b1752c55e5e49,	
	128'h90fb128d3a1af6e548521bb962bf1f05,	
	128'h26298e9c1db517c215fadfb7d2a8d691,	
	128'ha6cb761d61f8292d0df393a279ad0380,	
	128'h12acd89b13cd5f8726e34d44fd486108,	
	128'h95b1703fc57ba09fe0c3580febdd7ed4,	
	128'hde11722d893e9f9121c381becc1da59a,	
	128'h6d114ccb27bf391012e8974c546d9bf2,	
	128'h5ce37e17eb4646ecfac29b9cc38d9340,	
	128'h18c1b6e2157122056d0243d8a165cddb,	
	128'h99693e6a59d1366c74d823562d7e1431,	
	128'h6c7c64dc84a8bba758ed17eb025a57e3,	
	128'he17bc79f30eaab2fac2cbbe3458d687a,	
	128'h1114bc2028009b923f0b01915ce5e7c4,	
	128'h9c28524a16a1e1c1452971caa8d13476,	
	128'hed62e16363638360fdd6ad62112794f0,	
	128'h5a8688f0b2a2c16224c161658ffd4044,	
	128'h23f710842b9bb9c32f26648c786807ca,	
	128'h44a98bf11e163f632c47ec6a49683a89,	
	128'h0f18aff94274696d9b61848bd50ac5e5,	
	128'h82408571c3e2424540207f833b6dda69,	
	128'h303ff996947f0c7d1f43c8f3027b9b75,	
	128'h7df4daf4ad29a3615a9b6ece5c99518a,	
	128'hc72954a48d0774db0b4971c526260415,	
	128'h1df9b76112dc6531e07d2cfda04411f0,	
	128'h8e4d8e699119e1fc87545a647fb1d34f,	
	128'he6c4807ae11f36f091c57d9fb68548d1,	
	128'h8ebf73aad49c82007f77a5c1ccec6ab4,	
	128'h4fb288cc2040049001d2c7585ad123fc,	
	128'h04497110efb9dceb13e2b13fb4465564,	
	128'h75550e6cb5a88e49634c9ab69eda0430,	
	128'hb6768473ce9843ea66a81405dd50b345,	
	128'hcb2f430383f9084e03a653571e065de6,	
	128'hff4e66c07bae3e79fb7d210847a3b0ba,	
	128'h7b90785125505fad59b13c186dd66ce3,	
	128'h8b527a6aebdaec9eaef8eda2cb7783e5,	
	128'h43fdaf53ebbc9880c228617d6a9b548b,	
	128'h53786104b9744b98f052c46f1c850d0b,	
	128'hb5ab3013dd1e61df06cbaf34ca2aee78,	
	128'h7470469be9723030fdcc73a8cd4fbb10,	
	128'ha35a63f5343ebe9ef8167bcb48ad122e,	
	128'hfd8687f0757a210e9fdf181204c30863,	
	128'h7a181e84bd5457d26a88fbae96018fb0,	
	128'h653317b9362b6f9b9e1a580e68d494b5,	
	128'h995c9dc0b689f03c45867b5faa5c18d1,	
	128'h77a4d96d56dda398b9aabecfc75729fd,	
	128'h84be19e053635f09f2665e7bae85b42d,	
	128'h32cd652842926aea4aa6137bb2be2b5e,	
	128'h493d4a4f38ebb337d10aa84e9171a554,	
	128'hd9bff7ff454b0ec5a4a2a69566e2cb84,	
	128'h3535d565ace3f31eb249ba2cc6765d7a,	
	128'hf60e91fc3269eecf3231c6e9945697c6,	
	128'hab69cfadf51f8e604d9cc37182f6635a,	
	128'h7866373f24a0b6ed56e0d96fcdafb877,	
	128'h1ea448c2aac954f5d812e9d78494446a,	
	128'hacc5599dd8ac02239a0fef4a36dd1668,	
	128'hd8764468bb103828cf7e1473ce895073,	
	128'h1b0d02893683b9f180458e4aa6b73982,	
	128'h96d9b017d302df410a937dcdb8bb6e43,	
	128'hef1623cc44313cff440b1594a7e21cc6,	
	128'h284ca2fa35807b8b0ae4d19e11d7dbd7,	
	128'hf2e976875755f9401d54f36e2a23a594,	
	128'hec198a18e10e532403b7e20887c8dd80,	
	128'h545d50ebd919e4a6949d96ad47e46a80,	
	128'hdbdfb527060e0a71009c7bb0c68f1d44,	
	128'h9cfa1322ea33da2173a024f2ff0d896d,	
	128'h8785b1a75b0f3bd958dcd0e29318c521,	
	128'h38f67b9e98e4a97b6df030a9fcdd0104,	
	128'h192afffb2c880e82b05926d0fc6c448b,	
	128'h6a7980ce7b105cf530952d74daaf798c,	
	128'hea3695e1351b9d6858bd958cf513ef6c,	
	128'h6da0490ba0ba0343b935681d2cce5ba1,	
	128'hf0ea23af08534011c60009ab29ada2f1,	
	128'hff13806cf19cc38721554d7c0fcdcd4b,	
	128'h6838af1f4f69bae9d85dd188dcdf0688,	
	128'h36cf44c92d550bfb1ed28ef583ddf5d7,	
	128'hd06e3195b5376f109d5c4ec6c5d62ced,	
	128'hc440de014d3d610707279b13242a5c36,	
	128'hf0c5c6ffa5e0bd3a94c88f6b6f7c16b9,	
	128'h3e40c3901cd7effc22bffc35dee0b4d9,	
	128'hb63305c72bedfab97382c406d0c49bc6,	
	128'h36bbaab22a6bd4925a99a2b408d2dbae,	
	128'h307c5b8fcd0533ab98bc51e27a6ce461,	
	128'h829c04ff4c07513c0b3ef05c03e337b5,	
	128'hf17af0e895dda5eb98efc68066e84c54,	
	128'h277167f3812afff1ffacb4a934379fc3,	
	128'h2cb1dc3a9c72972e425ae2ef3eb597cd,	
	128'h36aeaa3a213e968d4b5b679d3a2c97fe,	
	128'h9241daca4fdd034a82372db50e1a0f3f,	
	128'hc14574d9cd00cf2b5a7f77e53cd57885,	
	128'h793de39236570aba83ab9b737cb521c9,	
	128'h16591c0f27d60e29b85a96c33861a7ef,	
	128'h44fb5c4d4f5cb79be5c174a3b1c97348,	
	128'h674d2b61633d162be59dde04222f4740,	
	128'hb4750ff263a65e1f9e924ccfd98f3e37,	
	128'h62d0662d6eaeddedebae7f7ea3a4f6b6,	
	128'h70c46bb30692be657f7eaa93ebad9897,	
	128'h323994cfb9da285a5d9642e1759b224a,	
	128'h1dbf57877b7b17385c85d0b54851e371,	
	128'hdfa5c097cdc1532ac071d57b1d28d1bd,	
	128'h3a0c53fa37311fc10bd2a9981f513174,	
	128'hba4f970c0a25c41814bdae2e506be3b4,	
	128'h2dce3acb727cd13ccd76d425ea56e4f6,	
	128'h5160474d504b9b3eefb68d35f245f4b3,	
	128'h41a8a947766635dec37553d9a6c0cbb7,	
	128'h25d6cfe6881f2bf497dd14cd4ddf445b,	
	128'h41c78c135ed9e98c096640647265da1e,	
	128'h5a4d404d8917e353e92a21072c3b2305,	
	128'h02bc96846b3fdc71643f384cd3cc3eaf,	
	128'h9ba4a9143f4e5d4048521c4f8877d88e,	
	128'ha1f6258c877d5fcd8964484538bfc92c
	};

	//--------------------------------------------------------
	//
	// 192-bit decryption test vectors
	//
	//--------------------------------------------------------
	
	// FIPS-197 Sample Vector 192-bit
	`define FIPS197_192_VEC_SIZE 1
	logic	[0:191]	FIPS197_192_kt[`FIPS197_192_VEC_SIZE] = {192'h000102030405060708090a0b0c0d0e0f1011121314151617};
	logic	[0:127]	FIPS197_192_pt[`FIPS197_192_VEC_SIZE] = {128'h00112233445566778899aabbccddeeff};
	logic	[0:127]	FIPS197_192_ct[`FIPS197_192_VEC_SIZE] = {128'hdda97ca4864cdfe06eaf70a0ec0d7191};
	
	// ECB-AES192.Decrypt sample vector test
	// SP800-38a appendix F.1.4
	`define ECB_DECRYPT_192_VEC_SIZE 4
	int	ECBDecrypt_192_failed = 0;
	logic	[0:191]	ECBDecrypt_192_kt = 192'h8e73b0f7da0e6452c810f32b809079e562f8ead2522c6b7b;	
	logic	[0:127]	ECBDecrypt_192_ct [`ECB_DECRYPT_192_VEC_SIZE] = {
	128'hbd334f1d6e45f25ff712a214571fa5cc,
	128'h974104846d0ad3ad7734ecb3ecee4eef,
	128'hef7afd2270e2e60adce0ba2face6444e,
	128'h9a4b41ba738d6c72fb16691603c18e0e
	};
	
	logic	[0:127]	ECBDecrypt_192_pt [`ECB_DECRYPT_192_VEC_SIZE] = {
	128'h6bc1bee22e409f96e93d7e117393172a,
	128'hae2d8a571e03ac9c9eb76fac45af8e51,
	128'h30c81c46a35ce411e5fbc1191a0a52ef,
	128'hf69f2445df4f9b17ad2b417be66c3710
	};
	
	// 192-bit GFSbox Known Answer Test vectors.
	// AESAVS appendix B.2
	`define GFSbox_192_VEC_SIZE 6
	int	GFSbox_192_failed=0;
	logic	[0:191]	GFSbox_192_kt = 'h0;
	logic	[0:127]	GFSbox_192_ct[`GFSbox_192_VEC_SIZE] = {
	128'h275cfc0413d8ccb70513c3859b1d0f72,
    128'hc9b8135ff1b5adc413dfd053b21bd96d,
    128'h4a3650c3371ce2eb35e389a171427440,
    128'h4f354592ff7c8847d2d0870ca9481b7c,
    128'hd5e08bf9a182e857cf40b3a36ee248cc,
    128'h067cd9d3749207791841562507fa9626
	};
										
	logic	[0:127]	GFSbox_192_pt[`GFSbox_192_VEC_SIZE] = {
	128'h1b077a6af4b7f98229de786d7516b639,
	128'h9c2d8842e5f48f57648205d39a239af1,
	128'hbff52510095f518ecca60af4205444bb,
	128'h51719783d3185a535bd75adc65071ce1,
	128'h26aa49dcfe7629a8901a69a9914e6dfd,
	128'h941a4773058224e1ef66d10e0a6ee782
	};

	// 192-bit KeySBox Known Answer Test vectors
	// AESAVS appendix C.2
	`define KEYSBOX_192_VEC_SIZE 24
	int	KeySbox_192_failed = 0;
	logic	[0:127]	KeySbox_192_pt = 'h0;
	logic	[0:127]	KeySbox_192_ct[`KEYSBOX_192_VEC_SIZE] = {
	128'h0956259c9cd5cfd0181cca53380cde06,
    128'h8e4e18424e591a3d5b6f0876f16f8594,
    128'h93f3270cfc877ef17e106ce938979cb0,
    128'h7f6c25ff41858561bb62f36492e93c29,
    128'h8e06556dcbb00b809a025047cff2a940,
    128'h3608c344868e94555d23a120f8a5502d,
    128'h77da2021935b840b7f5dcc39132da9e5,
    128'h3b7c24f825e3bf9873c9f14d39a0e6f4,
    128'h64ebf95686b353508c90ecd8b6134316,
    128'hff558c5d27210b7929b73fc708eb4cf1,
    128'ha2c3b2a818075490a7b4c14380f02702,
    128'hcfe4d74002696ccf7d87b14a2f9cafc9,
    128'hd2eafd86f63b109b91f5dbb3a3fb7e13,
	128'h9b9fdd1c5975655f539998b306a324af,
	128'hdd619e1cf204446112e0af2b9afa8f8c,
	128'hd4f0aae13c8fe9339fbf9e69ed0ad74d,
	128'h19c80ec4a6deb7e5ed1033dda933498f,
	128'h3cf5e1d21a17956d1dffad6a7c41c659,
	128'h69fd12e8505f8ded2fdcb197a121b362,
	128'h8aa584e2cc4d17417a97cb9a28ba29c8,
	128'habc786fb1edb504580c4d882ef29a0c7,
	128'h2e19fb60a3e1de0166f483c97824a978,
	128'h7656709538dd5fec41e0ce6a0f8e207d,
	128'ha67cf333b314d411d3c0ae6e1cfcd8f5
	};
									
	logic	[0:191]	KeySbox_192_kt[`KEYSBOX_192_VEC_SIZE] = {
	192'he9f065d7c13573587f7875357dfbb16c53489f6a4bd0f7cd,
    192'h15d20f6ebc7e649fd95b76b107e6daba967c8a9484797f29,
    192'ha8a282ee31c03fae4f8e9b8930d5473c2ed695a347e88b7c,
    192'hcd62376d5ebb414917f0c78f05266433dc9192a1ec943300,
    192'h502a6ab36984af268bf423c7f509205207fc1552af4a91e5,
    192'h25a39dbfd8034f71a81f9ceb55026e4037f8f6aa30ab44ce,
    192'he08c15411774ec4a908b64eadc6ac4199c7cd453f3aaef53,
    192'h3b375a1ff7e8d44409696e6326ec9dec86138e2ae010b980,
    192'h950bb9f22cc35be6fe79f52c320af93dec5bc9c0c2f9cd53,
    192'h7001c487cc3e572cfc92f4d0e697d982e8856fdcc957da40,
    192'hf029ce61d4e5a405b41ead0a883cc6a737da2cf50a6c92ae,
    192'h61257134a518a0d57d9d244d45f6498cbc32f2bafc522d79,
    192'hb0ab0a6a818baef2d11fa33eac947284fb7d748cfb75e570,
	192'hee053aa011c8b428cdcc3636313c54d6a03cac01c71579d6,
	192'hd2926527e0aa9f37b45e2ec2ade5853ef807576104c7ace3,
	192'h982215f4e173dfa0fcffe5d3da41c4812c7bcc8ed3540f93,
    192'h98c6b8e01e379fbd14e61af6af891596583565f2a27d59e9,
    192'hb3ad5cea1dddc214ca969ac35f37dae1a9a9d1528f89bb35,
    192'h45899367c3132849763073c435a9288a766c8b9ec2308516,
    192'hec250e04c3903f602647b85a401a1ae7ca2f02f67fa4253e,
    192'hd077a03bd8a38973928ccafe4a9d2f455130bd0af5ae46a9,
	192'hd184c36cf0dddfec39e654195006022237871a47c33d3198,
	192'h4c6994ffa9dcdc805b60c2c0095334c42d95a8fc0ca5b080,
	192'hc88f5b00a4ef9a6840e2acaf33f00a3bdc4e25895303fa72
	};
	
	// 192-bit VarTxt Known Answer Test vectors
	// AESAVS appendix D.2
	`define VARTXT_192_VEC_SIZE 128
	int	VarTxt_192_failed = 0;
	logic	[0:191]	VarTxt_192_kt = 'h0;
	logic	[0:127]	VarTxt_192_pt[`VARTXT_192_VEC_SIZE] = {
	128'h80000000000000000000000000000000, 
	128'hc0000000000000000000000000000000, 
	128'he0000000000000000000000000000000, 
	128'hf0000000000000000000000000000000, 
	128'hf8000000000000000000000000000000, 
	128'hfc000000000000000000000000000000, 
	128'hfe000000000000000000000000000000, 
	128'hff000000000000000000000000000000, 
	128'hff800000000000000000000000000000, 
	128'hffc00000000000000000000000000000, 
	128'hffe00000000000000000000000000000, 
	128'hfff00000000000000000000000000000, 
	128'hfff80000000000000000000000000000, 
	128'hfffc0000000000000000000000000000, 
	128'hfffe0000000000000000000000000000, 
	128'hffff0000000000000000000000000000, 
	128'hffff8000000000000000000000000000, 
	128'hffffc000000000000000000000000000, 
	128'hffffe000000000000000000000000000, 
	128'hfffff000000000000000000000000000, 
	128'hfffff800000000000000000000000000, 
	128'hfffffc00000000000000000000000000, 
	128'hfffffe00000000000000000000000000, 
	128'hffffff00000000000000000000000000, 
	128'hffffff80000000000000000000000000, 
	128'hffffffc0000000000000000000000000, 
	128'hffffffe0000000000000000000000000, 
	128'hfffffff0000000000000000000000000, 
	128'hfffffff8000000000000000000000000, 
	128'hfffffffc000000000000000000000000, 
	128'hfffffffe000000000000000000000000, 
	128'hffffffff000000000000000000000000, 
	128'hffffffff800000000000000000000000, 
	128'hffffffffc00000000000000000000000, 
	128'hffffffffe00000000000000000000000, 
	128'hfffffffff00000000000000000000000, 
	128'hfffffffff80000000000000000000000, 
	128'hfffffffffc0000000000000000000000, 
	128'hfffffffffe0000000000000000000000, 
	128'hffffffffff0000000000000000000000, 
	128'hffffffffff8000000000000000000000, 
	128'hffffffffffc000000000000000000000, 
	128'hffffffffffe000000000000000000000, 
	128'hfffffffffff000000000000000000000, 
	128'hfffffffffff800000000000000000000, 
	128'hfffffffffffc00000000000000000000, 
	128'hfffffffffffe00000000000000000000, 
	128'hffffffffffff00000000000000000000, 
	128'hffffffffffff80000000000000000000, 
	128'hffffffffffffc0000000000000000000, 
	128'hffffffffffffe0000000000000000000, 
	128'hfffffffffffff0000000000000000000, 
	128'hfffffffffffff8000000000000000000, 
	128'hfffffffffffffc000000000000000000, 
	128'hfffffffffffffe000000000000000000, 
	128'hffffffffffffff000000000000000000, 
	128'hffffffffffffff800000000000000000, 
	128'hffffffffffffffc00000000000000000, 
	128'hffffffffffffffe00000000000000000, 
	128'hfffffffffffffff00000000000000000, 
	128'hfffffffffffffff80000000000000000, 
	128'hfffffffffffffffc0000000000000000, 
	128'hfffffffffffffffe0000000000000000, 
	128'hffffffffffffffff0000000000000000, 
	128'hffffffffffffffff8000000000000000, 
	128'hffffffffffffffffc000000000000000, 
	128'hffffffffffffffffe000000000000000, 
	128'hfffffffffffffffff000000000000000, 
	128'hfffffffffffffffff800000000000000, 
	128'hfffffffffffffffffc00000000000000, 
	128'hfffffffffffffffffe00000000000000, 
	128'hffffffffffffffffff00000000000000, 
	128'hffffffffffffffffff80000000000000, 
	128'hffffffffffffffffffc0000000000000, 
	128'hffffffffffffffffffe0000000000000, 
	128'hfffffffffffffffffff0000000000000, 
	128'hfffffffffffffffffff8000000000000, 
	128'hfffffffffffffffffffc000000000000, 
	128'hfffffffffffffffffffe000000000000, 
	128'hffffffffffffffffffff000000000000, 
	128'hffffffffffffffffffff800000000000, 
	128'hffffffffffffffffffffc00000000000, 
	128'hffffffffffffffffffffe00000000000, 
	128'hfffffffffffffffffffff00000000000, 
	128'hfffffffffffffffffffff80000000000, 
	128'hfffffffffffffffffffffc0000000000, 
	128'hfffffffffffffffffffffe0000000000, 
	128'hffffffffffffffffffffff0000000000, 
	128'hffffffffffffffffffffff8000000000, 
	128'hffffffffffffffffffffffc000000000, 
	128'hffffffffffffffffffffffe000000000, 
	128'hfffffffffffffffffffffff000000000, 
	128'hfffffffffffffffffffffff800000000, 
	128'hfffffffffffffffffffffffc00000000, 
	128'hfffffffffffffffffffffffe00000000, 
	128'hffffffffffffffffffffffff00000000, 
	128'hffffffffffffffffffffffff80000000, 
	128'hffffffffffffffffffffffffc0000000, 
	128'hffffffffffffffffffffffffe0000000, 
	128'hfffffffffffffffffffffffff0000000, 
	128'hfffffffffffffffffffffffff8000000, 
	128'hfffffffffffffffffffffffffc000000, 
	128'hfffffffffffffffffffffffffe000000, 
	128'hffffffffffffffffffffffffff000000, 
	128'hffffffffffffffffffffffffff800000, 
	128'hffffffffffffffffffffffffffc00000, 
	128'hffffffffffffffffffffffffffe00000, 
	128'hfffffffffffffffffffffffffff00000, 
	128'hfffffffffffffffffffffffffff80000, 
	128'hfffffffffffffffffffffffffffc0000, 
	128'hfffffffffffffffffffffffffffe0000, 
	128'hffffffffffffffffffffffffffff0000, 
	128'hffffffffffffffffffffffffffff8000, 
	128'hffffffffffffffffffffffffffffc000, 
	128'hffffffffffffffffffffffffffffe000, 
	128'hfffffffffffffffffffffffffffff000, 
	128'hfffffffffffffffffffffffffffff800, 
	128'hfffffffffffffffffffffffffffffc00, 
	128'hfffffffffffffffffffffffffffffe00, 
	128'hffffffffffffffffffffffffffffff00, 
	128'hffffffffffffffffffffffffffffff80, 
	128'hffffffffffffffffffffffffffffffc0, 
	128'hffffffffffffffffffffffffffffffe0, 
	128'hfffffffffffffffffffffffffffffff0, 
	128'hfffffffffffffffffffffffffffffff8, 
	128'hfffffffffffffffffffffffffffffffc, 
	128'hfffffffffffffffffffffffffffffffe, 
	128'hffffffffffffffffffffffffffffffff
	}; 
	
	logic	[0:127]	VarTxt_192_ct[`VARTXT_192_VEC_SIZE] = {
	128'h6cd02513e8d4dc986b4afe087a60bd0c,
	128'h2ce1f8b7e30627c1c4519eada44bc436,
	128'h9946b5f87af446f5796c1fee63a2da24,
	128'h2a560364ce529efc21788779568d5555,
	128'h35c1471837af446153bce55d5ba72a0a,
	128'hce60bc52386234f158f84341e534cd9e,
	128'h8c7c27ff32bcf8dc2dc57c90c2903961,
	128'h32bb6a7ec84499e166f936003d55a5bb,
	128'ha5c772e5c62631ef660ee1d5877f6d1b,
	128'h030d7e5b64f380a7e4ea5387b5cd7f49,
	128'h0dc9a2610037009b698f11bb7e86c83e,
	128'h0046612c766d1840c226364f1fa7ed72,
	128'h4880c7e08f27befe78590743c05e698b,
	128'h2520ce829a26577f0f4822c4ecc87401,
	128'h8765e8acc169758319cb46dc7bcf3dca,
	128'he98f4ba4f073df4baa116d011dc24a28,
	128'hf378f68c5dbf59e211b3a659a7317d94,
	128'h283d3b069d8eb9fb432d74b96ca762b4,
	128'ha7e1842e8a87861c221a500883245c51,
	128'h77aa270471881be070fb52c7067ce732,
	128'h01b0f476d484f43f1aeb6efa9361a8ac,
	128'h1c3a94f1c052c55c2d8359aff2163b4f,
	128'he8a067b604d5373d8b0f2e05a03b341b,
	128'ha7876ec87f5a09bfea42c77da30fd50e,
	128'h0cf3e9d3a42be5b854ca65b13f35f48d,
	128'h6c62f6bbcab7c3e821c9290f08892dda,
	128'h7f5e05bd2068738196fee79ace7e3aec,
	128'h440e0d733255cda92fb46e842fe58054,
	128'haa5d5b1c4ea1b7a22e5583ac2e9ed8a7,
	128'h77e537e89e8491e8662aae3bc809421d,
	128'h997dd3e9f1598bfa73f75973f7e93b76,
	128'h1b38d4f7452afefcb7fc721244e4b72e,
	128'h0be2b18252e774dda30cdda02c6906e3,
	128'hd2695e59c20361d82652d7d58b6f11b2,
	128'h902d88d13eae52089abd6143cfe394e9,
	128'hd49bceb3b823fedd602c305345734bd2,
	128'h707b1dbb0ffa40ef7d95def421233fae,
	128'h7ca0c1d93356d9eb8aa952084d75f913,
	128'hf2cbf9cb186e270dd7bdb0c28febc57d,
	128'hc94337c37c4e790ab45780bd9c3674a0,
	128'h8e3558c135252fb9c9f367ed609467a1,
	128'h1b72eeaee4899b443914e5b3a57fba92,
	128'h011865f91bc56868d051e52c9efd59b7,
	128'he4771318ad7a63dd680f6e583b7747ea,
	128'h61e3d194088dc8d97e9e6db37457eac5,
	128'h36ff1ec9ccfbc349e5d356d063693ad6,
	128'h3cc9e9a9be8cc3f6fb2ea24088e9bb19,
	128'h1ee5ab003dc8722e74905d9a8fe3d350,
	128'h245339319584b0a412412869d6c2eada,
	128'h7bd496918115d14ed5380852716c8814,
	128'h273ab2f2b4a366a57d582a339313c8b1,
	128'h113365a9ffbe3b0ca61e98507554168b,
	128'hafa99c997ac478a0dea4119c9e45f8b1,
	128'h9216309a7842430b83ffb98638011512,
	128'h62abc792288258492a7cb45145f4b759,
	128'h534923c169d504d7519c15d30e756c50,
	128'hfa75e05bcdc7e00c273fa33f6ee441d2,
	128'h7d350fa6057080f1086a56b17ec240db,
	128'hf34e4a6324ea4a5c39a661c8fe5ada8f,
	128'h0882a16f44088d42447a29ac090ec17e,
	128'h3a3c15bfc11a9537c130687004e136ee,
	128'h22c0a7678dc6d8cf5c8a6d5a9960767c,
	128'hb46b09809d68b9a456432a79bdc2e38c,
	128'h93baaffb35fbe739c17c6ac22eecf18f,
	128'hc8aa80a7850675bc007c46df06b49868,
	128'h12c6f3877af421a918a84b775858021d,
	128'h33f123282c5d633924f7d5ba3f3cab11,
	128'ha8f161002733e93ca4527d22c1a0c5bb,
	128'hb72f70ebf3e3fda23f508eec76b42c02,
	128'h6a9d965e6274143f25afdcfc88ffd77c,
	128'ha0c74fd0b9361764ce91c5200b095357,
	128'h091d1fdc2bd2c346cd5046a8c6209146,
	128'he2a37580116cfb71856254496ab0aca8,
	128'he0b3a00785917c7efc9adba322813571,
	128'h733d41f4727b5ef0df4af4cf3cffa0cb,
	128'ha99ebb030260826f981ad3e64490aa4f,
	128'h73f34c7d3eae5e80082c1647524308ee,
	128'h40ebd5ad082345b7a2097ccd3464da02,
	128'h7cc4ae9a424b2cec90c97153c2457ec5,
	128'h54d632d03aba0bd0f91877ebdd4d09cb,
	128'hd3427be7e4d27cd54f5fe37b03cf0897,
	128'hb2099795e88cc158fd75ea133d7e7fbe,
	128'ha6cae46fb6fadfe7a2c302a34242817b,
	128'h026a7024d6a902e0b3ffccbaa910cc3f,
	128'h156f07767a85a4312321f63968338a01,
	128'h15eec9ebf42b9ca76897d2cd6c5a12e2,
	128'hdb0d3a6fdcc13f915e2b302ceeb70fd8,
	128'h71dbf37e87a2e34d15b20e8f10e48924,
	128'hc745c451e96ff3c045e4367c833e3b54,
	128'h340da09c2dd11c3b679d08ccd27dd595,
	128'h8279f7c0c2a03ee660c6d392db025d18,
	128'ha4b2c7d8eba531ff47c5041a55fbd1ec,
	128'h74569a2ca5a7bd5131ce8dc7cbfbf72f,
	128'h3713da0c0219b63454035613b5a403dd,
	128'h8827551ddcc9df23fa72a3de4e9f0b07,
	128'h2e3febfd625bfcd0a2c06eb460da1732,
	128'hee82e6ba488156f76496311da6941deb,
	128'h4770446f01d1f391256e85a1b30d89d3,
	128'haf04b68f104f21ef2afb4767cf74143c,
	128'hcf3579a9ba38c8e43653173e14f3a4c6,
	128'hb3bba904f4953e09b54800af2f62e7d4,
	128'hfc4249656e14b29eb9c44829b4c59a46,
	128'h9b31568febe81cfc2e65af1c86d1a308,
	128'h9ca09c25f273a766db98a480ce8dfedc,
	128'hb909925786f34c3c92d971883c9fbedf,
	128'h82647f1332fe570a9d4d92b2ee771d3b,
	128'h3604a7e80832b3a99954bca6f5b9f501,
	128'h884607b128c5de3ab39a529a1ef51bef,
	128'h670cfa093d1dbdb2317041404102435e,
	128'h7a867195f3ce8769cbd336502fbb5130,
	128'h52efcf64c72b2f7ca5b3c836b1078c15,
	128'h4019250f6eefb2ac5ccbcae044e75c7e,
	128'h022c4f6f5a017d292785627667ddef24,
	128'he9c21078a2eb7e03250f71000fa9e3ed,
	128'ha13eaeeb9cd391da4e2b09490b3e7fad,
	128'hc958a171dca1d4ed53e1af1d380803a9,
	128'h21442e07a110667f2583eaeeee44dc8c,
	128'h59bbb353cf1dd867a6e33737af655e99,
	128'h43cd3b25375d0ce41087ff9fe2829639,
	128'h6b98b17e80d1118e3516bd768b285a84,
	128'hae47ed3676ca0c08deea02d95b81db58,
	128'h34ec40dc20413795ed53628ea748720b,
	128'h4dc68163f8e9835473253542c8a65d46,
	128'h2aabb999f43693175af65c6c612c46fb,
	128'he01f94499dac3547515c5b1d756f0f58,
	128'h9d12435a46480ce00ea349f71799df9a,
	128'hcef41d16d266bdfe46938ad7884cc0cf,
	128'hb13db4da1f718bc6904797c82bcf2d32
	};

	// 192-bit VarKey Known Answer Test
	// AESAVS appendix E.2
	`define VARKEY_192_VEC_SIZE 192
	int	VarKey_192_failed = 0;
	logic	[0:127]	VarKey_192_pt = 'h0;
	logic	[0:191]	VarKey_192_kt[`VARKEY_192_VEC_SIZE] = {
	192'h800000000000000000000000000000000000000000000000,	
	192'hc00000000000000000000000000000000000000000000000,	
	192'he00000000000000000000000000000000000000000000000,	
	192'hf00000000000000000000000000000000000000000000000,	
	192'hf80000000000000000000000000000000000000000000000,	
	192'hfc0000000000000000000000000000000000000000000000,	
	192'hfe0000000000000000000000000000000000000000000000,	
	192'hff0000000000000000000000000000000000000000000000,	
	192'hff8000000000000000000000000000000000000000000000,	
	192'hffc000000000000000000000000000000000000000000000,	
	192'hffe000000000000000000000000000000000000000000000,	
	192'hfff000000000000000000000000000000000000000000000,	
	192'hfff800000000000000000000000000000000000000000000,	
	192'hfffc00000000000000000000000000000000000000000000,	
	192'hfffe00000000000000000000000000000000000000000000,	
	192'hffff00000000000000000000000000000000000000000000,	
	192'hffff80000000000000000000000000000000000000000000,	
	192'hffffc0000000000000000000000000000000000000000000,	
	192'hffffe0000000000000000000000000000000000000000000,	
	192'hfffff0000000000000000000000000000000000000000000,	
	192'hfffff8000000000000000000000000000000000000000000,	
	192'hfffffc000000000000000000000000000000000000000000,	
	192'hfffffe000000000000000000000000000000000000000000,	
	192'hffffff000000000000000000000000000000000000000000,	
	192'hffffff800000000000000000000000000000000000000000,	
	192'hffffffc00000000000000000000000000000000000000000,	
	192'hffffffe00000000000000000000000000000000000000000,	
	192'hfffffff00000000000000000000000000000000000000000,	
	192'hfffffff80000000000000000000000000000000000000000,	
	192'hfffffffc0000000000000000000000000000000000000000,	
	192'hfffffffe0000000000000000000000000000000000000000,	
	192'hffffffff0000000000000000000000000000000000000000,	
	192'hffffffff8000000000000000000000000000000000000000,	
	192'hffffffffc000000000000000000000000000000000000000,	
	192'hffffffffe000000000000000000000000000000000000000,	
	192'hfffffffff000000000000000000000000000000000000000,	
	192'hfffffffff800000000000000000000000000000000000000,	
	192'hfffffffffc00000000000000000000000000000000000000,	
	192'hfffffffffe00000000000000000000000000000000000000,	
	192'hffffffffff00000000000000000000000000000000000000,	
	192'hffffffffff80000000000000000000000000000000000000,	
	192'hffffffffffc0000000000000000000000000000000000000,	
	192'hffffffffffe0000000000000000000000000000000000000,	
	192'hfffffffffff0000000000000000000000000000000000000,	
	192'hfffffffffff8000000000000000000000000000000000000,	
	192'hfffffffffffc000000000000000000000000000000000000,	
	192'hfffffffffffe000000000000000000000000000000000000,	
	192'hffffffffffff000000000000000000000000000000000000,	
	192'hffffffffffff800000000000000000000000000000000000,	
	192'hffffffffffffc00000000000000000000000000000000000,	
	192'hffffffffffffe00000000000000000000000000000000000,	
	192'hfffffffffffff00000000000000000000000000000000000,	
	192'hfffffffffffff80000000000000000000000000000000000,	
	192'hfffffffffffffc0000000000000000000000000000000000,	
	192'hfffffffffffffe0000000000000000000000000000000000,	
	192'hffffffffffffff0000000000000000000000000000000000,	
	192'hffffffffffffff8000000000000000000000000000000000,	
	192'hffffffffffffffc000000000000000000000000000000000,	
	192'hffffffffffffffe000000000000000000000000000000000,	
	192'hfffffffffffffff000000000000000000000000000000000,	
	192'hfffffffffffffff800000000000000000000000000000000,	
	192'hfffffffffffffffc00000000000000000000000000000000,	
	192'hfffffffffffffffe00000000000000000000000000000000,	
	192'hffffffffffffffff00000000000000000000000000000000,	
	192'hffffffffffffffff80000000000000000000000000000000,	
	192'hffffffffffffffffc0000000000000000000000000000000,	
	192'hffffffffffffffffe0000000000000000000000000000000,	
	192'hfffffffffffffffff0000000000000000000000000000000,	
	192'hfffffffffffffffff8000000000000000000000000000000,	
	192'hfffffffffffffffffc000000000000000000000000000000,	
	192'hfffffffffffffffffe000000000000000000000000000000,	
	192'hffffffffffffffffff000000000000000000000000000000,	
	192'hffffffffffffffffff800000000000000000000000000000,	
	192'hffffffffffffffffffc00000000000000000000000000000,	
	192'hffffffffffffffffffe00000000000000000000000000000,	
	192'hfffffffffffffffffff00000000000000000000000000000,	
	192'hfffffffffffffffffff80000000000000000000000000000,	
	192'hfffffffffffffffffffc0000000000000000000000000000,	
	192'hfffffffffffffffffffe0000000000000000000000000000,	
	192'hffffffffffffffffffff0000000000000000000000000000,	
	192'hffffffffffffffffffff8000000000000000000000000000,	
	192'hffffffffffffffffffffc000000000000000000000000000,	
	192'hffffffffffffffffffffe000000000000000000000000000,	
	192'hfffffffffffffffffffff000000000000000000000000000,	
	192'hfffffffffffffffffffff800000000000000000000000000,	
	192'hfffffffffffffffffffffc00000000000000000000000000,	
	192'hfffffffffffffffffffffe00000000000000000000000000,	
	192'hffffffffffffffffffffff00000000000000000000000000,	
	192'hffffffffffffffffffffff80000000000000000000000000,	
	192'hffffffffffffffffffffffc0000000000000000000000000,	
	192'hffffffffffffffffffffffe0000000000000000000000000,	
	192'hfffffffffffffffffffffff0000000000000000000000000,	
	192'hfffffffffffffffffffffff8000000000000000000000000,	
	192'hfffffffffffffffffffffffc000000000000000000000000,	
	192'hfffffffffffffffffffffffe000000000000000000000000,	
	192'hffffffffffffffffffffffff000000000000000000000000,	
	192'hffffffffffffffffffffffff800000000000000000000000,	
	192'hffffffffffffffffffffffffc00000000000000000000000,	
	192'hffffffffffffffffffffffffe00000000000000000000000,	
	192'hfffffffffffffffffffffffff00000000000000000000000,	
	192'hfffffffffffffffffffffffff80000000000000000000000,	
	192'hfffffffffffffffffffffffffc0000000000000000000000,	
	192'hfffffffffffffffffffffffffe0000000000000000000000,	
	192'hffffffffffffffffffffffffff0000000000000000000000,	
	192'hffffffffffffffffffffffffff8000000000000000000000,	
	192'hffffffffffffffffffffffffffc000000000000000000000,	
	192'hffffffffffffffffffffffffffe000000000000000000000,	
	192'hfffffffffffffffffffffffffff000000000000000000000,	
	192'hfffffffffffffffffffffffffff800000000000000000000,	
	192'hfffffffffffffffffffffffffffc00000000000000000000,	
	192'hfffffffffffffffffffffffffffe00000000000000000000,	
	192'hffffffffffffffffffffffffffff00000000000000000000,	
	192'hffffffffffffffffffffffffffff80000000000000000000,	
	192'hffffffffffffffffffffffffffffc0000000000000000000,	
	192'hffffffffffffffffffffffffffffe0000000000000000000,	
	192'hfffffffffffffffffffffffffffff0000000000000000000,	
	192'hfffffffffffffffffffffffffffff8000000000000000000,	
	192'hfffffffffffffffffffffffffffffc000000000000000000,	
	192'hfffffffffffffffffffffffffffffe000000000000000000,	
	192'hffffffffffffffffffffffffffffff000000000000000000,	
	192'hffffffffffffffffffffffffffffff800000000000000000,	
	192'hffffffffffffffffffffffffffffffc00000000000000000,	
	192'hffffffffffffffffffffffffffffffe00000000000000000,	
	192'hfffffffffffffffffffffffffffffff00000000000000000,	
	192'hfffffffffffffffffffffffffffffff80000000000000000,	
	192'hfffffffffffffffffffffffffffffffc0000000000000000,	
	192'hfffffffffffffffffffffffffffffffe0000000000000000,	
	192'hffffffffffffffffffffffffffffffff0000000000000000,
	192'hffffffffffffffffffffffffffffffff8000000000000000,
	192'hffffffffffffffffffffffffffffffffc000000000000000,
	192'hffffffffffffffffffffffffffffffffe000000000000000,
	192'hfffffffffffffffffffffffffffffffff000000000000000,
	192'hfffffffffffffffffffffffffffffffff800000000000000,
	192'hfffffffffffffffffffffffffffffffffc00000000000000,
	192'hfffffffffffffffffffffffffffffffffe00000000000000,
	192'hffffffffffffffffffffffffffffffffff00000000000000,
	192'hffffffffffffffffffffffffffffffffff80000000000000,
	192'hffffffffffffffffffffffffffffffffffc0000000000000,
	192'hffffffffffffffffffffffffffffffffffe0000000000000,
	192'hfffffffffffffffffffffffffffffffffff0000000000000,
	192'hfffffffffffffffffffffffffffffffffff8000000000000,
	192'hfffffffffffffffffffffffffffffffffffc000000000000,
	192'hfffffffffffffffffffffffffffffffffffe000000000000,
	192'hffffffffffffffffffffffffffffffffffff000000000000,
	192'hffffffffffffffffffffffffffffffffffff800000000000,
	192'hffffffffffffffffffffffffffffffffffffc00000000000,
	192'hffffffffffffffffffffffffffffffffffffe00000000000,
	192'hfffffffffffffffffffffffffffffffffffff00000000000,
	192'hfffffffffffffffffffffffffffffffffffff80000000000,
	192'hfffffffffffffffffffffffffffffffffffffc0000000000,
	192'hfffffffffffffffffffffffffffffffffffffe0000000000,
	192'hffffffffffffffffffffffffffffffffffffff0000000000,
	192'hffffffffffffffffffffffffffffffffffffff8000000000,
	192'hffffffffffffffffffffffffffffffffffffffc000000000,
	192'hffffffffffffffffffffffffffffffffffffffe000000000,
	192'hfffffffffffffffffffffffffffffffffffffff000000000,
	192'hfffffffffffffffffffffffffffffffffffffff800000000,
	192'hfffffffffffffffffffffffffffffffffffffffc00000000,
	192'hfffffffffffffffffffffffffffffffffffffffe00000000,
	192'hffffffffffffffffffffffffffffffffffffffff00000000,
	192'hffffffffffffffffffffffffffffffffffffffff80000000,
	192'hffffffffffffffffffffffffffffffffffffffffc0000000,
	192'hffffffffffffffffffffffffffffffffffffffffe0000000,
	192'hfffffffffffffffffffffffffffffffffffffffff0000000,
	192'hfffffffffffffffffffffffffffffffffffffffff8000000,
	192'hfffffffffffffffffffffffffffffffffffffffffc000000,
	192'hfffffffffffffffffffffffffffffffffffffffffe000000,
	192'hffffffffffffffffffffffffffffffffffffffffff000000,
	192'hffffffffffffffffffffffffffffffffffffffffff800000,
	192'hffffffffffffffffffffffffffffffffffffffffffc00000,
	192'hffffffffffffffffffffffffffffffffffffffffffe00000,
	192'hfffffffffffffffffffffffffffffffffffffffffff00000,
	192'hfffffffffffffffffffffffffffffffffffffffffff80000,
	192'hfffffffffffffffffffffffffffffffffffffffffffc0000,
	192'hfffffffffffffffffffffffffffffffffffffffffffe0000,
	192'hffffffffffffffffffffffffffffffffffffffffffff0000,
	192'hffffffffffffffffffffffffffffffffffffffffffff8000,
	192'hffffffffffffffffffffffffffffffffffffffffffffc000,
	192'hffffffffffffffffffffffffffffffffffffffffffffe000,
	192'hfffffffffffffffffffffffffffffffffffffffffffff000,
	192'hfffffffffffffffffffffffffffffffffffffffffffff800,
	192'hfffffffffffffffffffffffffffffffffffffffffffffc00,
	192'hfffffffffffffffffffffffffffffffffffffffffffffe00,
	192'hffffffffffffffffffffffffffffffffffffffffffffff00,
	192'hffffffffffffffffffffffffffffffffffffffffffffff80,
	192'hffffffffffffffffffffffffffffffffffffffffffffffc0,
	192'hffffffffffffffffffffffffffffffffffffffffffffffe0,
	192'hfffffffffffffffffffffffffffffffffffffffffffffff0,
	192'hfffffffffffffffffffffffffffffffffffffffffffffff8,
	192'hfffffffffffffffffffffffffffffffffffffffffffffffc,
	192'hfffffffffffffffffffffffffffffffffffffffffffffffe,
	192'hffffffffffffffffffffffffffffffffffffffffffffffff
	};                                   
	
	logic	[0:127]	VarKey_192_ct[`VARKEY_192_VEC_SIZE] = {
	128'hde885dc87f5a92594082d02cc1e1b42c,	
	128'h132b074e80f2a597bf5febd8ea5da55e,	
	128'h6eccedf8de592c22fb81347b79f2db1f,	
	128'h180b09f267c45145db2f826c2582d35c,	
	128'hedd807ef7652d7eb0e13c8b5e15b3bc0,	
	128'h9978bcf8dd8fd72241223ad24b31b8a4,	
	128'h5310f654343e8f27e12c83a48d24ff81,	
	128'h833f71258d53036b02952c76c744f5a1,	
	128'heba83ff200cff9318a92f8691a06b09f,	
	128'hff620ccbe9f3292abdf2176b09f04eba,	
	128'h7ababc4b3f516c9aafb35f4140b548f9,	
	128'haa187824d9c4582b0916493ecbde8c57,	
	128'h1c0ad553177fd5ea1092c9d626a29dc4,	
	128'ha5dc46c37261194124ecaebd680408ec,	
	128'he4f2f2ae23e9b10bacfa58601531ba54,	
	128'hb7d67cf1a1e91e8ff3a57a172c7bf412,	
	128'h26706be06967884e847d137128ce47b3,	
	128'hb2f8b409b0585909aad3a7b5a219072a,	
	128'h5e4b7bff0290c78344c54a23b722cd20,	
	128'h07093657552d4414227ce161e9ebf7dd,	
	128'he1af1e7d8bc225ed4dffb771ecbb9e67,	
	128'hef6555253635d8432156cfd9c11b145a,	
	128'hfb4035074a5d4260c90cbd6da6c3fceb,	
	128'h446ee416f9ad1c103eb0cc96751c88e1,	
	128'h198ae2a4637ac0a7890a8fd1485445c9,	
	128'h562012ec8faded0825fb2fa70ab30cbd,	
	128'hcc8a64b46b5d88bf7f247d4dbaf38f05,	
	128'ha168253762e2cc81b42d1e5001762699,	
	128'h1b41f83b38ce5032c6cd7af98cf62061,	
	128'h61a89990cd1411750d5fb0dc988447d4,	
	128'hb5accc8ed629edf8c68a539183b1ea82,	
	128'hb16fa71f846b81a13f361c43a851f290,	
	128'h4fad6efdff5975aee7692234bcd54488,	
	128'hebfdb05a783d03082dfe5fdd80a00b17,	
	128'heb81b584766997af6ba5529d3bdd8609,	
	128'h0cf4ff4f49c8a0ca060c443499e29313,	
	128'hcc4ba8a8e029f8b26d8afff9df133bb6,	
	128'hfefebf64360f38e4e63558f0ffc550c3,	
	128'h12ad98cbf725137d6a8108c2bed99322,	
	128'h6afaa996226198b3e2610413ce1b3f78,	
	128'h2a8ce6747a7e39367828e290848502d9,	
	128'h223736e8b8f89ca1e37b6deab40facf1,	
	128'hc0f797e50418b95fa6013333917a9480,	
	128'ha758de37c2ece2a02c73c01fedc9a132,	
	128'h3a9b87ae77bae706803966c66c73adbd,	
	128'hd365ab8df8ffd782e358121a4a4fc541,	
	128'hc8dcd9e6f75e6c36c8daee0466f0ed74,	
	128'hc79a637beb1c0304f14014c037e736dd,	
	128'h105f0a25e84ac930d996281a5f954dd9,	
	128'h42e4074b2927973e8d17ffa92f7fe615,	
	128'h4fe2a9d2c1824449c69e3e0398f12963,	
	128'hb7f29c1e1f62847a15253b28a1e9d712,	
	128'h36ed5d29b903f31e8983ef8b0a2bf990,	
	128'h27b8070270810f9d023f9dd7ff3b4aa2,	
	128'h94d46e155c1228f61d1a0db4815ecc4b,	
	128'hca6108d1d98071428eeceef1714b96dd,	
	128'hdc5b25b71b6296cf73dd2cdcac2f70b1,	
	128'h44aba95e8a06a2d9d3530d2677878c80,	
	128'ha570d20e89b467e8f5176061b81dd396,	
	128'h758f4467a5d8f1e7307dc30b34e404f4,	
	128'hbcea28e9071b5a2302970ff352451bc5,	
	128'h7523c00bc177d331ad312e09c9015c1c,	
	128'hccac61e3183747b3f5836da21a1bc4f4,	
	128'h707b075791878880b44189d3522b8c30,	
	128'h7132d0c0e4a07593cf12ebb12be7688c,	
	128'heffbac1644deb0c784275fe56e19ead3,	
	128'ha005063f30f4228b374e2459738f26bb,	
	128'h29975b5f48bb68fcbbc7cea93b452ed7,	
	128'hcf3f2576e2afedc74bb1ca7eeec1c0e7,	
	128'h07c403f5f966e0e3d9f296d6226dca28,	
	128'hc8c20908249ab4a34d6dd0a31327ff1a,	
	128'hc0541329ecb6159ab23b7fc5e6a21bca,	
	128'h7aa1acf1a2ed9ba72bc6deb31d88b863,	
	128'h808bd8eddabb6f3bf0d5a8a27be1fe8a,	
	128'h273c7d7685e14ec66bbb96b8f05b6ddd,	
	128'h32752eefc8c2a93f91b6e73eb07cca6e,	
	128'hd893e7d62f6ce502c64f75e281f9c000,	
	128'h8dfd999be5d0cfa35732c0ddc88ff5a5,	
	128'h02647c76a300c3173b841487eb2bae9f,	
	128'h172df8b02f04b53adab028b4e01acd87,	
	128'h054b3bf4998aeb05afd87ec536533a36,	
	128'h3783f7bf44c97f065258a666cae03020,	
	128'haad4c8a63f80954104de7b92cede1be1,	
	128'hcbfe61810fd5467ccdacb75800f3ac07,	
	128'h830d8a2590f7d8e1b55a737f4af45f34,	
	128'hfffcd4683f858058e74314671d43fa2c,	
	128'h523d0babbb82f46ebc9e70b1cd41ddd0,	
	128'h344aab37080d7486f7d542a309e53eed,	
	128'h56c5609d0906b23ab9caca816f5dbebd,	
	128'h7026026eedd91adc6d831cdf9894bdc6,	
	128'h88330baa4f2b618fc9d9b021bf503d5a,	
	128'hfc9e0ea22480b0bac935c8a8ebefcdcf,	
	128'h29ca779f398fb04f867da7e8a44756cb,	
	128'h51f89c42985786bfc43c6df8ada36832,	
	128'h6ac1de5fb8f21d874e91c53b560c50e3,	
	128'h03aa9058490eda306001a8a9f48d0ca7,	
	128'he34ec71d6128d4871865d617c30b37e3,	
	128'h14be1c535b17cabd0c4d93529d69bf47,	
	128'hc9ef67756507beec9dd3862883478044,	
	128'h40e231fa5a5948ce2134e92fc0664d4b,	
	128'h03194b8e5dda5530d0c678c0b48f5d92,	
	128'h90bd086f237cc4fd99f4d76bde6b4826,	
	128'h19259761ca17130d6ed86d57cd7951ee,	
	128'hd7cbb3f34b9b450f24b0e8518e54da6d,	
	128'h725b9caebe9f7f417f4068d0d2ee20b3,	
	128'h9d924b934a90ce1fd39b8a9794f82672,	
	128'hc50562bf094526a91c5bc63c0c224995,	
	128'hd2f11805046743bd74f57188d9188df7,	
	128'h8dd274bd0f1b58ae345d9e7233f9b8f3,	
	128'h9d6bdc8f4ce5feb0f3bed2e4b9a9bb0b,	
	128'hfd5548bcf3f42565f7efa94562528d46,	
	128'hd2ccaebd3a4c3e80b063748131ba4a71,	
	128'he03cb23d9e11c9d93f117e9c0a91b576,	
	128'h78f933a2081ac1db84f69d10f4523fe0,	
	128'h4061f7412ed320de0edc8851c2e2436f,	
	128'h9064ba1cd04ce6bab98474330814b4d4,	
	128'h48391bffb9cfff80ac238c886ef0a461,	
	128'hb8d2a67df5a999fdbf93edd0343296c9,	
	128'haaca7367396b69a221bd632bea386eec,	
	128'ha80fd5020dfe65f5f16293ec92c6fd89,	
	128'h2162995b8217a67f1abc342e146406f8,	
	128'hc6a6164b7a60bae4e986ffac28dfadd9,	
	128'h64e0d7f900e3d9c83e4b8f96717b2146,	
	128'h1ad2561de8c1232f5d8dbab4739b6cbb,	
	128'h279689e9a557f58b1c3bf40c97a90964,	
	128'hc4637e4a5e6377f9cc5a8638045de029,	
	128'h492e607e5aea4688594b45f3aee3df90,	
	128'he8c4e4381feec74054954c05b777a00a,
	128'h91549514605f38246c9b724ad839f01d,
    128'h74b24e3b6fefe40a4f9ef7ac6e44d76a,
	128'h2437a683dc5d4b52abb4a123a8df86c6,
	128'hbb2852c891c5947d2ed44032c421b85f,
	128'h1b9f5fbd5e8a4264c0a85b80409afa5e,
	128'h30dab809f85a917fe924733f424ac589,
	128'heaef5c1f8d605192646695ceadc65f32,
	128'hb8aa90040b4c15a12316b78e0f9586fc,
	128'h97fac8297ceaabc87d454350601e0673,
	128'h9b47ef567ac28dfe488492f157e2b2e0,
	128'h1b8426027ddb962b5c5ba7eb8bc9ab63,
	128'he917fc77e71992a12dbe4c18068bec82,
	128'hdceebbc98840f8ae6daf76573b7e56f4,
	128'h4e11a9f74205125b61e0aee047eca20d,
	128'hf60467f55a1f17eab88e800120cbc284,
	128'hd436649f600b449ee276530f0cd83c11,
	128'h3bc0e3656a9e3ac7cd378a737f53b637,
	128'h6bacae63d33b928aa8380f8d54d88c17,
	128'h8935ffbc75ae6251bf8e859f085adcb9,
	128'h93dc4970fe35f67747cb0562c06d875a,
	128'h14f9df858975851797ba604fb0d16cc7,
	128'h02ea0c98dca10b38c21b3b14e8d1b71f,
	128'h8f091b1b5b0749b2adc803e63dda9b72,
	128'h05b389e3322c6da08384345a4137fd08,
	128'h381308c438f35b399f10ad71b05027d8,
	128'h68c230fcfa9279c3409fc423e2acbe04,
	128'h1c84a475acb011f3f59f4f46b76274c0,
	128'h45119b68cb3f8399ee60066b5611a4d7,
	128'h9423762f527a4060ffca312dcca22a16,
	128'hf361a2745a33f056a5ac6ace2f08e344,
	128'h5ef145766eca849f5d011536a6557fdb,
	128'hc9af27b2c89c9b4cf4a0c4106ac80318,
	128'hfb9c4f16c621f4eab7e9ac1d7551dd57,
	128'h138e06fba466fa70854d8c2e524cffb2,
	128'hfb4bc78b225070773f04c40466d4e90c,
	128'h8b2cbff1ed0150feda8a4799be94551f,
	128'h08b30d7b3f27962709a36bcadfb974bd,
	128'hfdf6d32e044d77adcf37fb97ac213326,
	128'h93cb284ecdcfd781a8afe32077949e88,
	128'h7b017bb02ec87b2b94c96e40a26fc71a,
	128'hc5c038b6990664ab08a3aaa5df9f3266,
	128'h4b7020be37fab6259b2a27f4ec551576,
	128'h60136703374f64e860b48ce31f930716,
	128'h8d63a269b14d506ccc401ab8a9f1b591,
	128'hd317f81dc6aa454aee4bd4a5a5cff4bd,
	128'hdddececd5354f04d530d76ed884246eb,
	128'h41c5205cc8fd8eda9a3cffd2518f365a,
	128'hcf42fb474293d96eca9db1b37b1ba676,
	128'ha231692607169b4ecdead5cd3b10db3e,
	128'hace4b91c9c669e77e7acacd19859ed49,
	128'h75db7cfd4a7b2b62ab78a48f3ddaf4af,
	128'hc1faba2d46e259cf480d7c38e4572a58,
	128'h241c45bc6ae16dee6eb7bea128701582,
	128'h8fd03057cf1364420c2b78069a3e2502,
	128'hddb505e6cc1384cbaec1df90b80beb20,
	128'h5674a3bed27bf4bd3622f9f5fe208306,
	128'hb687f26a89cfbfbb8e5eeac54055315e,
	128'h0547dd32d3b29ab6a4caeb606c5b6f78,
	128'h186861f8bc5386d31fb77f720c3226e6,
	128'heacf1e6c4224efb38900b185ab1dfd42,
	128'hd241aab05a42d319de81d874f5c7b90d,
	128'h5eb9bc759e2ad8d2140a6c762ae9e1ab,
	128'h018596e15e78e2c064159defce5f3085,
	128'hdd8a493514231cbf56eccee4c40889fb
	};
	
	//--------------------------------------------------------
	//
	// 256-bit decryption test vectors
	//
	//--------------------------------------------------------
	
		
	// FIPS-197 appendix C.3 Sample Vector 256-bit
	`define FIPS197_256_VEC_SIZE 1
	logic	[0:255]	FIPS197_256_kt[`FIPS197_256_VEC_SIZE] = {256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f};
	logic	[0:127]	FIPS197_256_pt[`FIPS197_256_VEC_SIZE] = {128'h00112233445566778899aabbccddeeff};
	logic	[0:127]	FIPS197_256_ct[`FIPS197_256_VEC_SIZE] = {128'h8ea2b7ca516745bfeafc49904b496089};
	
	// ECB-AES256.Decrypt sample vector test
	// SP800-38a appendix F.1.6
	`define ECB_DECRYPT_256_VEC_SIZE 4
	int	ECBDecrypt_256_failed = 0;
	logic	[0:255]	ECBDecrypt_256_kt = 256'h603deb1015ca71be2b73aef0857d77811f352c073b6108d72d9810a30914dff4;	
	logic	[0:127]	ECBDecrypt_256_ct [`ECB_DECRYPT_256_VEC_SIZE] = {
	128'hf3eed1bdb5d2a03c064b5a7e3db181f8,
	128'h591ccb10d410ed26dc5ba74a31362870,
	128'hb6ed21b99ca6f4f9f153e7b1beafed1d,
	128'h23304b7a39f9f3ff067d8d8f9e24ecc7
	};
	
	logic	[0:127]	ECBDecrypt_256_pt [`ECB_DECRYPT_256_VEC_SIZE] = {
	128'h6bc1bee22e409f96e93d7e117393172a,
	128'hae2d8a571e03ac9c9eb76fac45af8e51,
	128'h30c81c46a35ce411e5fbc1191a0a52ef,
	128'hf69f2445df4f9b17ad2b417be66c3710
	};
	
	// 256-bit GFSbox Known Answer Test vectors.
	// AESAVS appendix B.2
	`define GFSbox_256_VEC_SIZE 5
	int	GFSbox_256_failed=0;
	logic	[0:255]	GFSbox_256_kt = 'h0;
	logic	[0:127]	GFSbox_256_ct[`GFSbox_256_VEC_SIZE] = {
	128'h5c9d844ed46f9885085e5d6a4f94c7d7,
    128'ha9ff75bd7cf6613d3731c77c3b6d0c04,
    128'h623a52fcea5d443e48d9181ab32c7421,
    128'h38f2c7ae10612415d27ca190d27da8b4,
    128'h1bc704f1bce135ceb810341b216d7abe
	};
										
	logic	[0:127]	GFSbox_256_pt[`GFSbox_256_VEC_SIZE] = {
	128'h014730f80ac625fe84f026c60bfd547d,
	128'h0b24af36193ce4665f2825d7b4749c98,
	128'h761c1fe41a18acf20d241650611d90f1,
	128'h8a560769d605868ad80d819bdba03771,
	128'h91fbef2d15a97816060bee1feaa49afe
	};
	
	// 256-bit KeySBox Known Answer Test vectors
	// AESAVS appendix C.2
	`define KEYSBOX_256_VEC_SIZE 16
	int	KeySbox_256_failed = 0;
	logic	[0:127]	KeySbox_256_pt = 'h0;
	logic	[0:127]	KeySbox_256_ct[`KEYSBOX_256_VEC_SIZE] = {
	128'h46f2fb342d6f0ab477476fc501242c5f,
    128'h4bf3b0a69aeb6657794f2901b1440ad4,
    128'h352065272169abf9856843927d0674fd,
    128'h4307456a9e67813b452e15fa8fffe398,
    128'h4663446607354989477a5c6f0f007ef4,
    128'h531c2c38344578b84d50b3c917bbb6e1,
    128'hfc6aec906323480005c58e7e1ab004ad,
    128'ha3944b95ca0b52043584ef02151926a8,
    128'ha74289fe73a4c123ca189ea1e1b49ad5,
    128'hb91d4ea4488644b56cf0812fa7fcf5fc,
    128'h304f81ab61a80c2e743b94d5002a126b,
    128'h649a71545378c783e368c9ade7114f6c,
    128'h47cb030da2ab051dfc6c4bf6910d12bb,
	128'h798c7c005dee432b2c8ea5dfa381ecc3,
	128'h637c31dc2591a07636f646b72daabbe7,
	128'h179a49c712154bbffbe6e7a84a18e220
	};
									
	logic	[0:255]	KeySbox_256_kt[`KEYSBOX_256_VEC_SIZE] = {
	256'hc47b0294dbbbee0fec4757f22ffeee3587ca4730c3d33b691df38bab076bc558,
    256'h28d46cffa158533194214a91e712fc2b45b518076675affd910edeca5f41ac64,
    256'hc1cc358b449909a19436cfbb3f852ef8bcb5ed12ac7058325f56e6099aab1a1c,
    256'h984ca75f4ee8d706f46c2d98c0bf4a45f5b00d791c2dfeb191b5ed8e420fd627,
    256'hb43d08a447ac8609baadae4ff12918b9f68fc1653f1269222f123981ded7a92f,
    256'h1d85a181b54cde51f0e098095b2962fdc93b51fe9b88602b3f54130bf76a5bd9,
    256'hdc0eba1f2232a7879ded34ed8428eeb8769b056bbaf8ad77cb65c3541430b4cf,
    256'hf8be9ba615c5a952cabbca24f68f8593039624d524c816acda2c9183bd917cb9,
    256'h797f8b3d176dac5b7e34a2d539c4ef367a16f8635f6264737591c5c07bf57a3e,
    256'h6838d40caf927749c13f0329d331f448e202c73ef52c5f73a37ca635d4c47707,
    256'hccd1bc3c659cd3c59bc437484e3c5c724441da8d6e90ce556cd57d0752663bbc,
    256'h13428b5e4c005e0636dd338405d173ab135dec2a25c22c5df0722d69dcc43887,
    256'h07eb03a08d291d1b07408bf3512ab40c91097ac77461aad4bb859647f74f00ee,
	256'h90143ae20cd78c5d8ebdd6cb9dc1762427a96c78c639bccc41a61424564eafe1,
	256'hb7a5794d52737475d53d5a377200849be0260a67a2b22ced8bbef12882270d07,
	256'hfca02f3d5011cfc5c1e23165d413a049d4526a991827424d896fe3435e0bf68e
	};

	// 256-bit VarTxt Known Answer Test vectors
	// AESAVS appendix D.3
	`define VARTXT_256_VEC_SIZE 128
	int	VarTxt_256_failed = 0;
	logic	[0:255]	VarTxt_256_kt = 'h0;
	logic	[0:127]	VarTxt_256_pt[`VARTXT_256_VEC_SIZE] = {
	128'h80000000000000000000000000000000, 
	128'hc0000000000000000000000000000000, 
	128'he0000000000000000000000000000000, 
	128'hf0000000000000000000000000000000, 
	128'hf8000000000000000000000000000000, 
	128'hfc000000000000000000000000000000, 
	128'hfe000000000000000000000000000000, 
	128'hff000000000000000000000000000000, 
	128'hff800000000000000000000000000000, 
	128'hffc00000000000000000000000000000, 
	128'hffe00000000000000000000000000000, 
	128'hfff00000000000000000000000000000, 
	128'hfff80000000000000000000000000000, 
	128'hfffc0000000000000000000000000000, 
	128'hfffe0000000000000000000000000000, 
	128'hffff0000000000000000000000000000, 
	128'hffff8000000000000000000000000000, 
	128'hffffc000000000000000000000000000, 
	128'hffffe000000000000000000000000000, 
	128'hfffff000000000000000000000000000, 
	128'hfffff800000000000000000000000000, 
	128'hfffffc00000000000000000000000000, 
	128'hfffffe00000000000000000000000000, 
	128'hffffff00000000000000000000000000, 
	128'hffffff80000000000000000000000000, 
	128'hffffffc0000000000000000000000000, 
	128'hffffffe0000000000000000000000000, 
	128'hfffffff0000000000000000000000000, 
	128'hfffffff8000000000000000000000000, 
	128'hfffffffc000000000000000000000000, 
	128'hfffffffe000000000000000000000000, 
	128'hffffffff000000000000000000000000, 
	128'hffffffff800000000000000000000000, 
	128'hffffffffc00000000000000000000000, 
	128'hffffffffe00000000000000000000000, 
	128'hfffffffff00000000000000000000000, 
	128'hfffffffff80000000000000000000000, 
	128'hfffffffffc0000000000000000000000, 
	128'hfffffffffe0000000000000000000000, 
	128'hffffffffff0000000000000000000000, 
	128'hffffffffff8000000000000000000000, 
	128'hffffffffffc000000000000000000000, 
	128'hffffffffffe000000000000000000000, 
	128'hfffffffffff000000000000000000000, 
	128'hfffffffffff800000000000000000000, 
	128'hfffffffffffc00000000000000000000, 
	128'hfffffffffffe00000000000000000000, 
	128'hffffffffffff00000000000000000000, 
	128'hffffffffffff80000000000000000000, 
	128'hffffffffffffc0000000000000000000, 
	128'hffffffffffffe0000000000000000000, 
	128'hfffffffffffff0000000000000000000, 
	128'hfffffffffffff8000000000000000000, 
	128'hfffffffffffffc000000000000000000, 
	128'hfffffffffffffe000000000000000000, 
	128'hffffffffffffff000000000000000000, 
	128'hffffffffffffff800000000000000000, 
	128'hffffffffffffffc00000000000000000, 
	128'hffffffffffffffe00000000000000000, 
	128'hfffffffffffffff00000000000000000, 
	128'hfffffffffffffff80000000000000000, 
	128'hfffffffffffffffc0000000000000000, 
	128'hfffffffffffffffe0000000000000000, 
	128'hffffffffffffffff0000000000000000, 
	128'hffffffffffffffff8000000000000000, 
	128'hffffffffffffffffc000000000000000, 
	128'hffffffffffffffffe000000000000000, 
	128'hfffffffffffffffff000000000000000, 
	128'hfffffffffffffffff800000000000000, 
	128'hfffffffffffffffffc00000000000000, 
	128'hfffffffffffffffffe00000000000000, 
	128'hffffffffffffffffff00000000000000, 
	128'hffffffffffffffffff80000000000000, 
	128'hffffffffffffffffffc0000000000000, 
	128'hffffffffffffffffffe0000000000000, 
	128'hfffffffffffffffffff0000000000000, 
	128'hfffffffffffffffffff8000000000000, 
	128'hfffffffffffffffffffc000000000000, 
	128'hfffffffffffffffffffe000000000000, 
	128'hffffffffffffffffffff000000000000, 
	128'hffffffffffffffffffff800000000000, 
	128'hffffffffffffffffffffc00000000000, 
	128'hffffffffffffffffffffe00000000000, 
	128'hfffffffffffffffffffff00000000000, 
	128'hfffffffffffffffffffff80000000000, 
	128'hfffffffffffffffffffffc0000000000, 
	128'hfffffffffffffffffffffe0000000000, 
	128'hffffffffffffffffffffff0000000000, 
	128'hffffffffffffffffffffff8000000000, 
	128'hffffffffffffffffffffffc000000000, 
	128'hffffffffffffffffffffffe000000000, 
	128'hfffffffffffffffffffffff000000000, 
	128'hfffffffffffffffffffffff800000000, 
	128'hfffffffffffffffffffffffc00000000, 
	128'hfffffffffffffffffffffffe00000000, 
	128'hffffffffffffffffffffffff00000000, 
	128'hffffffffffffffffffffffff80000000, 
	128'hffffffffffffffffffffffffc0000000, 
	128'hffffffffffffffffffffffffe0000000, 
	128'hfffffffffffffffffffffffff0000000, 
	128'hfffffffffffffffffffffffff8000000, 
	128'hfffffffffffffffffffffffffc000000, 
	128'hfffffffffffffffffffffffffe000000, 
	128'hffffffffffffffffffffffffff000000, 
	128'hffffffffffffffffffffffffff800000, 
	128'hffffffffffffffffffffffffffc00000, 
	128'hffffffffffffffffffffffffffe00000, 
	128'hfffffffffffffffffffffffffff00000, 
	128'hfffffffffffffffffffffffffff80000, 
	128'hfffffffffffffffffffffffffffc0000, 
	128'hfffffffffffffffffffffffffffe0000, 
	128'hffffffffffffffffffffffffffff0000, 
	128'hffffffffffffffffffffffffffff8000, 
	128'hffffffffffffffffffffffffffffc000, 
	128'hffffffffffffffffffffffffffffe000, 
	128'hfffffffffffffffffffffffffffff000, 
	128'hfffffffffffffffffffffffffffff800, 
	128'hfffffffffffffffffffffffffffffc00, 
	128'hfffffffffffffffffffffffffffffe00, 
	128'hffffffffffffffffffffffffffffff00, 
	128'hffffffffffffffffffffffffffffff80, 
	128'hffffffffffffffffffffffffffffffc0, 
	128'hffffffffffffffffffffffffffffffe0, 
	128'hfffffffffffffffffffffffffffffff0, 
	128'hfffffffffffffffffffffffffffffff8, 
	128'hfffffffffffffffffffffffffffffffc, 
	128'hfffffffffffffffffffffffffffffffe, 
	128'hffffffffffffffffffffffffffffffff
	}; 
	
	logic	[0:127]	VarTxt_256_ct[`VARTXT_256_VEC_SIZE] = {
	128'hddc6bf790c15760d8d9aeb6f9a75fd4e,
	128'h0a6bdc6d4c1e6280301fd8e97ddbe601,
	128'h9b80eefb7ebe2d2b16247aa0efc72f5d,
	128'h7f2c5ece07a98d8bee13c51177395ff7,
	128'h7818d800dcf6f4be1e0e94f403d1e4c2,
	128'he74cd1c92f0919c35a0324123d6177d3,
	128'h8092a4dcf2da7e77e93bdd371dfed82e,
	128'h49af6b372135acef10132e548f217b17,
	128'h8bcd40f94ebb63b9f7909676e667f1e7,
	128'hfe1cffb83f45dcfb38b29be438dbd3ab,
	128'h0dc58a8d886623705aec15cb1e70dc0e,
	128'hc218faa16056bd0774c3e8d79c35a5e4,
	128'h047bba83f7aa841731504e012208fc9e,
	128'hdc8f0e4915fd81ba70a331310882f6da,
	128'h1569859ea6b7206c30bf4fd0cbfac33c,
	128'h300ade92f88f48fa2df730ec16ef44cd,
	128'h1fe6cc3c05965dc08eb0590c95ac71d0,
	128'h59e858eaaa97fec38111275b6cf5abc0,
	128'h2239455e7afe3b0616100288cc5a723b,
	128'h3ee500c5c8d63479717163e55c5c4522,
	128'hd5e38bf15f16d90e3e214041d774daa8,
	128'hb1f4066e6f4f187dfe5f2ad1b17819d0,
	128'h6ef4cc4de49b11065d7af2909854794a,
	128'hac86bc606b6640c309e782f232bf367f,
	128'h36aff0ef7bf3280772cf4cac80a0d2b2,
	128'h1f8eedea0f62a1406d58cfc3ecea72cf,
	128'habf4154a3375a1d3e6b1d454438f95a6,
	128'h96f96e9d607f6615fc192061ee648b07,
	128'hcf37cdaaa0d2d536c71857634c792064,
	128'hfbd6640c80245c2b805373f130703127,
	128'h8d6a8afe55a6e481badae0d146f436db,
	128'h6a4981f2915e3e68af6c22385dd06756,
	128'h42a1136e5f8d8d21d3101998642d573b,
	128'h9b471596dc69ae1586cee6158b0b0181,
	128'h753665c4af1eff33aa8b628bf8741cfd,
	128'h9a682acf40be01f5b2a4193c9a82404d,
	128'h54fafe26e4287f17d1935f87eb9ade01,
	128'h49d541b2e74cfe73e6a8e8225f7bd449,
	128'h11a45530f624ff6f76a1b3826626ff7b,
	128'hf96b0c4a8bc6c86130289f60b43b8fba,
	128'h48c7d0e80834ebdc35b6735f76b46c8b,
	128'h2463531ab54d66955e73edc4cb8eaa45,
	128'hac9bd8e2530469134b9d5b065d4f565b,
	128'h3f5f9106d0e52f973d4890e6f37e8a00,
	128'h20ebc86f1304d272e2e207e59db639f0,
	128'he67ae6426bf9526c972cff072b52252c,
	128'h1a518dddaf9efa0d002cc58d107edfc8,
	128'head731af4d3a2fe3b34bed047942a49f,
	128'hb1d4efe40242f83e93b6c8d7efb5eae9,
	128'hcd2b1fec11fd906c5c7630099443610a,
	128'ha1853fe47fe29289d153161d06387d21,
	128'h4632154179a555c17ea604d0889fab14,
	128'hdd27cac6401a022e8f38f9f93e774417,
	128'hc090313eb98674f35f3123385fb95d4d,
	128'hcc3526262b92f02edce548f716b9f45c,
	128'hc0838d1a2b16a7c7f0dfcc433c399c33,
	128'h0d9ac756eb297695eed4d382eb126d26,
	128'h56ede9dda3f6f141bff1757fa689c3e1,
	128'h768f520efe0f23e61d3ec8ad9ce91774,
	128'hb1144ddfa75755213390e7c596660490,
	128'h1d7c0c4040b355b9d107a99325e3b050,
	128'hd8e2bb1ae8ee3dcf5bf7d6c38da82a1a,
	128'hfaf82d178af25a9886a47e7f789b98d7,
	128'h9b58dbfd77fe5aca9cfc190cd1b82d19,
	128'h77f392089042e478ac16c0c86a0b5db5,
	128'h19f08e3420ee69b477ca1420281c4782,
	128'ha1b19beee4e117139f74b3c53fdcb875,
	128'ha37a5869b218a9f3a0868d19aea0ad6a,
	128'hbc3594e865bcd0261b13202731f33580,
	128'h811441ce1d309eee7185e8c752c07557,
	128'h959971ce4134190563518e700b9874d1,
	128'h76b5614a042707c98e2132e2e805fe63,
	128'h7d9fa6a57530d0f036fec31c230b0cc6,
	128'h964153a83bf6989a4ba80daa91c3e081,
	128'ha013014d4ce8054cf2591d06f6f2f176,
	128'hd1c5f6399bf382502e385eee1474a869,
	128'h0007e20b8298ec354f0f5fe7470f36bd,
	128'hb95ba05b332da61ef63a2b31fcad9879,
	128'h4620a49bd967491561669ab25dce45f4,
	128'h12e71214ae8e04f0bb63d7425c6f14d5,
	128'h4cc42fc1407b008fe350907c092e80ac,
	128'h08b244ce7cbc8ee97fbba808cb146fda,
	128'h39b333e8694f21546ad1edd9d87ed95b,
	128'h3b271f8ab2e6e4a20ba8090f43ba78f3,
	128'h9ad983f3bf651cd0393f0a73cccdea50,
	128'h8f476cbff75c1f725ce18e4bbcd19b32,
	128'h905b6267f1d6ab5320835a133f096f2a,
	128'h145b60d6d0193c23f4221848a892d61a,
	128'h55cfb3fb6d75cad0445bbc8dafa25b0f,
	128'h7b8e7098e357ef71237d46d8b075b0f5,
	128'h2bf27229901eb40f2df9d8398d1505ae,
	128'h83a63402a77f9ad5c1e931a931ecd706,
	128'h6f8ba6521152d31f2bada1843e26b973,
	128'he5c3b8e30fd2d8e6239b17b44bd23bbd,
	128'h1ac1f7102c59933e8b2ddc3f14e94baa,
	128'h21d9ba49f276b45f11af8fc71a088e3d,
	128'h649f1cddc3792b4638635a392bc9bade,
	128'he2775e4b59c1bc2e31a2078c11b5a08c,
	128'h2be1fae5048a25582a679ca10905eb80,
	128'hda86f292c6f41ea34fb2068df75ecc29,
	128'h220df19f85d69b1b562fa69a3c5beca5,
	128'h1f11d5d0355e0b556ccdb6c7f5083b4d,
	128'h62526b78be79cb384633c91f83b4151b,
	128'h90ddbcb950843592dd47bbef00fdc876,
	128'h2fd0e41c5b8402277354a7391d2618e2,
	128'h3cdf13e72dee4c581bafec70b85f9660,
	128'hafa2ffc137577092e2b654fa199d2c43,
	128'h8d683ee63e60d208e343ce48dbc44cac,
	128'h705a4ef8ba2133729c20185c3d3a4763,
	128'h0861a861c3db4e94194211b77ed761b9,
	128'h4b00c27e8b26da7eab9d3a88dec8b031,
	128'h5f397bf03084820cc8810d52e5b666e9,
	128'h63fafabb72c07bfbd3ddc9b1203104b8,
	128'h683e2140585b18452dd4ffbb93c95df9,
	128'h286894e48e537f8763b56707d7d155c8,
	128'ha423deabc173dcf7e2c4c53e77d37cd1,
	128'heb8168313e1cfdfdb5e986d5429cf172,
	128'h27127daafc9accd2fb334ec3eba52323,
	128'hee0715b96f72e3f7a22a5064fc592f4c,
	128'h29ee526770f2a11dcfa989d1ce88830f,
	128'h0493370e054b09871130fe49af730a5a,
	128'h9b7b940f6c509f9e44a4ee140448ee46,
	128'h2915be4a1ecfdcbe3e023811a12bb6c7,
	128'h7240e524bc51d8c4d440b1be55d1062c,
	128'hda63039d38cb4612b2dc36ba26684b93,
	128'h0f59cb5a4b522e2ac56c1a64f558ad9a,
	128'h7bfe9d876c6d63c1d035da8fe21c409d,
	128'hacdace8078a32b1a182bfa4987ca1347
	};
	
	// 256-bit VarKey Known Answer Test
	// AESAVS appendix E.2
	`define VARKEY_256_VEC_SIZE 256
	int	VarKey_256_failed = 0;
	logic	[0:127]	VarKey_256_pt = 'h0;
	logic	[0:255]	VarKey_256_kt[`VARKEY_256_VEC_SIZE] = {
	256'h8000000000000000000000000000000000000000000000000000000000000000,	
	256'hc000000000000000000000000000000000000000000000000000000000000000,	
	256'he000000000000000000000000000000000000000000000000000000000000000,	
	256'hf000000000000000000000000000000000000000000000000000000000000000,	
	256'hf800000000000000000000000000000000000000000000000000000000000000,	
	256'hfc00000000000000000000000000000000000000000000000000000000000000,	
	256'hfe00000000000000000000000000000000000000000000000000000000000000,	
	256'hff00000000000000000000000000000000000000000000000000000000000000,	
	256'hff80000000000000000000000000000000000000000000000000000000000000,	
	256'hffc0000000000000000000000000000000000000000000000000000000000000,	
	256'hffe0000000000000000000000000000000000000000000000000000000000000,	
	256'hfff0000000000000000000000000000000000000000000000000000000000000,	
	256'hfff8000000000000000000000000000000000000000000000000000000000000,	
	256'hfffc000000000000000000000000000000000000000000000000000000000000,	
	256'hfffe000000000000000000000000000000000000000000000000000000000000,	
	256'hffff000000000000000000000000000000000000000000000000000000000000,	
	256'hffff800000000000000000000000000000000000000000000000000000000000,	
	256'hffffc00000000000000000000000000000000000000000000000000000000000,	
	256'hffffe00000000000000000000000000000000000000000000000000000000000,	
	256'hfffff00000000000000000000000000000000000000000000000000000000000,	
	256'hfffff80000000000000000000000000000000000000000000000000000000000,	
	256'hfffffc0000000000000000000000000000000000000000000000000000000000,	
	256'hfffffe0000000000000000000000000000000000000000000000000000000000,	
	256'hffffff0000000000000000000000000000000000000000000000000000000000,	
	256'hffffff8000000000000000000000000000000000000000000000000000000000,	
	256'hffffffc000000000000000000000000000000000000000000000000000000000,	
	256'hffffffe000000000000000000000000000000000000000000000000000000000,	
	256'hfffffff000000000000000000000000000000000000000000000000000000000,	
	256'hfffffff800000000000000000000000000000000000000000000000000000000,	
	256'hfffffffc00000000000000000000000000000000000000000000000000000000,	
	256'hfffffffe00000000000000000000000000000000000000000000000000000000,	
	256'hffffffff00000000000000000000000000000000000000000000000000000000,	
	256'hffffffff80000000000000000000000000000000000000000000000000000000,	
	256'hffffffffc0000000000000000000000000000000000000000000000000000000,	
	256'hffffffffe0000000000000000000000000000000000000000000000000000000,	
	256'hfffffffff0000000000000000000000000000000000000000000000000000000,	
	256'hfffffffff8000000000000000000000000000000000000000000000000000000,	
	256'hfffffffffc000000000000000000000000000000000000000000000000000000,	
	256'hfffffffffe000000000000000000000000000000000000000000000000000000,	
	256'hffffffffff000000000000000000000000000000000000000000000000000000,	
	256'hffffffffff800000000000000000000000000000000000000000000000000000,	
	256'hffffffffffc00000000000000000000000000000000000000000000000000000,	
	256'hffffffffffe00000000000000000000000000000000000000000000000000000,	
	256'hfffffffffff00000000000000000000000000000000000000000000000000000,	
	256'hfffffffffff80000000000000000000000000000000000000000000000000000,	
	256'hfffffffffffc0000000000000000000000000000000000000000000000000000,	
	256'hfffffffffffe0000000000000000000000000000000000000000000000000000,	
	256'hffffffffffff0000000000000000000000000000000000000000000000000000,	
	256'hffffffffffff8000000000000000000000000000000000000000000000000000,	
	256'hffffffffffffc000000000000000000000000000000000000000000000000000,	
	256'hffffffffffffe000000000000000000000000000000000000000000000000000,	
	256'hfffffffffffff000000000000000000000000000000000000000000000000000,	
	256'hfffffffffffff800000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffc00000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffe00000000000000000000000000000000000000000000000000,	
	256'hffffffffffffff00000000000000000000000000000000000000000000000000,	
	256'hffffffffffffff80000000000000000000000000000000000000000000000000,	
	256'hffffffffffffffc0000000000000000000000000000000000000000000000000,	
	256'hffffffffffffffe0000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffff0000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffff8000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffc000000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffe000000000000000000000000000000000000000000000000,	
	256'hffffffffffffffff000000000000000000000000000000000000000000000000,	
	256'hffffffffffffffff800000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffc00000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffe00000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffff00000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffff80000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffc0000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffe0000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffff0000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffff8000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffc000000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffe000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffff000000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffff800000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffc00000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffe00000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffff00000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffff80000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffc0000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffe0000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffff0000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffff8000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffc000000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffe000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffff000000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffff800000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffc00000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffe00000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffff00000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffff80000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffc0000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffe0000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffff0000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffff8000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffc000000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffe000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffff000000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffff800000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffc00000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffe00000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffff00000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffff80000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffc0000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffe0000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffff0000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffff8000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffc000000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffe000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffff000000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffff800000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffc00000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffe00000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffff00000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffff80000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffc0000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffe0000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffff0000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffff8000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffffc000000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffffe000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffff000000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffff800000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffffc00000000000000000000000000000000,	
	256'hfffffffffffffffffffffffffffffffe00000000000000000000000000000000,	
	256'hffffffffffffffffffffffffffffffff00000000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffff80000000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffc0000000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffe0000000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffff0000000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffff8000000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffc000000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffe000000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffff000000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffff800000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffc00000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffe00000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffff00000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffff80000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffc0000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffe0000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffff0000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffff8000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffc000000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffe000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffff000000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffff800000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffc00000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffe00000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffff00000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffff80000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffc0000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffe0000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffff0000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffff8000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffc000000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffe000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffff000000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffff800000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffc00000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffe00000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffff00000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffff80000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffc0000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffe0000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffff0000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffff8000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffc000000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffe000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffff000000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffff800000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffc00000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffe00000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffff00000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffff80000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffc0000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffe0000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffff0000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffff8000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffc000000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffe000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffff000000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffff800000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffc00000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffe00000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffff00000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffff80000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffc0000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffe0000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffc000000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffe000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffff000000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffff800000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffc00000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffe00000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffff00000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffff80000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffc0000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffe0000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffc000000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffe000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffff800000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffff00000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffff80000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffc0000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffe0000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffff800000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc000,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff800,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc00,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe00,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff00,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff80,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc0,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe0,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff0,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff8,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc,
	256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe,
	256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
	};                                   
	
	logic	[0:127]	VarKey_256_ct[`VARKEY_256_VEC_SIZE] = {
	128'he35a6dcb19b201a01ebcfa8aa22b5759,
	128'hb29169cdcf2d83e838125a12ee6aa400,
	128'hd8f3a72fc3cdf74dfaf6c3e6b97b2fa6,
	128'h1c777679d50037c79491a94da76a9a35,
	128'h9cf4893ecafa0a0247a898e040691559,
	128'h8fbb413703735326310a269bd3aa94b2,
	128'h60e32246bed2b0e859e55c1cc6b26502,
	128'hec52a212f80a09df6317021bc2a9819e,
	128'hf23e5b600eb70dbccf6c0b1d9a68182c,
	128'ha3f599d63a82a968c33fe26590745970,
	128'hd1ccb9b1337002cbac42c520b5d67722,
	128'hcc111f6c37cf40a1159d00fb59fb0488,
	128'hdc43b51ab609052372989a26e9cdd714,
	128'h4dcede8da9e2578f39703d4433dc6459,
	128'h1a4c1c263bbccfafc11782894685e3a8,
	128'h937ad84880db50613423d6d527a2823d,
	128'h610b71dfc688e150d8152c5b35ebc14d,
	128'h27ef2495dabf323885aab39c80f18d8b,
	128'h633cafea395bc03adae3a1e2068e4b4e,
	128'h6e1b482b53761cf631819b749a6f3724,
	128'h976e6f851ab52c771998dbb2d71c75a9,
	128'h85f2ba84f8c307cf525e124c3e22e6cc,
	128'h6bcca98bf6a835fa64955f72de4115fe,
	128'h2c75e2d36eebd65411f14fd0eb1d2a06,
	128'hbd49295006250ffca5100b6007a0eade,
	128'ha190527d0ef7c70f459cd3940df316ec,
	128'hbbd1097a62433f79449fa97d4ee80dbf,
	128'h07058e408f5b99b0e0f061a1761b5b3b,
	128'h5fd1f13fa0f31e37fabde328f894eac2,
	128'hfc4af7c948df26e2ef3e01c1ee5b8f6f,
	128'h829fd7208fb92d44a074a677ee9861ac,
	128'had9fc613a703251b54c64a0e76431711,
	128'h33ac9eccc4cc75e2711618f80b1548e8,
	128'h2025c74b8ad8f4cda17ee2049c4c902d,
	128'hf85ca05fe528f1ce9b790166e8d551e7,
	128'h6f6238d8966048d4967154e0dad5a6c9,
	128'hf2b21b4e7640a9b3346de8b82fb41e49,
	128'hf836f251ad1d11d49dc344628b1884e1,
	128'h077e9470ae7abea5a9769d49182628c3,
	128'he0dcc2d27fc9865633f85223cf0d611f,
	128'hbe66cfea2fecd6bf0ec7b4352c99bcaa,
	128'hdf31144f87a2ef523facdcf21a427804,
	128'hb5bb0f5629fb6aae5e1839a3c3625d63,
	128'h3c9db3335306fe1ec612bdbfae6b6028,
	128'h3dd5c34634a79d3cfcc8339760e6f5f4,
	128'h82bda118a3ed7af314fa2ccc5c07b761,
	128'h2937a64f7d4f46fe6fea3b349ec78e38,
	128'h225f068c28476605735ad671bb8f39f3,
	128'hae682c5ecd71898e08942ac9aa89875c,
	128'h5e031cb9d676c3022d7f26227e85c38f,
	128'ha78463fb064db5d52bb64bfef64f2dda,
	128'h8aa9b75e784593876c53a00eae5af52b,
	128'h3f84566df23da48af692722fe980573a,
	128'h31690b5ed41c7eb42a1e83270a7ff0e6,
	128'h77dd7702646d55f08365e477d3590eda,
	128'h4c022ac62b3cb78d739cc67b3e20bb7e,
	128'h092fa137ce18b5dfe7906f550bb13370,
	128'h3e0cdadf2e68353c0027672c97144dd3,
	128'hd8c4b200b383fc1f2b2ea677618a1d27,
	128'h11825f99b0e9bb3477c1c0713b015aac,
	128'hf8b9fffb5c187f7ddc7ab10f4fb77576,
	128'hffb4e87a32b37d6f2c8328d3b5377802,
	128'hd276c13a5d220f4da9224e74896391ce,
	128'h94efe7a0e2e031e2536da01df799c927,
	128'h8f8fd822680a85974e53a5a8eb9d38de,
	128'he0f0a91b2e45f8cc37b7805a3042588d,
	128'h597a6252255e46d6364dbeeda31e279c,
	128'hf51a0f694442b8f05571797fec7ee8bf,
	128'h9ff071b165b5198a93dddeebc54d09b5,
	128'hc20a19fd5758b0c4bc1a5df89cf73877,
	128'h97120166307119ca2280e9315668e96f,
	128'h4b3b9f1e099c2a09dc091e90e4f18f0a,
	128'heb040b891d4b37f6851f7ec219cd3f6d,
	128'h9f0fdec08b7fd79aa39535bea42db92a,
	128'h2e70f168fc74bf911df240bcd2cef236,
	128'h462ccd7f5fd1108dbc152f3cacad328b,
	128'ha4af534a7d0b643a01868785d86dfb95,
	128'hab980296197e1a5022326c31da4bf6f3,
	128'hf97d57b3333b6281b07d486db2d4e20c,
	128'hf33fa36720231afe4c759ade6bd62eb6,
	128'hfdcfac0c02ca538343c68117e0a15938,
	128'had4916f5ee5772be764fc027b8a6e539,
	128'h2e16873e1678610d7e14c02d002ea845,
	128'h4e6e627c1acc51340053a8236d579576,
	128'hab0c8410aeeead92feec1eb430d652cb,
	128'he86f7e23e835e114977f60e1a592202e,
	128'he68ad5055a367041fade09d9a70a794b,
	128'h0791823a3c666bb6162825e78606a7fe,
	128'hdcca366a9bf47b7b868b77e25c18a364,
	128'h684c9efc237e4a442965f84bce20247a,
	128'ha858411ffbe63fdb9c8aa1bfaed67b52,
	128'h04bc3da2179c3015498b0e03910db5b8,
	128'h40071eeab3f935dbc25d00841460260f,
	128'h0ebd7c30ed2016e08ba806ddb008bcc8,
	128'h15c6becf0f4cec7129cbd22d1a79b1b8,
	128'h0aeede5b91f721700e9e62edbf60b781,
	128'h266581af0dcfbed1585e0a242c64b8df,
	128'h6693dc911662ae473216ba22189a511a,
	128'h7606fa36d86473e6fb3a1bb0e2c0adf5,
	128'h112078e9e11fbb78e26ffb8899e96b9a,
	128'h40b264e921e9e4a82694589ef3798262,
	128'h8d4595cb4fa7026715f55bd68e2882f9,
	128'hb588a302bdbc09197df1edae68926ed9,
	128'h33f7502390b8a4a221cfecd0666624ba,
	128'h3d20253adbce3be2373767c4d822c566,
	128'ha42734a3929bf84cf0116c9856a3c18c,
	128'he3abc4939457422bb957da3c56938c6d,
	128'h972bdd2e7c525130fadc8f76fc6f4b3f,
	128'h84a83d7b94c699cbcb8a7d9b61f64093,
	128'hce61d63514aded03d43e6ebfc3a9001f,
	128'h6c839dd58eeae6b8a36af48ed63d2dc9,
	128'hcd5ece55b8da3bf622c4100df5de46f9,
	128'h3b6f46f40e0ac5fc0a9c1105f800f48d,
	128'hba26d47da3aeb028de4fb5b3a854a24b,
	128'h87f53bf620d3677268445212904389d5,
	128'h10617d28b5e0f4605492b182a5d7f9f6,
	128'h9aaec4fabbf6fae2a71feff02e372b39,
	128'h3a90c62d88b5c42809abf782488ed130,
	128'hf1f1c5a40899e15772857ccb65c7a09a,
	128'h190843d29b25a3897c692ce1dd81ee52,
	128'ha866bc65b6941d86e8420a7ffb0964db,
	128'h8193c6ff85225ced4255e92f6e078a14,
	128'h9661cb2424d7d4a380d547f9e7ec1cb9,
	128'h86f93d9ec08453a071e2e2877877a9c8,
	128'h27eefa80ce6a4a9d598e3fec365434d2,
	128'hd62068444578e3ab39ce7ec95dd045dc,
	128'hb5f71d4dd9a71fe5d8bc8ba7e6ea3048,
	128'h6825a347ac479d4f9d95c5cb8d3fd7e9,
	128'he3714e94a5778955cc0346358e94783a,
	128'hd836b44bb29e0c7d89fa4b2d4b677d2a,
	128'h5d454b75021d76d4b84f873a8f877b92,
	128'hc3498f7eced2095314fc28115885b33f,
	128'h6e668856539ad8e405bd123fe6c88530,
	128'h8680db7f3a87b8605543cfdbe6754076,
	128'h6c5d03b13069c3658b3179be91b0800c,
	128'hef1b384ac4d93eda00c92add0995ea5f,
	128'hbf8115805471741bd5ad20a03944790f,
	128'hc64c24b6894b038b3c0d09b1df068b0b,
	128'h3967a10cffe27d0178545fbf6a40544b,
	128'h7c85e9c95de1a9ec5a5363a8a053472d,
	128'ha9eec03c8abec7ba68315c2c8c2316e0,
	128'hcac8e414c2f388227ae14986fc983524,
	128'h5d942b7f4622ce056c3ce3ce5f1dd9d6,
	128'hd240d648ce21a3020282c3f1b528a0b6,
	128'h45d089c36d5c5a4efc689e3b0de10dd5,
	128'hb4da5df4becb5462e03a0ed00d295629,
	128'hdcf4e129136c1a4b7a0f38935cc34b2b,
	128'hd9a4c7618b0ce48a3d5aee1a1c0114c4,
	128'hca352df025c65c7b0bf306fbee0f36ba,
	128'h238aca23fd3409f38af63378ed2f5473,
	128'h59836a0e06a79691b36667d5380d8188,
	128'h33905080f7acf1cdae0a91fc3e85aee4,
	128'h72c9e4646dbc3d6320fc6689d93e8833,
	128'hba77413dea5925b7f5417ea47ff19f59,
	128'h6cae8129f843d86dc786a0fb1a184970,
	128'hfcfefb534100796eebbd990206754e19,
	128'h8c791d5fdddf470da04f3e6dc4a5b5b5,
	128'hc93bbdc07a4611ae4bb266ea5034a387,
	128'hc102e38e489aa74762f3efc5bb23205a,
	128'h93201481665cbafc1fcc220bc545fb3d,
	128'h4960757ec6ce68cf195e454cfd0f32ca,
	128'hfeec7ce6a6cbd07c043416737f1bbb33,
	128'h11c5413904487a805d70a8edd9c35527,
	128'h347846b2b2e36f1f0324c86f7f1b98e2,
	128'h332eee1a0cbd19ca2d69b426894044f0,
	128'h866b5b3977ba6efa5128efbda9ff03cd,
	128'hcc1445ee94c0f08cdee5c344ecd1e233,
	128'hbe288319029363c2622feba4b05dfdfe,
	128'hcfd1875523f3cd21c395651e6ee15e56,
	128'hcb5a408657837c53bf16f9d8465dce19,
	128'hca0bf42cb107f55ccff2fc09ee08ca15,
	128'hfdd9bbb4a7dc2e4a23536a5880a2db67,
	128'hede447b362c484993dec9442a3b46aef,
	128'h10dffb05904bff7c4781df780ad26837,
	128'hc33bc13e8de88ac25232aa7496398783,
	128'hca359c70803a3b2a3d542e8781dea975,
	128'hbcc65b526f88d05b89ce8a52021fdb06,
	128'hdb91a38855c8c4643851fbfb358b0109,
	128'hca6e8893a114ae8e27d5ab03a5499610,
	128'h6629d2b8df97da728cdd8b1e7f945077,
	128'h4570a5a18cfc0dd582f1d88d5c9a1720,
	128'h72bc65aa8e89562e3f274d45af1cd10b,
	128'h98551da1a6503276ae1c77625f9ea615,
	128'h0ddfe51ced7e3f4ae927daa3fe452cee,
	128'hdb826251e4ce384b80218b0e1da1dd4c,
	128'h2cacf728b88abbad7011ed0e64a1680c,
	128'h330d8ee7c5677e099ac74c9994ee4cfb,
	128'hedf61ae362e882ddc0167474a7a77f3a,
	128'h6168b00ba7859e0970ecfd757efecf7c,
	128'hd1415447866230d28bb1ea18a4cdfd02,
	128'h516183392f7a8763afec68a060264141,
	128'h77565c8d73cfd4130b4aa14d8911710f,
	128'h37232a4ed21ccc27c19c9610078cabac,
	128'h804f32ea71828c7d329077e712231666,
	128'hd64424f23cb97215e9c2c6f28d29eab7,
	128'h023e82b533f68c75c238cebdb2ee89a2,
	128'h193a3d24157a51f1ee0893f6777417e7,
	128'h84ecacfcd400084d078612b1945f2ef5,
	128'h1dcd8bb173259eb33a5242b0de31a455,
	128'h35e9eddbc375e792c19992c19165012b,
	128'h8a772231c01dfdd7c98e4cfddcc0807a,
	128'h6eda7ff6b8319180ff0d6e65629d01c3,
	128'hc267ef0e2d01a993944dd397101413cb,
	128'he9f80e9d845bcc0f62926af72eabca39,
	128'h6702990727aa0878637b45dcd3a3b074,
	128'h2e2e647d5360e09230a5d738ca33471e,
	128'h1f56413c7add6f43d1d56e4f02190330,
	128'h69cd0606e15af729d6bca143016d9842,
	128'ha085d7c1a500873a20099c4caa3c3f5b,
	128'h4fc0d230f8891415b87b83f95f2e09d1,
	128'h4327d08c523d8eba697a4336507d1f42,
	128'h7a15aab82701efa5ae36ab1d6b76290f,
	128'h5bf0051893a18bb30e139a58fed0fa54,
	128'h97e8adf65638fd9cdf3bc22c17fe4dbd,
	128'h1ee6ee326583a0586491c96418d1a35d,
	128'h26b549c2ec756f82ecc48008e529956b,
	128'h70377b6da669b072129e057cc28e9ca5,
	128'h9c94b8b0cb8bcc919072262b3fa05ad9,
	128'h2fbb83dfd0d7abcb05cd28cad2dfb523,
	128'h96877803de77744bb970d0a91f4debae,
	128'h7379f3370cf6e5ce12ae5969c8eea312,
	128'h02dc99fa3d4f98ce80985e7233889313,
	128'h1e38e759075ba5cab6457da51844295a,
	128'h70bed8dbf615868a1f9d9b05d3e7a267,
	128'h234b148b8cb1d8c32b287e896903d150,
	128'h294b033df4da853f4be3e243f7e513f4,
	128'h3f58c950f0367160adec45f2441e7411,
	128'h37f655536a704e5ace182d742a820cf4,
	128'hea7bd6bb63418731aeac790fe42d61e8,
	128'he74a4c999b4c064e48bb1e413f51e5ea,
	128'hba9ebefdb4ccf30f296cecb3bc1943e8,
	128'h3194367a4898c502c13bb7478640a72d,
	128'hda797713263d6f33a5478a65ef60d412,
	128'hd1ac39bb1ef86b9c1344f214679aa376,
	128'h2fdea9e650532be5bc0e7325337fd363,
	128'hd3a204dbd9c2af158b6ca67a5156ce4a,
	128'h3a0a0e75a8da36735aee6684d965a778,
	128'h52fc3e620492ea99641ea168da5b6d52,
	128'hd2e0c7f15b4772467d2cfc873000b2ca,
	128'h563531135e0c4d70a38f8bdb190ba04e,
	128'ha8a39a0f5663f4c0fe5f2d3cafff421a,
	128'hd94b5e90db354c1e42f61fabe167b2c0,
	128'h50e6d3c9b6698a7cd276f96b1473f35a,
	128'h9338f08e0ebee96905d8f2e825208f43,
	128'h8b378c86672aa54a3a266ba19d2580ca,
	128'hcca7c3086f5f9511b31233da7cab9160,
	128'h5b40ff4ec9be536ba23035fa4f06064c,
	128'h60eb5af8416b257149372194e8b88749,
	128'h2f005a8aed8a361c92e440c15520cbd1,
	128'h7b03627611678a997717578807a800e2,
	128'hcf78618f74f6f3696e0a4779b90b5a77,
	128'h03720371a04962eaea0a852e69972858,
	128'h1f8a8133aa8ccf70e2bd3285831ca6b7,
	128'h27936bd27fb1468fc8b48bc483321725,
	128'hb07d4f3e2cd2ef2eb545980754dfea0f,
	128'h4bf85f1b5d54adbc307b0a048389adcb
	};