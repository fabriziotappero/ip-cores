-------------------------------------------------------------------------------
--
-- The Timer/Counter unit.
--
-- $Id: timer-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_timer_rtl_c0 of t48_timer is

  for rtl
  end for;

end t48_timer_rtl_c0;
