-------------------------------------------------------------------------------
--
-- The reset generation unit.
--
-- $Id: t400_reset-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_reset_rtl_c0 of t400_reset is

  for rtl
  end for;

end t400_reset_rtl_c0;
