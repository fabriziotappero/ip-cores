----------------------------------------------------------------------------
--  This file is a part of the LM VHDL IP LIBRARY
--  Copyright (C) 2009 Jose Nunez-Yanez
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  See the file COPYING for the full details of the license.
--
--  The license allows free and unlimited use of the library and tools for research and education purposes. 
--  The full LM core supports many more advanced motion estimation features and it is available under a 
--  low-cost commercial license. See the readme file to learn more or contact us at 
--  eejlny@byacom.co.uk or www.byacom.co.uk
-----------------------------------------------------------------------------
-- Entity: 	
-- File:	reference_data.vhd
-- Author:	Jose Luis Nunez 
-- Description:	reference data 5x5 macroblocks 
------------------------------------------------------------------------------



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.Numeric_STD.all;
use IEEE.std_logic_unsigned."<";

entity reference_data1 is
    port(
      clk : in std_logic;
      reset : in std_logic;
      clear : in std_logic;
      addr : in std_logic_vector (9 downto 0);
      data : out std_logic_vector (63 downto 0)
      );
end;


architecture rtl of reference_data1 is

signal data_int: std_logic_vector(63 downto 0);

subtype word is integer range 0 to 255;
type mem is array (0 to 6399) of word;

signal memory : mem := ( 
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#53#,16#4C#,16#49#,16#4C#,16#50#,16#53#,16#4E#,16#50#,16#56#,16#46#,16#A2#,16#DF#,16#CA#,16#DC#,16#F5#,16#FD#,16#87#,16#1D#,16#47#,16#C3#,16#D5#,16#C8#,16#DB#,16#EC#,16#E5#,16#82#,16#35#,16#43#,16#47#,16#5C#,16#C9#,16#D7#,16#C6#,16#CF#,16#D7#,16#D7#,16#E6#,16#E2#,16#DF#,16#F3#,16#D2#,16#43#,16#39#,16#BC#,16#EE#,16#EB#,16#DD#,16#91#,16#32#,16#03#,16#57#,16#E9#,16#E9#,16#AE#,16#A8#,16#B3#,16#B2#,16#A5#,16#B0#,16#BD#,16#54#,16#3D#,16#CE#,16#D8#,16#A7#,16#6F#,16#22#,16#1F#,
16#49#,16#47#,16#48#,16#4B#,16#4B#,16#4B#,16#49#,16#49#,16#4A#,16#4B#,16#4C#,16#4C#,16#4F#,16#4A#,16#48#,16#4C#,16#4B#,16#51#,16#42#,16#40#,16#4B#,16#3C#,16#4B#,16#59#,16#5A#,16#95#,16#B6#,16#D6#,16#E3#,16#56#,16#33#,16#C8#,16#DD#,16#C3#,16#D2#,16#D0#,16#D0#,16#E2#,16#C9#,16#6D#,16#28#,16#4A#,16#C7#,16#D9#,16#C3#,16#C9#,16#CB#,16#C8#,16#CA#,16#D1#,16#E2#,16#BD#,16#45#,16#66#,16#CE#,16#D9#,16#D1#,16#D1#,16#D0#,16#DA#,16#BD#,16#4A#,16#15#,16#74#,16#DE#,16#C0#,16#9F#,16#B2#,16#AF#,16#A6#,16#B0#,16#8C#,16#1C#,16#4A#,16#C6#,16#B7#,16#A6#,16#BB#,16#A1#,16#69#,
16#4A#,16#43#,16#43#,16#4A#,16#4C#,16#4A#,16#49#,16#49#,16#4A#,16#4B#,16#4B#,16#4B#,16#49#,16#45#,16#47#,16#4C#,16#4E#,16#4A#,16#37#,16#4E#,16#48#,16#34#,16#58#,16#4B#,16#38#,16#5E#,16#53#,16#5D#,16#ED#,16#AF#,16#3C#,16#C3#,16#D8#,16#C1#,16#C9#,16#BD#,16#C6#,16#E9#,16#FC#,16#CB#,16#43#,16#2F#,16#BA#,16#DA#,16#C3#,16#C9#,16#CB#,16#C8#,16#C6#,16#DA#,16#BC#,16#48#,16#3B#,16#C8#,16#FF#,16#CC#,16#BD#,16#CD#,16#C9#,16#E2#,16#FE#,16#C1#,16#2E#,16#0A#,16#92#,16#D0#,16#AC#,16#A7#,16#A9#,16#A8#,16#B6#,16#69#,16#10#,16#5C#,16#B4#,16#AC#,16#A8#,16#C7#,16#DE#,16#C9#,
16#4B#,16#44#,16#44#,16#4A#,16#4C#,16#4A#,16#49#,16#49#,16#4A#,16#4B#,16#4B#,16#4A#,16#48#,16#44#,16#46#,16#4D#,16#53#,16#2E#,16#34#,16#8D#,16#58#,16#2C#,16#8E#,16#82#,16#6A#,16#61#,16#48#,16#37#,16#7B#,16#C3#,16#BB#,16#BE#,16#CC#,16#C4#,16#C8#,16#C7#,16#C2#,16#BC#,16#CA#,16#FE#,16#AC#,16#2E#,16#A7#,16#E5#,16#C6#,16#CF#,16#D7#,16#D7#,16#D9#,16#A3#,16#55#,16#2B#,16#74#,16#DA#,16#CD#,16#B2#,16#C1#,16#CC#,16#C8#,16#C3#,16#CC#,16#ED#,16#A9#,16#1B#,16#31#,16#B6#,16#BC#,16#A1#,16#A7#,16#A9#,16#B5#,16#75#,16#1D#,16#66#,16#C1#,16#C4#,16#B5#,16#95#,16#7B#,16#8F#,
16#4B#,16#49#,16#45#,16#4A#,16#4A#,16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4A#,16#4A#,16#48#,16#48#,16#49#,16#58#,16#3E#,16#2F#,16#6B#,16#93#,16#67#,16#54#,16#79#,16#6F#,16#6B#,16#6E#,16#75#,16#78#,16#4A#,16#6C#,16#CF#,16#EB#,16#CC#,16#C0#,16#CC#,16#CB#,16#CC#,16#C7#,16#C6#,16#D9#,16#E6#,16#7E#,16#92#,16#E0#,16#C7#,16#CB#,16#BE#,16#A9#,16#82#,16#36#,16#30#,16#49#,16#48#,16#B1#,16#D9#,16#BB#,16#C7#,16#C7#,16#CF#,16#D8#,16#D9#,16#EE#,16#FA#,16#9E#,16#19#,16#6E#,16#CE#,16#AE#,16#A1#,16#AB#,16#B4#,16#6C#,16#28#,16#82#,16#AC#,16#7D#,16#72#,16#5A#,16#3A#,16#3C#,
16#48#,16#48#,16#48#,16#49#,16#4A#,16#4A#,16#4A#,16#4A#,16#4B#,16#4B#,16#4B#,16#4B#,16#4A#,16#4C#,16#4F#,16#44#,16#2D#,16#5F#,16#8E#,16#75#,16#6C#,16#6C#,16#74#,16#6A#,16#6D#,16#6D#,16#6C#,16#6B#,16#70#,16#58#,16#69#,16#C2#,16#E3#,16#C6#,16#BF#,16#C8#,16#C8#,16#C6#,16#C1#,16#C0#,16#DC#,16#B8#,16#A2#,16#C7#,16#D2#,16#A2#,16#5A#,16#46#,16#2E#,16#1F#,16#3A#,16#33#,16#5B#,16#BF#,16#D0#,16#B9#,16#C0#,16#EA#,16#E6#,16#D3#,16#C7#,16#C0#,16#D7#,16#DA#,16#52#,16#24#,16#B1#,16#DF#,16#AC#,16#B0#,16#C1#,16#5B#,16#19#,16#71#,16#6E#,16#30#,16#31#,16#3E#,16#4C#,16#53#,
16#46#,16#47#,16#49#,16#4A#,16#4A#,16#4A#,16#4A#,16#4A#,16#4B#,16#4C#,16#4B#,16#4B#,16#47#,16#54#,16#51#,16#32#,16#4C#,16#8B#,16#83#,16#58#,16#6F#,16#76#,16#69#,16#68#,16#6B#,16#6B#,16#67#,16#64#,16#6F#,16#6E#,16#47#,16#53#,16#BE#,16#DC#,16#C3#,16#BD#,16#C2#,16#C5#,16#C3#,16#BE#,16#C8#,16#DB#,16#C6#,16#C4#,16#CD#,16#85#,16#1B#,16#11#,16#1A#,16#30#,16#37#,16#28#,16#76#,16#D7#,16#C4#,16#C3#,16#C2#,16#C0#,16#AF#,16#80#,16#62#,16#4B#,16#50#,16#88#,16#6F#,16#07#,16#51#,16#C7#,16#BF#,16#B1#,16#97#,16#3F#,16#17#,16#41#,16#49#,16#44#,16#4A#,16#52#,16#5A#,16#59#,
16#45#,16#47#,16#49#,16#4A#,16#4A#,16#4A#,16#4A#,16#4A#,16#4B#,16#4C#,16#4B#,16#4C#,16#4C#,16#4C#,16#3F#,16#41#,16#7D#,16#83#,16#66#,16#62#,16#6D#,16#6A#,16#63#,16#68#,16#6A#,16#6A#,16#69#,16#69#,16#69#,16#74#,16#69#,16#41#,16#68#,16#C4#,16#D8#,16#BA#,16#BE#,16#C5#,16#C8#,16#C6#,16#C2#,16#C7#,16#CF#,16#C8#,16#CC#,16#95#,16#35#,16#2B#,16#32#,16#3A#,16#3D#,16#24#,16#7D#,16#E0#,16#C0#,16#CB#,16#A7#,16#49#,16#31#,16#2F#,16#28#,16#24#,16#1E#,16#34#,16#51#,16#3A#,16#19#,16#3B#,16#A5#,16#A4#,16#40#,16#30#,16#49#,16#48#,16#52#,16#5C#,16#5C#,16#5C#,16#5A#,16#59#,
16#45#,16#47#,16#48#,16#4A#,16#4A#,16#4A#,16#4A#,16#4A#,16#4C#,16#4D#,16#4A#,16#48#,16#4E#,16#40#,16#2E#,16#73#,16#87#,16#67#,16#6A#,16#69#,16#6B#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#68#,16#69#,16#6B#,16#6D#,16#46#,16#5E#,16#B9#,16#EA#,16#D4#,16#CA#,16#CA#,16#CA#,16#CA#,16#CC#,16#C6#,16#C3#,16#CF#,16#A2#,16#3D#,16#3F#,16#48#,16#36#,16#36#,16#12#,16#79#,16#EB#,16#C5#,16#AF#,16#70#,16#24#,16#20#,16#33#,16#39#,16#3E#,16#43#,16#43#,16#42#,16#50#,16#32#,16#0A#,16#44#,16#4C#,16#27#,16#45#,16#69#,16#60#,16#55#,16#5B#,16#57#,16#57#,16#59#,16#57#,
16#44#,16#47#,16#49#,16#4A#,16#49#,16#4A#,16#4A#,16#4A#,16#47#,16#4C#,16#47#,16#53#,16#44#,16#2B#,16#59#,16#8E#,16#73#,16#62#,16#6F#,16#69#,16#69#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#68#,16#69#,16#6B#,16#6D#,16#6A#,16#48#,16#59#,16#90#,16#C0#,16#D0#,16#D8#,16#D3#,16#CB#,16#CB#,16#CA#,16#C5#,16#CF#,16#C5#,16#50#,16#01#,16#21#,16#11#,16#11#,16#56#,16#D0#,16#CA#,16#87#,16#59#,16#3E#,16#49#,16#53#,16#4A#,16#4C#,16#4C#,16#4C#,16#4C#,16#49#,16#42#,16#44#,16#39#,16#18#,16#20#,16#37#,16#63#,16#71#,16#52#,16#55#,16#55#,16#56#,16#56#,16#58#,16#57#,
16#43#,16#47#,16#48#,16#4A#,16#49#,16#4A#,16#4A#,16#4A#,16#46#,16#4C#,16#4E#,16#4F#,16#2F#,16#4A#,16#80#,16#73#,16#62#,16#69#,16#6C#,16#65#,16#68#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#68#,16#6A#,16#6C#,16#6C#,16#6B#,16#6B#,16#4A#,16#3E#,16#7F#,16#95#,16#AC#,16#C5#,16#E0#,16#D7#,16#CC#,16#C5#,16#C0#,16#E0#,16#B2#,16#5B#,16#48#,16#43#,16#76#,16#D1#,16#D1#,16#79#,16#3B#,16#34#,16#3E#,16#48#,16#47#,16#48#,16#47#,16#46#,16#46#,16#46#,16#47#,16#43#,16#3C#,16#3E#,16#41#,16#3F#,16#2E#,16#3C#,16#5E#,16#6A#,16#5D#,16#53#,16#57#,16#57#,16#58#,16#57#,
16#43#,16#47#,16#48#,16#4A#,16#49#,16#49#,16#4A#,16#4A#,16#4A#,16#4E#,16#58#,16#3C#,16#36#,16#78#,16#7A#,16#5E#,16#63#,16#68#,16#67#,16#66#,16#67#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6B#,16#6B#,16#6B#,16#6B#,16#6A#,16#65#,16#5E#,16#59#,16#5B#,16#7D#,16#AD#,16#BF#,16#D7#,16#E0#,16#C9#,16#BD#,16#D2#,16#E7#,16#D4#,16#D0#,16#EC#,16#B3#,16#6D#,16#41#,16#3D#,16#43#,16#43#,16#41#,16#4A#,16#48#,16#47#,16#46#,16#46#,16#46#,16#45#,16#44#,16#3E#,16#3D#,16#3E#,16#3D#,16#3A#,16#2A#,16#3B#,16#5D#,16#64#,16#61#,16#57#,16#57#,16#59#,16#57#,
16#43#,16#47#,16#48#,16#49#,16#49#,16#4A#,16#4A#,16#49#,16#49#,16#4E#,16#44#,16#2D#,16#64#,16#83#,16#6B#,16#66#,16#65#,16#68#,16#67#,16#67#,16#67#,16#67#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#69#,16#68#,16#63#,16#5E#,16#58#,16#54#,16#45#,16#70#,16#AD#,16#C8#,16#DA#,16#D6#,16#D4#,16#FE#,16#FF#,16#DA#,16#9F#,16#58#,16#2D#,16#3A#,16#47#,16#49#,16#44#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#44#,16#3E#,16#3D#,16#3E#,16#3D#,16#3D#,16#37#,16#32#,16#2D#,16#46#,16#5D#,16#56#,16#5D#,16#5B#,16#59#,
16#41#,16#45#,16#47#,16#49#,16#4B#,16#4A#,16#48#,16#44#,16#4C#,16#47#,16#32#,16#55#,16#86#,16#6C#,16#64#,16#6A#,16#66#,16#68#,16#67#,16#67#,16#67#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#69#,16#68#,16#67#,16#64#,16#4F#,16#56#,16#50#,16#5A#,16#B5#,16#DD#,16#C4#,16#BE#,16#96#,16#4B#,16#2F#,16#33#,16#3C#,16#47#,16#4B#,16#46#,16#44#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3E#,16#3D#,16#3D#,16#3B#,16#39#,16#2B#,16#2E#,16#36#,16#41#,16#58#,16#5B#,16#5A#,
16#47#,16#4B#,16#4C#,16#4B#,16#4B#,16#4A#,16#49#,16#48#,16#52#,16#37#,16#3F#,16#84#,16#7A#,16#62#,16#68#,16#68#,16#67#,16#68#,16#68#,16#68#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6B#,16#6B#,16#6B#,16#6B#,16#6A#,16#73#,16#65#,16#4E#,16#49#,16#4E#,16#8C#,16#AD#,16#58#,16#29#,16#1C#,16#2B#,16#43#,16#4A#,16#4C#,16#4A#,16#45#,16#44#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3E#,16#3E#,16#3D#,16#3D#,16#3D#,16#3C#,16#44#,16#36#,16#27#,16#2E#,16#3B#,16#3A#,16#3A#,
16#22#,16#26#,16#28#,16#27#,16#26#,16#2A#,16#30#,16#33#,16#35#,16#28#,16#6E#,16#7F#,16#5E#,16#67#,16#68#,16#63#,16#67#,16#68#,16#68#,16#68#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6B#,16#6B#,16#6B#,16#6B#,16#6A#,16#6A#,16#6B#,16#72#,16#71#,16#46#,16#50#,16#46#,16#0A#,16#26#,16#4C#,16#4C#,16#48#,16#49#,16#45#,16#45#,16#45#,16#44#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3E#,16#3E#,16#3D#,16#3D#,16#3D#,16#3C#,16#45#,16#3F#,16#40#,16#37#,16#2C#,16#31#,16#2D#,
16#3C#,16#3D#,16#34#,16#37#,16#38#,16#37#,16#36#,16#34#,16#2E#,16#57#,16#7C#,16#72#,16#63#,16#69#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6F#,16#62#,16#3A#,16#1D#,16#39#,16#50#,16#44#,16#48#,16#48#,16#48#,16#47#,16#46#,16#45#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3D#,16#3C#,16#3C#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#80#,16#83#,16#6C#,16#6F#,16#76#,16#6F#,16#6F#,16#5A#,16#4D#,16#7F#,16#77#,16#65#,16#66#,16#67#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#63#,16#70#,16#77#,16#51#,16#29#,16#41#,16#4B#,16#48#,16#48#,16#48#,16#47#,16#46#,16#45#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3D#,16#3C#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#94#,16#89#,16#76#,16#73#,16#75#,16#6D#,16#79#,16#6E#,16#5B#,16#69#,16#6F#,16#70#,16#6A#,16#68#,16#67#,16#67#,16#68#,16#68#,16#68#,16#69#,16#68#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6C#,16#77#,16#7F#,16#45#,16#35#,16#4A#,16#4A#,16#48#,16#48#,16#47#,16#47#,16#45#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#46#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3A#,
16#83#,16#69#,16#6A#,16#65#,16#6D#,16#64#,16#66#,16#71#,16#64#,16#4D#,16#5E#,16#70#,16#68#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#69#,16#68#,16#68#,16#68#,16#6A#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6F#,16#67#,16#7C#,16#70#,16#37#,16#40#,16#4E#,16#48#,16#49#,16#48#,16#47#,16#45#,16#41#,16#4A#,16#48#,16#47#,16#47#,16#47#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#41#,16#2F#,16#5D#,16#73#,16#73#,16#68#,16#66#,16#70#,16#73#,16#62#,16#42#,16#3F#,16#66#,16#6E#,16#6C#,16#6F#,16#6F#,16#67#,16#65#,16#6B#,16#70#,16#73#,16#70#,16#69#,16#69#,16#73#,16#72#,16#72#,16#72#,16#73#,16#69#,16#60#,16#5A#,16#5B#,16#5E#,16#60#,16#5F#,16#5E#,16#67#,16#6B#,16#77#,16#76#,16#74#,16#74#,16#73#,16#71#,16#6C#,16#75#,16#67#,16#46#,16#47#,16#4B#,16#49#,16#48#,16#48#,16#48#,16#46#,16#42#,16#49#,16#47#,16#47#,16#47#,16#47#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3A#,
16#60#,16#53#,16#41#,16#37#,16#35#,16#45#,16#4A#,16#3F#,16#40#,16#4D#,16#51#,16#59#,16#4D#,16#3C#,16#48#,16#44#,16#4A#,16#57#,16#69#,16#6D#,16#63#,16#57#,16#5A#,16#69#,16#66#,16#66#,16#50#,16#3D#,16#3C#,16#38#,16#49#,16#5F#,16#61#,16#60#,16#5D#,16#5C#,16#5B#,16#54#,16#4D#,16#51#,16#68#,16#60#,16#64#,16#6B#,16#6F#,16#70#,16#75#,16#6C#,16#58#,16#48#,16#49#,16#4A#,16#49#,16#49#,16#48#,16#48#,16#46#,16#42#,16#49#,16#47#,16#47#,16#47#,16#47#,16#46#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#DE#,16#CD#,16#94#,16#72#,16#57#,16#54#,16#55#,16#59#,16#55#,16#6C#,16#9D#,16#BF#,16#8B#,16#5F#,16#5B#,16#5E#,16#77#,16#78#,16#62#,16#53#,16#5D#,16#51#,16#54#,16#63#,16#5A#,16#4A#,16#72#,16#88#,16#68#,16#69#,16#85#,16#A1#,16#A9#,16#A8#,16#A5#,16#A3#,16#A4#,16#94#,16#8A#,16#6F#,16#3A#,16#3C#,16#4F#,16#4E#,16#4D#,16#4D#,16#53#,16#4A#,16#45#,16#4A#,16#49#,16#4A#,16#49#,16#49#,16#48#,16#48#,16#46#,16#43#,16#49#,16#47#,16#47#,16#47#,16#47#,16#47#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#DB#,16#E4#,16#F3#,16#F0#,16#ED#,16#CF#,16#B4#,16#B7#,16#BC#,16#CD#,16#D0#,16#D5#,16#D5#,16#CA#,16#CC#,16#C8#,16#AE#,16#94#,16#62#,16#4D#,16#65#,16#68#,16#65#,16#5F#,16#5E#,16#51#,16#84#,16#DC#,16#FF#,16#F8#,16#DF#,16#CE#,16#D3#,16#D5#,16#D7#,16#D9#,16#D9#,16#D0#,16#E4#,16#B1#,16#1C#,16#2E#,16#48#,16#3B#,16#3B#,16#3B#,16#35#,16#3E#,16#47#,16#49#,16#49#,16#4A#,16#4A#,16#48#,16#48#,16#48#,16#46#,16#44#,16#49#,16#47#,16#47#,16#47#,16#47#,16#47#,16#45#,16#43#,16#3D#,16#3D#,16#3D#,16#3C#,16#3B#,16#3B#,16#3B#,16#3B#,16#3A#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#8D#,16#A1#,16#B6#,16#B6#,16#DD#,16#F5#,16#FB#,16#EF#,16#DF#,16#DD#,16#CC#,16#CB#,16#D6#,16#E8#,16#F4#,16#CF#,16#86#,16#71#,16#6E#,16#66#,16#6C#,16#6B#,16#6A#,16#6A#,16#6A#,16#6E#,16#52#,16#82#,16#D3#,16#E9#,16#ED#,16#DD#,16#CE#,16#CD#,16#CD#,16#D3#,16#D8#,16#CF#,16#E5#,16#CD#,16#37#,16#15#,16#45#,16#46#,16#45#,16#42#,16#3F#,16#4A#,16#47#,16#48#,16#49#,16#49#,16#4A#,16#49#,16#48#,16#47#,16#46#,16#46#,16#4F#,16#54#,16#42#,16#3C#,16#39#,16#3B#,16#46#,16#46#,16#47#,16#44#,16#41#,16#3C#,16#3D#,16#43#,16#39#,16#39#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,16#3B#,
16#47#,16#4B#,16#46#,16#3B#,16#51#,16#94#,16#C8#,16#D0#,16#CA#,16#C2#,16#C1#,16#C5#,16#C8#,16#CE#,16#9D#,16#64#,16#65#,16#65#,16#6B#,16#6D#,16#6C#,16#69#,16#67#,16#68#,16#68#,16#70#,16#59#,16#49#,16#3A#,16#4C#,16#B3#,16#D2#,16#BC#,16#C0#,16#C2#,16#C7#,16#CA#,16#C5#,16#BC#,16#DD#,16#A4#,16#2B#,16#29#,16#4B#,16#53#,16#4C#,16#48#,16#4E#,16#4D#,16#4C#,16#4A#,16#49#,16#48#,16#4A#,16#4A#,16#48#,16#46#,16#45#,16#43#,16#44#,16#3C#,16#33#,16#30#,16#35#,16#39#,16#40#,16#42#,16#3E#,16#3C#,16#40#,16#3F#,16#3A#,16#40#,16#3F#,16#3C#,16#3B#,16#3B#,16#3B#,16#3C#,16#3C#,
16#52#,16#51#,16#4B#,16#47#,16#3E#,16#3E#,16#48#,16#75#,16#BC#,16#E3#,16#D5#,16#C6#,16#C7#,16#84#,16#4B#,16#54#,16#68#,16#6E#,16#66#,16#65#,16#65#,16#68#,16#68#,16#68#,16#68#,16#67#,16#6E#,16#68#,16#3B#,16#3A#,16#50#,16#A3#,16#DE#,16#C6#,16#C5#,16#CA#,16#C3#,16#C4#,16#C2#,16#D3#,16#E3#,16#B0#,16#3F#,16#18#,16#22#,16#3F#,16#4B#,16#4D#,16#4E#,16#4F#,16#50#,16#51#,16#50#,16#4E#,16#4C#,16#4B#,16#45#,16#2A#,16#16#,16#1F#,16#44#,16#5B#,16#6A#,16#62#,16#4F#,16#31#,16#19#,16#24#,16#29#,16#35#,16#3D#,16#39#,16#3E#,16#3F#,16#3E#,16#3D#,16#3C#,16#3C#,16#3B#,16#3B#,
16#6E#,16#6E#,16#70#,16#73#,16#71#,16#53#,16#38#,16#44#,16#67#,16#81#,16#B4#,16#E1#,16#99#,16#54#,16#51#,16#75#,16#6E#,16#69#,16#69#,16#68#,16#68#,16#68#,16#69#,16#69#,16#63#,16#67#,16#6A#,16#71#,16#81#,16#75#,16#3D#,16#47#,16#AD#,16#E4#,16#C8#,16#BB#,16#C0#,16#C1#,16#C1#,16#C0#,16#DC#,16#FB#,16#B9#,16#79#,16#54#,16#27#,16#1C#,16#1E#,16#1F#,16#24#,16#2D#,16#32#,16#3B#,16#36#,16#2D#,16#28#,16#18#,16#4B#,16#80#,16#80#,16#AF#,16#C4#,16#D2#,16#CD#,16#B9#,16#8A#,16#5F#,16#5A#,16#3D#,16#2A#,16#14#,16#19#,16#29#,16#32#,16#3E#,16#42#,16#3B#,16#3B#,16#3B#,16#3C#,
16#67#,16#67#,16#67#,16#67#,16#6A#,16#6E#,16#6E#,16#6A#,16#45#,16#39#,16#76#,16#91#,16#56#,16#72#,16#79#,16#64#,16#6F#,16#6B#,16#69#,16#69#,16#68#,16#69#,16#69#,16#69#,16#69#,16#68#,16#68#,16#6A#,16#6C#,16#70#,16#73#,16#56#,16#49#,16#B1#,16#F3#,16#CC#,16#BB#,16#C5#,16#C0#,16#C8#,16#C2#,16#CA#,16#E5#,16#EE#,16#C6#,16#83#,16#61#,16#57#,16#4C#,16#42#,16#40#,16#36#,16#36#,16#33#,16#39#,16#42#,16#4D#,16#B0#,16#FB#,16#EE#,16#E6#,16#E6#,16#E6#,16#E6#,16#E7#,16#DB#,16#C2#,16#B4#,16#95#,16#6D#,16#56#,16#4C#,16#3C#,16#1F#,16#14#,16#1B#,16#1E#,16#2E#,16#3A#,16#36#,
16#67#,16#67#,16#67#,16#67#,16#6D#,16#69#,16#69#,16#6D#,16#65#,16#68#,16#5F#,16#40#,16#43#,16#65#,16#6D#,16#65#,16#72#,16#6F#,16#69#,16#68#,16#68#,16#69#,16#69#,16#69#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6B#,16#66#,16#73#,16#55#,16#45#,16#AD#,16#EF#,16#CD#,16#BC#,16#BD#,16#C1#,16#C6#,16#C7#,16#C3#,16#C8#,16#E0#,16#E9#,16#E9#,16#D4#,16#C1#,16#B4#,16#A3#,16#96#,16#8D#,16#90#,16#9C#,16#A5#,16#C9#,16#D6#,16#D5#,16#C3#,16#C2#,16#C2#,16#C2#,16#C2#,16#C4#,16#B5#,16#AF#,16#B6#,16#BD#,16#BF#,16#BF#,16#AE#,16#89#,16#5A#,16#34#,16#2A#,16#26#,16#22#,16#1C#,16#1B#,
16#67#,16#67#,16#67#,16#67#,16#6A#,16#68#,16#68#,16#6A#,16#6D#,16#74#,16#67#,16#5A#,16#56#,16#48#,16#4E#,16#63#,16#67#,16#69#,16#69#,16#68#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#69#,16#69#,16#69#,16#69#,16#69#,16#65#,16#71#,16#71#,16#41#,16#48#,16#B6#,16#E0#,16#D1#,16#BF#,16#C4#,16#C8#,16#C7#,16#C3#,16#BF#,16#D1#,16#E1#,16#E6#,16#E3#,16#ED#,16#EF#,16#E9#,16#EB#,16#EC#,16#ED#,16#E7#,16#E1#,16#DC#,16#D3#,16#C4#,16#BC#,16#C1#,16#C1#,16#C1#,16#C1#,16#C3#,16#AE#,16#A3#,16#AE#,16#B5#,16#BB#,16#C1#,16#BA#,16#BA#,16#BD#,16#B9#,16#97#,16#74#,16#61#,16#4A#,16#45#,
16#67#,16#67#,16#67#,16#67#,16#64#,16#67#,16#67#,16#64#,16#68#,16#66#,16#68#,16#74#,16#6A#,16#5C#,16#61#,16#61#,16#50#,16#5D#,16#6B#,16#6B#,16#6B#,16#6A#,16#6A#,16#6A#,16#6A#,16#69#,16#69#,16#69#,16#69#,16#69#,16#6B#,16#61#,16#6F#,16#76#,16#3F#,16#46#,16#AC#,16#D9#,16#C3#,16#C6#,16#C7#,16#C7#,16#C6#,16#C6#,16#C4#,16#C1#,16#CB#,16#C5#,16#CC#,16#D6#,16#D8#,16#E2#,16#E8#,16#E8#,16#DC#,16#D0#,16#C7#,16#C9#,16#C8#,16#C8#,16#C8#,16#C9#,16#CA#,16#CA#,16#C9#,16#B7#,16#A8#,16#AD#,16#AE#,16#A2#,16#A5#,16#A6#,16#B5#,16#C2#,16#CB#,16#BE#,16#BA#,16#B5#,16#AF#,16#AD#,
16#67#,16#67#,16#67#,16#67#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#69#,16#6B#,16#6F#,16#71#,16#6B#,16#63#,16#5F#,16#56#,16#52#,16#6D#,16#6F#,16#6D#,16#6A#,16#6A#,16#6A#,16#69#,16#69#,16#6A#,16#69#,16#69#,16#69#,16#68#,16#6B#,16#76#,16#6B#,16#49#,16#48#,16#B4#,16#E6#,16#C3#,16#C5#,16#C8#,16#C7#,16#CB#,16#C8#,16#C8#,16#C7#,16#C7#,16#C6#,16#C6#,16#C5#,16#C4#,16#C4#,16#C3#,16#C3#,16#C3#,16#C4#,16#CA#,16#CC#,16#C8#,16#CE#,16#CC#,16#C9#,16#C8#,16#CA#,16#BD#,16#A8#,16#AE#,16#B0#,16#AB#,16#A8#,16#A8#,16#A6#,16#A4#,16#A2#,16#A1#,16#B3#,16#BB#,16#C4#,16#C1#,
16#67#,16#67#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#68#,16#68#,16#69#,16#68#,16#68#,16#6A#,16#6D#,16#6D#,16#74#,16#68#,16#58#,16#58#,16#69#,16#69#,16#6A#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#69#,16#69#,16#69#,16#69#,16#68#,16#61#,16#6E#,16#75#,16#40#,16#4B#,16#BD#,16#DB#,16#BD#,16#C8#,16#CC#,16#CB#,16#C9#,16#C9#,16#C8#,16#C8#,16#C7#,16#C7#,16#C7#,16#C8#,16#C8#,16#C8#,16#C9#,16#C9#,16#C8#,16#CC#,16#CC#,16#C8#,16#CC#,16#CB#,16#C8#,16#C7#,16#C9#,16#BB#,16#A7#,16#AE#,16#AE#,16#AB#,16#A7#,16#A6#,16#A4#,16#A3#,16#A3#,16#A3#,16#A3#,16#A5#,16#A0#,16#A0#,
16#67#,16#67#,16#67#,16#67#,16#67#,16#68#,16#68#,16#69#,16#68#,16#69#,16#69#,16#68#,16#69#,16#68#,16#67#,16#6A#,16#67#,16#71#,16#71#,16#5A#,16#58#,16#65#,16#6D#,16#63#,16#65#,16#65#,16#66#,16#66#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#6A#,16#6B#,16#6F#,16#6E#,16#3E#,16#62#,16#D8#,16#D8#,16#BD#,16#C6#,16#C7#,16#C8#,16#C8#,16#C8#,16#C8#,16#C8#,16#C9#,16#C9#,16#C9#,16#C9#,16#C9#,16#CA#,16#CA#,16#C7#,16#CB#,16#CC#,16#C8#,16#C8#,16#C7#,16#C4#,16#C3#,16#C6#,16#B8#,16#A4#,16#AB#,16#AD#,16#AB#,16#A7#,16#A4#,16#A5#,16#A5#,16#A5#,16#A5#,16#A6#,16#A6#,16#A1#,16#A5#,
16#67#,16#67#,16#67#,16#67#,16#68#,16#68#,16#68#,16#69#,16#69#,16#6A#,16#6A#,16#6A#,16#6A#,16#68#,16#6B#,16#6A#,16#68#,16#67#,16#74#,16#6A#,16#58#,16#74#,16#78#,16#70#,16#6E#,16#6E#,16#6D#,16#6C#,16#6A#,16#6B#,16#6B#,16#6C#,16#6C#,16#6C#,16#6B#,16#67#,16#74#,16#6D#,16#49#,16#82#,16#D7#,16#C7#,16#BF#,16#CC#,16#C8#,16#C9#,16#C9#,16#CA#,16#CA#,16#CB#,16#CA#,16#CA#,16#CA#,16#C9#,16#CA#,16#C9#,16#C6#,16#CB#,16#CB#,16#C9#,16#C7#,16#C7#,16#C4#,16#C1#,16#C5#,16#B8#,16#A2#,16#AB#,16#AC#,16#A9#,16#A7#,16#A5#,16#A7#,16#A7#,16#A7#,16#A7#,16#A7#,16#A7#,16#A5#,16#A5#,
16#67#,16#67#,16#68#,16#68#,16#68#,16#68#,16#69#,16#6A#,16#69#,16#69#,16#69#,16#6B#,16#69#,16#69#,16#6A#,16#70#,16#69#,16#6D#,16#67#,16#48#,16#49#,16#5D#,16#56#,16#5C#,16#58#,16#5A#,16#5F#,16#63#,16#6A#,16#6F#,16#71#,16#6F#,16#69#,16#6D#,16#6C#,16#67#,16#67#,16#78#,16#63#,16#4C#,16#A0#,16#DF#,16#C4#,16#C3#,16#C8#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CA#,16#C9#,16#C9#,16#C5#,16#CA#,16#CC#,16#C9#,16#CB#,16#CA#,16#C8#,16#C4#,16#CE#,16#BB#,16#A2#,16#AB#,16#AC#,16#A9#,16#A8#,16#A6#,16#A7#,16#A7#,16#A7#,16#A8#,16#A8#,16#A7#,16#AA#,16#A8#,
16#69#,16#69#,16#69#,16#69#,16#69#,16#69#,16#6A#,16#6A#,16#69#,16#68#,16#67#,16#67#,16#67#,16#69#,16#6B#,16#6C#,16#6E#,16#70#,16#57#,16#3C#,16#40#,16#43#,16#4B#,16#4C#,16#47#,16#4C#,16#53#,16#55#,16#69#,16#6B#,16#70#,16#70#,16#6D#,16#6C#,16#6F#,16#6F#,16#68#,16#70#,16#7C#,16#54#,16#69#,16#CD#,16#CA#,16#BF#,16#C9#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CA#,16#CA#,16#CA#,16#C6#,16#CB#,16#CD#,16#CA#,16#CF#,16#C9#,16#CB#,16#CA#,16#CA#,16#BD#,16#B2#,16#AF#,16#AE#,16#AA#,16#A7#,16#A7#,16#A7#,16#A7#,16#A7#,16#A8#,16#A8#,16#A8#,16#AA#,16#A8#,
16#6C#,16#6C#,16#6C#,16#6C#,16#6B#,16#6B#,16#6C#,16#6E#,16#6F#,16#70#,16#71#,16#70#,16#71#,16#69#,16#67#,16#6E#,16#73#,16#4E#,16#4B#,16#A5#,16#A9#,16#92#,16#8F#,16#8D#,16#8E#,16#91#,16#8A#,16#7F#,16#64#,16#5B#,16#4B#,16#49#,16#66#,16#6B#,16#6F#,16#6D#,16#72#,16#6E#,16#7A#,16#5D#,16#3E#,16#AE#,16#D8#,16#B6#,16#C9#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CC#,16#CC#,16#CA#,16#C5#,16#CC#,16#CD#,16#CB#,16#D3#,16#D9#,16#D7#,16#D8#,16#C8#,16#AD#,16#B1#,16#B8#,16#B3#,16#AB#,16#A6#,16#A6#,16#A6#,16#A6#,16#A7#,16#A8#,16#A8#,16#A8#,16#A9#,16#A8#,
16#37#,16#37#,16#36#,16#36#,16#35#,16#35#,16#34#,16#34#,16#38#,16#45#,16#53#,16#52#,16#5F#,16#6A#,16#66#,16#57#,16#37#,16#51#,16#9D#,16#EA#,16#F5#,16#DE#,16#D4#,16#DC#,16#D2#,16#DA#,16#D4#,16#C7#,16#A5#,16#9C#,16#86#,16#74#,16#5F#,16#4D#,16#37#,16#3C#,16#41#,16#44#,16#42#,16#4A#,16#71#,16#B7#,16#D1#,16#C7#,16#CA#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#CD#,16#CD#,16#CB#,16#C4#,16#CD#,16#CD#,16#CC#,16#B0#,16#AF#,16#C9#,16#AC#,16#99#,16#9B#,16#68#,16#7A#,16#BA#,16#AC#,16#A6#,16#A7#,16#A6#,16#A6#,16#A7#,16#A8#,16#A8#,16#A8#,16#A8#,16#A8#,
16#6B#,16#6B#,16#6B#,16#6B#,16#6A#,16#6F#,16#6F#,16#6A#,16#5F#,16#56#,16#56#,16#4D#,16#3F#,16#40#,16#54#,16#67#,16#64#,16#A4#,16#D8#,16#C3#,16#C4#,16#CB#,16#CF#,16#CB#,16#CD#,16#CE#,16#D2#,16#D4#,16#D3#,16#DF#,16#D8#,16#C6#,16#A2#,16#85#,16#6A#,16#61#,16#61#,16#5C#,16#62#,16#8F#,16#CB#,16#CB#,16#CB#,16#CB#,16#CA#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#CE#,16#CE#,16#CB#,16#C4#,16#CC#,16#CB#,16#CC#,16#93#,16#5D#,16#6F#,16#7D#,16#99#,16#A6#,16#6B#,16#4A#,16#A0#,16#B5#,16#A5#,16#A5#,16#A6#,16#A6#,16#A6#,16#A7#,16#A7#,16#A7#,16#A8#,16#A6#,
16#D7#,16#D7#,16#D8#,16#D8#,16#D9#,16#DC#,16#DD#,16#DA#,16#D3#,16#C2#,16#A7#,16#96#,16#7C#,16#6C#,16#88#,16#B3#,16#CF#,16#CF#,16#D0#,16#C4#,16#C7#,16#CB#,16#CB#,16#C9#,16#C8#,16#C9#,16#C9#,16#CA#,16#CA#,16#CC#,16#CD#,16#CB#,16#DF#,16#E0#,16#DA#,16#D5#,16#C6#,16#BF#,16#C9#,16#D6#,16#C9#,16#C9#,16#C9#,16#C9#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#CF#,16#CF#,16#CB#,16#C4#,16#CC#,16#CB#,16#CA#,16#85#,16#2A#,16#43#,16#AD#,16#BE#,16#7F#,16#94#,16#8C#,16#68#,16#AE#,16#AD#,16#A3#,16#A6#,16#A7#,16#A7#,16#A8#,16#A8#,16#A8#,16#A8#,16#A6#,
16#E0#,16#E0#,16#DF#,16#DF#,16#DE#,16#DB#,16#DB#,16#DD#,16#DE#,16#DE#,16#D6#,16#D6#,16#E2#,16#D9#,16#D4#,16#D9#,16#E6#,16#EA#,16#DD#,16#D5#,16#CD#,16#C9#,16#C9#,16#C8#,16#C9#,16#C7#,16#C5#,16#C4#,16#C3#,16#C1#,16#C6#,16#CB#,16#D8#,16#DC#,16#DC#,16#E0#,16#DE#,16#D7#,16#DE#,16#D4#,16#C7#,16#C7#,16#C8#,16#C9#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#CF#,16#CF#,16#CB#,16#C5#,16#C8#,16#CF#,16#C9#,16#7A#,16#2F#,16#5A#,16#D2#,16#BF#,16#66#,16#87#,16#AA#,16#68#,16#A2#,16#B7#,16#9F#,16#A7#,16#A8#,16#A8#,16#A8#,16#A8#,16#A8#,16#A8#,16#A6#,
16#C5#,16#C5#,16#C5#,16#C5#,16#C6#,16#C1#,16#C1#,16#C6#,16#C3#,16#CC#,16#CC#,16#D5#,16#E1#,16#E5#,16#DC#,16#CF#,16#CE#,16#DC#,16#C9#,16#BA#,16#D1#,16#C9#,16#C5#,16#C7#,16#CC#,16#CA#,16#C7#,16#C4#,16#C4#,16#C5#,16#C6#,16#C6#,16#C5#,16#C5#,16#C4#,16#C3#,16#CE#,16#CA#,16#C8#,16#C8#,16#C8#,16#C8#,16#C8#,16#C8#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#D0#,16#D0#,16#CB#,16#C6#,16#C7#,16#CF#,16#C9#,16#CE#,16#B0#,16#85#,16#B7#,16#BE#,16#98#,16#8C#,16#9C#,16#8E#,16#9A#,16#B2#,16#AD#,16#AA#,16#A9#,16#A9#,16#A9#,16#A9#,16#A8#,16#A8#,16#A6#,
16#C4#,16#C4#,16#C4#,16#C5#,16#C5#,16#C5#,16#C6#,16#C6#,16#C1#,16#C6#,16#C6#,16#C0#,16#C3#,16#BD#,16#D2#,16#E0#,16#AB#,16#87#,16#52#,16#5C#,16#CC#,16#D6#,16#C2#,16#C6#,16#BF#,16#C7#,16#C0#,16#C8#,16#C9#,16#C7#,16#C6#,16#C6#,16#C5#,16#C5#,16#C5#,16#C6#,16#C5#,16#C5#,16#C2#,16#CE#,16#C8#,16#C8#,16#C8#,16#C9#,16#C9#,16#CA#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#D0#,16#D0#,16#CB#,16#C5#,16#C8#,16#CE#,16#C8#,16#E6#,16#F4#,16#9D#,16#86#,16#C2#,16#B4#,16#96#,16#99#,16#94#,16#71#,16#98#,16#B7#,16#AB#,16#AA#,16#A9#,16#A9#,16#A9#,16#A8#,16#A6#,16#A5#,
16#C8#,16#C8#,16#C7#,16#C7#,16#C7#,16#C6#,16#C5#,16#C5#,16#C4#,16#C5#,16#C7#,16#C4#,16#CE#,16#E2#,16#BD#,16#95#,16#7B#,16#52#,16#33#,16#5B#,16#CE#,16#D3#,16#C3#,16#C6#,16#C5#,16#CC#,16#E1#,16#E8#,16#D9#,16#D7#,16#DE#,16#E7#,16#F0#,16#EA#,16#EA#,16#D0#,16#C6#,16#C4#,16#C3#,16#CB#,16#C8#,16#C8#,16#C7#,16#C8#,16#C8#,16#C9#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#D0#,16#D0#,16#CB#,16#C5#,16#C8#,16#CD#,16#C9#,16#CA#,16#D1#,16#A7#,16#99#,16#BB#,16#AD#,16#91#,16#95#,16#95#,16#75#,16#7A#,16#A1#,16#B4#,16#AF#,16#A7#,16#A8#,16#AA#,16#A8#,16#A7#,16#A5#,
16#C8#,16#C9#,16#C8#,16#C8#,16#C7#,16#C7#,16#C6#,16#C5#,16#C5#,16#C4#,16#C8#,16#CE#,16#DB#,16#BB#,16#7F#,16#5F#,16#5E#,16#80#,16#76#,16#85#,16#D3#,16#CC#,16#C3#,16#C6#,16#DE#,16#DB#,16#B5#,16#B2#,16#D1#,16#CD#,16#BB#,16#AC#,16#AF#,16#B5#,16#C0#,16#C9#,16#CB#,16#C4#,16#C4#,16#C6#,16#C6#,16#C6#,16#C7#,16#C7#,16#C8#,16#C9#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#D0#,16#D0#,16#CB#,16#C6#,16#C9#,16#CD#,16#C9#,16#D0#,16#AF#,16#94#,16#BC#,16#B4#,16#AA#,16#90#,16#96#,16#9D#,16#9E#,16#89#,16#7C#,16#9E#,16#B3#,16#AF#,16#A6#,16#AB#,16#A8#,16#A7#,16#A5#,
16#C8#,16#C8#,16#C8#,16#C8#,16#C6#,16#C8#,16#C6#,16#C5#,16#C5#,16#C3#,16#C9#,16#D2#,16#B4#,16#6F#,16#69#,16#76#,16#7D#,16#8E#,16#63#,16#94#,16#D5#,16#C9#,16#C4#,16#C6#,16#CC#,16#AC#,16#68#,16#48#,16#92#,16#96#,16#74#,16#4F#,16#53#,16#63#,16#64#,16#A6#,16#CE#,16#C4#,16#C4#,16#C6#,16#C6#,16#C6#,16#C7#,16#C7#,16#C8#,16#C9#,16#CA#,16#CA#,16#CB#,16#CB#,16#CB#,16#CB#,16#CB#,16#D0#,16#D0#,16#CB#,16#C6#,16#C8#,16#CC#,16#CB#,16#CB#,16#97#,16#93#,16#B8#,16#B4#,16#AA#,16#94#,16#9B#,16#98#,16#9D#,16#97#,16#7D#,16#7C#,16#A3#,16#B9#,16#AB#,16#AA#,16#A8#,16#A7#,16#A7#
);

--attribute syn_romstyle : string;
--attribute syn_romstyle of memory : signal is "logic";


begin

  p : process(addr)
	variable vaddr1 : integer range 0 to 6399;
	variable vaddr2 : integer range 0 to 6399;
	variable vaddr3 : integer range 0 to 6399;
	variable vaddr4 : integer range 0 to 6399;
	variable vaddr5 : integer range 0 to 6399;
	variable vaddr6 : integer range 0 to 6399;
	variable vaddr7 : integer range 0 to 6399;
	variable vaddr8 : integer range 0 to 6399;
	begin
			if addr < 800 then
			vaddr1 := To_integer(unsigned(addr&"000"));
			vaddr2 := To_integer(unsigned(addr&"001"));
			vaddr3 := To_integer(unsigned(addr&"010"));
			vaddr4 := To_integer(unsigned(addr&"011"));
			vaddr5 := To_integer(unsigned(addr&"100"));
			vaddr6 := To_integer(unsigned(addr&"101"));
			vaddr7 := To_integer(unsigned(addr&"110"));
			vaddr8 := To_integer(unsigned(addr&"111"));
			end if;
			data_int <= (std_logic_vector(to_unsigned(memory(vaddr1),8)) &  std_logic_vector(to_unsigned(memory(vaddr2),8)) &  std_logic_vector(to_unsigned(memory(vaddr3),8)) & std_logic_vector(to_unsigned(memory(vaddr4),8)) & std_logic_vector(to_unsigned(memory(vaddr5),8)) & std_logic_vector(to_unsigned(memory(vaddr6),8)) & std_logic_vector(to_unsigned(memory(vaddr7),8)) & std_logic_vector(to_unsigned(memory(vaddr8),8)));
		--	data_int(23 downto 16) <= std_logic_vector(to_unsigned(memory(vaddr2),8));
		--	data_int(15 downto 8) <= std_logic_vector(to_unsigned(memory(vaddr3),8));
		--	data_int(7 downto 0) <= std_logic_vector(to_unsigned(memory(vaddr4),8));
  end process;
  
  
  ff: process(clear,clk)
  begin
  	if (clear = '1') then
			data <= (others => '0');    			
	elsif rising_edge(clk) then 
			if (reset = '1') then
			     data <= (others => '0');  
			else 
			     data <= data_int;
 			end if;
 	end if;
  end process;
  




end rtl;
