----------------------------------------------------------------------------------
--
--  This file is a part of Technica Corporation Wizardry Project
--
--  Copyright (C) 2004-2009, Technica Corporation  
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- Module Name: lengthsaver - Behavioral 
-- Project Name: Wizardry
-- Target Devices: Virtex 4 ML401
-- Description: This component calculates the length of each packet.
-- Revision: 1.0
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
USE ieee.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all;
use work.EmPAC_constants.all;

ENTITY lengthsaver IS 
PORT( 
	clock	: IN	std_logic;
	field_data	: IN       std_logic_vector (31 DOWNTO 0);
	length_indicator	: IN       std_logic;
	field_type : IN       std_logic_vector (7 DOWNTO 0);
	reset	: IN       std_logic;
	optional	:	OUT     std_logic;
	length1	: OUT	std_logic_vector (17 DOWNTO 0)
);
END lengthsaver ;
-- VHDL Architecture ProtocolAnalyzer.length_block.struct
-- Generated by Mentor Graphics' HDL Designer(TM) 2003.1 (Build 399)

 

ARCHITECTURE struct OF lengthsaver IS 
-- Architecture declarations 
-- Internal signal declarations
-- SIGNAL IP_header_len	: std_logic_vector(15 DOWNTO 0);
-- SIGNAL opt            : std_logic := '0';
 SIGNAL length1_tmp	: std_logic_vector(17 DOWNTO 0) := (others => '0');
-- signal ip_total_len : std_logic_vector(15 downto 0);
-- signal tcp_header_len : std_logic_vector(15 downto 0);
-- signal no_app_layer : std_logic;
-- signal app_layer_len : std_logic_vector(15 downto 0);
-- signal tcp_head : std_logic_vector(15 downto 0);
-- signal ip_packet_len : std_logic_vector(15 downto 0);
signal IPv4_header_len : std_logic_vector(17 downto 0) := (others => '0');
signal app_layer: std_logic := '0';
signal tcp_header_len : std_logic_Vector(17 downto 0) := (others => '0');
signal transport_layer_len : std_logic_Vector(17 downto 0) := (others => '0');
signal padding : std_logic_Vector(17 downto 0) := (others => '0');
signal total_length : std_logic_Vector(17 downto 0) := (others => '0');
signal IPv6transp_true : std_logic := '1';
signal opt : std_logic := '0';
signal padded : std_logic := '0';
signal pad_data,udp_length : std_logic_vector(17 downto 0) := (others => '0');

BEGIN
 
-- Architecture concurrent statements
 
-- HDL Embedded Text Block	1 len_calc
 
-- The field_type bus indicates what packet field is currently coming
 
-- in on field_data. If the field contains information that will be used to
 
-- calculate a dynamic field length, the information is registered and/or used
 
-- in calculations accordingly.
 --tcp_head <= "0000000000" & tcp_header_len;
-- tcp_head <= "0000000000"&(unsigned(field_data(15 downto 12)) - 5)&"00";

set_len:process(reset,tcp_header_len,field_type,IPv4_header_len,opt,app_layer,clock,transport_layer_len,
					 pad_data)
begin
--if reset = '1' then
--	length1_tmp <= "000000000000000000";

if rising_edge(clock) then
	if reset = '1' then
		length1_tmp <= (others => '0');
	elsif field_type = X"02" then
		length1_tmp <= (others => '0');
	elsif opt = '1' then
		if field_type = X"1C" then
			length1_tmp <= IPv4_header_len - "000000000000010100";--x14,   dec_20 
		elsif field_type = X"29" then
			length1_tmp <= TCP_header_len - "000000000000010100";--x14,    dec_20
		elsif field_type = X"37" then
			length1_tmp <= transport_layer_len;
		elsif field_type = X"30" then
			length1_tmp <= "00"&(unsigned(field_data(15 downto 0)) - 8);
		else
			length1_tmp <= length1_tmp;
		end if;
	elsif app_layer = '1' then
		if field_type = X"29" then
			length1_tmp <= Transport_layer_len - TCP_header_len;
		elsif field_type = X"31" then
--			if padded = '1' then--field_data(15 downto 0) < X"001A" then
--				length1_tmp <= (X"001A" - field_data(15 downto 0)) + ("00"&(unsigned(field_data(15 downto 0)) - 8));
--			else
				length1_tmp <= udp_length + pad_data;
--				length1_tmp <= ("00"&(unsigned(field_data(15 downto 0)) - 8)) + pad_data;--+ padding;--changed 3-26-08
--			end if;
		else
			length1_tmp <= length1_tmp;
		end if;
	elsif opt = '0' and app_layer = '0' then
		if field_type = X"29" then
			length1_tmp <= "000000000000000110";
		elsif field_type = X"31" then
--			if padded = '1' then --field_data(15 downto 0) < X"001A" then
--				length1_tmp <= (X"001A" - field_data(15 downto 0)) + ("00"&(unsigned(field_data(15 downto 0)) - 8));
--			else
				length1_tmp <= udp_length + pad_data;
--				length1_tmp <= ("00"&(unsigned(field_data(15 downto 0)) - 8)) + pad_data;--+ padding;--changed 3-26-08
--			end if;
--			length1_tmp <= "0000000000"&(unsigned(field_data(7 downto 0)) - 8);--original_wrong
		else
			length1_tmp <= length1_tmp;
		end if;
	else
		length1_tmp <= length1_tmp;
	end if;
else
	length1_tmp <= length1_tmp;
end if;
end process;

length1 <= length1_tmp;-- when padded = '0' else 
--			  (length1_tmp + padding) when padded = '1';

process(clock,length_indicator,field_data,field_type)
begin
	if rising_edge(clock) then
		if reset = '1' then
			padded <= '0';
			pad_data <= (others => '0');
			udp_length <= (others => '0');
		else
			if length_indicator = '1' then
				if field_type = X"30" then
					udp_length <= ("00"&(unsigned(field_data(15 downto 0)) - 8));
					if field_data(15 downto 0) < X"001A" then
						padded <= '1';
						pad_data <= "00" & (X"001A" - field_data(15 downto 0));
					else
--						udp_length <= udp_length;
						padded <= '0';
						pad_data <= (others => '0');
					end if;
				elsif field_type = X"17" then
					udp_length <= (others => '0');
					padded <= '0';
					pad_data <= (others => '0');
				else
					udp_length <= udp_length;
					padded <= padded;
					pad_data <= pad_data;
				end if;
			else
				udp_length <= udp_length;
				padded <= padded;
				pad_data <= pad_data;
			end if;
		end if;
	end if;
					
				
end process;


process(clock,reset,length_indicator,field_type)
begin
	if rising_edge(clock) then
		if reset = '1' then
			TCP_header_len <= (others => '0');
		else
			if length_indicator = '1' then
				if field_type = X"17" then
					TCP_header_len <= (others => '0');
				elsif field_type = X"28" then
					TCP_header_len <= "000000000000" & field_data(15 downto 12) & "00";
				else
					TCP_header_len <= TCP_header_len;
				end if;
			else
				TCP_header_len <= TCP_header_len;
			end if;
		end if;
	end if;
end process;


process(clock,reset,length_indicator,field_type)
begin
	if rising_edge(clock) then
		if reset = '1' then
			transport_layer_len <= (others => '0');
		else
			if length_indicator = '1' then
				if field_type = X"17" then
					transport_layer_len <= (others => '0');
				elsif field_type = X"1B" then
					transport_layer_len <= (("00" & field_data(15 downto 0)) - IPv4_header_len);
				elsif field_type = X"36" then
					transport_layer_len <= field_data(15 downto 0) & "00";
				else
					transport_layer_len <= transport_layer_len;
				end if;
			else
				transport_layer_len <= transport_layer_len;
			end if;
		end if;
	end if;
end process;


process(clock,reset,length_indicator,field_type)
begin
	if rising_edge(clock) then
		if reset = '1' then
			IPv4_header_len <= (others => '0');
		else
			if length_indicator = '1' then
				if field_type = X"17" then
					IPv4_header_len <= (others => '0');
				elsif field_type = X"19" then
					IPv4_header_len <= "000000000000" & field_data(3 downto 0) & "00";
				else
					IPv4_header_len <= IPv4_header_len;
				end if;
			else
				IPv4_header_len <= IPv4_header_len;
			end if;
		end if;
	end if;
end process;

process(clock,reset,field_type,field_data)
begin
	if rising_edge(clock) then
		if reset = '1' then
			IPv6transp_true <= '1';
		else
			if field_type = X"37" then
				if ((field_data(7 downto 0) = X"06") or (field_data(7 downto 0) = X"11")) then
					IPv6transp_true <= '1';
				else 	
					IPv6transp_true <= '0';
				end if; 
			elsif field_type = X"17" then
				IPv6transp_true <= '1';
			else
				IPv6transp_true <= IPv6transp_true;
			end if;
		end if;
	end if;
end process;

process(clock,reset,field_type,field_data,length_indicator)
begin
	if rising_edge(clock) then
		if reset = '1' then
			total_length <= (others => '0');
		else
			if field_type = X"1B" then
				Total_length <= (("00" & field_data(15 downto 0)) + X"12"); 
			elsif field_type = X"02" then
				total_length <= (others => '0');
			else
				total_length <= total_length;
			end if;
		end if;
	end if;
end process;

--process(clock,reset,total_length,field_type)
--begin
--	if rising_edge(clock) then
--		if reset = '1' then
--			padded <= '0';
--		else
--			if field_type >= X"1C" then
--				if (total_length < "000000000001000000") then --"X"40") then
--					padded <= '1';
--				else
--					padded <= '0';
--				end if;
--			else
--				padded <= '0';
--			end if;
--		end if;
--	end if;
--end process;


--process(clock,reset,padded)
--begin
--	if rising_edge(clock) then
--		if reset = '1' then
--			padding <= (others => '0');
--		else
--			if padded = '1' then
--				padding <= "000000000001000000" - total_length;
--			else
--				padding <= (others => '0');
--			end if;
--		end if;
--	end if;
--end process;
--transp_len: process(clock,reset,IPv4_header_len,field_type,length_indicator,field_data)
--begin
--if reset = '1' then
----	TCP_header_len <= "000000000000000000";
----	transport_layer_len <= "000000000000000000";
----	IPv4_header_len <= "000000000000000000";
--	IPv6transp_true <= '1';
--elsif rising_edge(clock) then
--	if length_indicator = '1' then
--		if field_type = X"17" then
----			TCP_header_len <= "000000000000000000";
----			transport_layer_len <= "000000000000000000";
----			IPv4_header_len <= "000000000000000000";
--			IPv6transp_true <= '1';
----		elsif field_type = X"19" then
----			IPv4_header_len <= "000000000000" & field_data(3 downto 0) & "00";
----			TCP_header_len <= TCP_header_len;
----			transport_layer_len <= transport_layer_len;
--			IPv6transp_true <= IPv6transp_true;
----		elsif field_type = X"1B" then
----			transport_layer_len <= (("00" & field_data(15 downto 0)) - IPv4_header_len); 
----			IPv4_header_len <= IPv4_header_len;
----			TCP_header_len <= TCP_header_len;
--			IPv6transp_true <= IPv6transp_true;
--		elsif field_type = X"28" then
----			TCP_header_len <= "000000000000" & field_data(15 downto 12) & "00";
----			IPv4_header_len <= IPv4_header_len;
----			transport_layer_len <= transport_layer_len;
--			IPv6transp_true <= IPv6transp_true;
----		elsif field_type = X"36" then
----			transport_layer_len <= field_data(15 downto 0) & "00";
----			IPv4_header_len <= IPv4_header_len;
----			TCP_header_len <= TCP_header_len;
--			IPv6transp_true <= IPv6transp_true;
--		elsif field_type = X"37" then
--			if ((field_data(7 downto 0) = X"06") or (field_data(7 downto 0) = X"11")) then
--				IPv6transp_true <= '1';
--			else 	
--				IPv6transp_true <= '0';
--			end if;
----			transport_layer_len <= transport_layer_len;
----			IPv4_header_len <= IPv4_header_len;
----			TCP_header_len <= TCP_header_len;
--		else
----			IPv4_header_len <= IPv4_header_len;
----			transport_layer_len <= transport_layer_len;
----			TCP_header_len <= TCP_header_len;
--			IPv6transp_true <= IPv6transp_true;
--		end if;
--	else
----		IPv4_header_len <= IPv4_header_len;
----			transport_layer_len <= transport_layer_len;
----			TCP_header_len <= TCP_header_len;
--			IPv6transp_true <= IPv6transp_true;
--	end if;
--else
----	IPv4_header_len <= IPv4_header_len;
----		transport_layer_len <= transport_layer_len;
----		TCP_header_len <= TCP_header_len;
--		IPv6transp_true <= IPv6transp_true;
--end if;
--end process;		

app_lay: process(clock,transport_layer_len,TCP_header_len)
begin
--if rising_edge(clock) then
	if (transport_layer_len - TCP_header_len) > "000000000000000000" then
		app_layer <= '1';
	else
		app_layer <= '0';
	end if;
--end if;
end process;

--app_layer <= '1' when 

options: process(clock,TCP_header_len,IPv4_header_len,IPv6transp_true)
begin
--if rising_edge(clock) then
--	if field_type = X"16" or field_type = X"17" then --X"2B" or field_type = X"22" or field_type = X"40" then
--		opt <= '0';
--	els
	if (((TCP_header_len > "000000000000010100") or (IPv4_header_len > "000000000000010100")) or (IPv6transp_true = '0')) then
		opt <= '1';
--	elsif IPv6transp_true = '1' then
--		opt <= '1';
	else
		opt <= '0';
	end if;
--end if;
end process;
optional <= opt;

END struct; 