-------------------------------------------------------------------------------
-- Title      : LUT to transform HIBI address into mesh address
-- Project    : 
-------------------------------------------------------------------------------
-- File       : addr_lut_example.vhd
-- Author     : 
-- Company    : 
-- Created    : 2006-08-07
-- Last update: 2011-12-01
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: This is an example file that is meant to be copied to somewhere
--              else and edited there. Do not edit this file directly.
-------------------------------------------------------------------------------
-- Copyright (c) 2006 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2006-08-07  1.0      rasmusa Created
-------------------------------------------------------------------------------


-------------------------------------------------------------------------------
-- Funbase IP library Copyright (C) 2011 TUT Department of Computer Systems
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--use ieee.std_logic_arith.all;

-- net_type_g: 0 - 2D MESH
--             1 - Octagon

entity addr_lut is  
  generic (
    in_addr_w_g  : integer := 32;
    out_addr_w_g : integer := 36;
    cmp_high_g   : integer := 31;
    cmp_low_g    : integer := 0;
    net_type_g   : integer := 0;
    lut_en_g     : integer := 1         -- if disabled, out <= in
    );
  port (
    addr_in  : in  std_logic_vector (in_addr_w_g-1 downto 0);
    addr_out : out std_logic_vector (out_addr_w_g-1 downto 0)
    );
end addr_lut;

architecture rtl of addr_lut is

  -- Number of net types
  constant n_net_types_c   : integer := 3;
  constant addr_w_c        : integer := 36;
  constant n_addr_ranges_c : integer := 17;

  
  type addr_rec is record
    in_addr : std_logic_vector (addr_w_c-1 downto 0);
    mask    : std_logic_vector (addr_w_c-1 downto 0);
  end record;
  type address_array is array (0 to n_addr_ranges_c-1) of addr_rec;

  type number_record is record
    x : integer;
    y : integer;
    z : integer;
  end record;
  type number_array is array (0 to n_net_types_c-1, 0 to n_addr_ranges_c-1) of number_record;

  type res_addr_array is array (0 to n_addr_ranges_c-1) of std_logic_vector (out_addr_w_g-1 downto 0);
  
  -- Function for initializing address table
  -- nodes have at most three coordinates (x,y,z)
  -- that are translated differently according to net_type.
  -- All nets do not have 3 coordinates, e.g. 2D-mesh has only 2
  function gen_result_addresses (
    constant numb_arr : number_array;
    constant net_type : integer range 0 to n_net_types_c-1)
    return res_addr_array is
    variable x, y, z : integer;
    variable results : res_addr_array;
  begin  -- gen_addr

    for i in 0 to n_addr_ranges_c-1 loop

      x := numb_arr(net_type, i).x;
      y := numb_arr(net_type, i).y;
      z := numb_arr(net_type, i).z;

      case net_type is

        when 0 =>                       -- MESH: Uses X and Y
          assert out_addr_w_g mod 2 = 0 report "out_addr_w_g must be even" severity failure;
          results(i) := conv_std_logic_vector (x + y*(2**(out_addr_w_g/2)), out_addr_w_g);

        when 1 =>
          results(i) := conv_std_logic_vector (x+y+z, out_addr_w_g);

        when 2 =>
          results(i) := conv_std_logic_vector (z, out_addr_w_g);

          
      end case;

    end loop;  -- i

    return results;
    
  end gen_result_addresses;

  -- Input addresses: received addr is compared against this table.
  constant addr_table_c : address_array :=
    (
      (x"00b000100", x"0ffffff00"),
      (x"00b000300", x"0ffffff00"),
      (x"00b000500", x"0ffffff00"),
      (x"00b000700", x"0ffffff00"),
      
      (x"00b000900", x"1ffffff00"),
      (x"01b000900", x"1ffffff00"),--14.10.06 es, orig value does not fit into integer(x"10b000900", x"1ffffff00"),
      (x"00b000b00", x"0ffffff00"),
      (x"00b000d00", x"0ffffff00"),

      (x"00b000f00", x"0ffffff00"),      
      (x"00b001100", x"0ffffff00"),
      (x"00b001300", x"0ffffff00"),
      (x"00bfffe00", x"0fffffe00"),
      
      (x"009000000", x"0ff000000"),
      (x"00bfedd00", x"0ffffff00"),
      (x"00bfedf00", x"0ffffff00"),
      (x"00bfefd00", x"0ffffff00"),
      
      (x"00bfeff00", x"0ffffff00")
      );

  

  constant num_table_c : number_array :=
    (
      (                                 -- MESH:      
        (0, 0, -1),                     --MASTER     
        (1, 0, -1),                     --Slave1
        (2, 0, -1),                     --Slave2
        (3, 0, -1),                     --Slave3
        (0, 1, -1),                     --Slave4
        (1, 1, -1),                     --Slave5
        (2, 1, -1),                     --Slave6
        (3, 1, -1),                     --Slave7
        (0, 2, -1),                     --Slave8
        (1, 2, -1),                     --Slave9
        (2, 2, -1),                     --SDRAM_msg
        (3, 2, -1),                     --SDRAM_data
        (0, 3, -1),                     --RTM
        (1, 3, -1),                     --ME 2
        (2, 3, -1),                     --ME 1
        (3, 3, -1),                     --dctQidct 2
        (0, 4, -1)                      --dctQidct 1      
        ),
      (                                 -- Octagon:
        (0, 0, 0),                     --MASTER     
        (0, 0, 0),                     --Slave1
        (0, 0, 0),                     --Slave2
        (0, 0, 0),                     --Slave3
        (0, 0, 0),                     --Slave4
        (0, 0, 0),                     --Slave5
        (0, 0, 0),                     --Slave6
        (0, 0, 0),                     --Slave7
        (0, 0, 0),                     --Slave8
        (0, 0, 0),                     --Slave9
        (0, 0, 0),                     --RTM
        (0, 0, 0),                     --SDRAM_msg
        (0, 0, 0),                     --SDRAM_data
        (0, 0, 0),                     --ME 2
        (0, 0, 0),                     --ME 1
        (0, 0, 0),                     --dctQidct 2
        (0, 0, 0)                      --dctQidct 1 
        ),
      (                                 -- Crossbar:
        (0, 0, 0),                      --MASTER     
        (0, 0, 1),                      --Slave1
        (0, 0, 2),                      --Slave2
        (0, 0, 3),                      --Slave3
        (0, 0, 4),                      --Slave4
        (0, 0, 5),                      --Slave5
        (0, 0, 6),                      --Slave6
        (0, 0, 7),                      --Slave7
        (0, 0, 8),                      --Slave8
        (0, 0, 9),                      --Slave9
        (0, 0, 10),                     --RTM
        (0, 0, 11),                     --SDRAM_msg
        (0, 0, 12),                     --SDRAM_data
        (0, 0, 13),                     --ME 2
        (0, 0, 14),                     --ME 1
        (0, 0, 15),                     --dctQidct 2
        (0, 0, 16)                      --dctQidct 1 
        )
      );
  
  constant res_addr_table_c : res_addr_array := gen_result_addresses(num_table_c, net_type_g);

  
begin  -- rtl

  -- Prosessin koodi n�ytt�� ihan j�rkev�lt�.
  -- Kuitenkin jos ulostulo-osoite on _kapeampi_
  -- simulaation k�ynnistys kuolee if-haaraan, johon
  -- ei pit�isi ikin� menn� 8ehto on genericeill�!)
--   cmp_proc : process (addr_in)
--   begin  -- process cmp_proc
--     addr_out <= (others => '0');
--     -- if LUT is disabled
--     if lut_en_g = 0 then
--       if in_addr_w_g > out_addr_w_g then
--         -- Sis��nmeno leve�mpi
--         addr_out                                    <= addr_in(out_addr_w_g-1 downto 0);
--       else
--         -- Ulostulo leve�mpi
--         -- T�� est�� simuloinnin vaikka lut_en_g=1
--         --  Ei voi tajuta. 20.09.2006 es
--         --addr_out (in_addr_w_g-1 downto 0)            <= addr_in(in_addr_w_g-1 downto 0);
--         --addr_out (out_addr_w_g-1 downto in_addr_w_g) <= (others => '0');
--         --assert false report "addr_lut_example: Suurta h�m�ryytt� ilmassa" severity note;
--       end if;
--     else
--       -- if LUT is enabled
--       for i in 0 to n_addr_ranges_c-1 loop
--          if ((addr_in (cmp_high_g downto cmp_low_g)
--               and addr_table_c(i).mask (cmp_high_g downto cmp_low_g))
--               = addr_table_c (i).in_addr (cmp_high_g downto cmp_low_g))
--          then
--            addr_out <= res_addr_table_c(i);
--          end if;
--       end loop;  -- i
--     end if;   
--   end process cmp_proc;


  -- Fix: make tow processes with if-generate
  in_ad_narrower: if in_addr_w_g <= out_addr_w_g generate
    cmp_proc1 : process (addr_in)
    begin  -- process cmp_proc
      addr_out <= (others => '0');

      -- if LUT is disabled
      if lut_en_g = 0 then
          addr_out (out_addr_w_g-1 downto in_addr_w_g) <= (others => '0');
          addr_out (in_addr_w_g-1 downto 0)            <= addr_in(in_addr_w_g-1 downto 0);
          -- The above line was troublesome with regualr if (works with if-generate)
      else
        -- if LUT is enabled

        for i in 0 to n_addr_ranges_c-1 loop
          if ((addr_in (cmp_high_g downto cmp_low_g)
               and addr_table_c(i).mask (cmp_high_g downto cmp_low_g))
              = addr_table_c (i).in_addr (cmp_high_g downto cmp_low_g))
          then
            addr_out <= res_addr_table_c(i);
          end if;
        end loop;  -- i

      end if;
      
    end process cmp_proc1;

  end generate in_ad_narrower;

  

  in_ad_wider: if in_addr_w_g > out_addr_w_g generate
    cmp_proc1 : process (addr_in)
    begin  -- process cmp_proc
      addr_out <= (others => '0');

      -- if LUT is disabled
      if lut_en_g = 0 then
        -- Sis��nmeno leve�mpi
        addr_out <= addr_in(out_addr_w_g-1 downto 0);

      else
        -- if LUT is enabled

        for i in 0 to n_addr_ranges_c-1 loop
          if ((addr_in (cmp_high_g downto cmp_low_g)
               and addr_table_c(i).mask (cmp_high_g downto cmp_low_g))
              = addr_table_c (i).in_addr (cmp_high_g downto cmp_low_g))
          then
            addr_out <= res_addr_table_c(i);
          end if;
        end loop;  -- i

      end if;
      
    end process cmp_proc1;

  end generate in_ad_wider;


  
end rtl;
