// --------------------------------------------------------------------
//
// --------------------------------------------------------------------


module tb_top();

  // --------------------------------------------------------------------
  // test bench clock & reset
  wire clk_50mhz;
  wire tb_clk = clk_50mhz;
  wire tb_rst;

  tb_base #( .PERIOD(20_000) ) tb( clk_50mhz, tb_rst );
  
  
  // --------------------------------------------------------------------
  // 


  // --------------------------------------------------------------------
  // sim models
  //  |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   | 
  // \|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/
  //  '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   ' 



  

  //  '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   ' 
  // /|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\
  //  |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   | 
  // sim models 
  // --------------------------------------------------------------------


  // --------------------------------------------------------------------
  //  debug wires



  // --------------------------------------------------------------------
  // test
  the_test test( tb_clk, tb_rst );

  initial
    begin

      test.run_the_test();

      $display("^^^---------------------------------");
      $display("^^^ %16.t | Testbench done.", $time);
      $display("^^^---------------------------------");

      $display("^^^---------------------------------");

`ifdef MAKEFILE_TEST_RUN
      $finish();
`else
      $stop();
`endif

    end

endmodule



