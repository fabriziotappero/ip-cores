-- Copyright 2015, J�rgen Defurne
--
-- This file is part of the Experimental Unstable CPU System.
--
-- The Experimental Unstable CPU System Is free software: you can redistribute
-- it and/or modify it under the terms of the GNU Lesser General Public License
-- as published by the Free Software Foundation, either version 3 of the
-- License, or (at your option) any later version.
--
-- The Experimental Unstable CPU System is distributed in the hope that it will
-- be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU Lesser
-- General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with Experimental Unstable CPU System. If not, see
-- http://www.gnu.org/licenses/lgpl.txt.


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY dp_000 IS
END dp_000;

ARCHITECTURE behavior OF dp_000 IS

  -- Component Declaration for the Unit Under Test (UUT)
  
  COMPONENT dp
    PORT(
      reset     : IN  STD_LOGIC;
      clock     : IN  STD_LOGIC;
      reg_a     : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
      reg_b     : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
      reg_input : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
      op_sel    : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
      we        : IN  STD_LOGIC;
      pc_input  : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
      pc_load   : IN  STD_LOGIC;
      dr_load   : IN  STD_LOGIC;
      ar_load   : IN  STD_LOGIC;
      aa_load   : IN  STD_LOGIC;
      ab_load   : IN  STD_LOGIC;
      addr_sel  : IN  STD_LOGIC;
      zero      : OUT STD_LOGIC;
      n_zero    : OUT STD_LOGIC;
      data_in   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
      data_out  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
      addr_out  : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
      );
  END COMPONENT;

  -- purpose: Convert a register number into a STD_LOGIC_VECTOR
  FUNCTION reg (reg_nr, len : NATURAL)
    RETURN STD_LOGIC_VECTOR IS
  BEGIN  -- reg
    RETURN STD_LOGIC_VECTOR(to_unsigned(reg_nr, len));
  END reg;


  --Inputs
  -- These two are master signals
  -- There should also be a reset generated by the test code FOR
  -- resetting the data path.
  SIGNAL reset : STD_LOGIC := '0';
  SIGNAL clock : STD_LOGIC := '0';

  SIGNAL dp_rst    : STD_LOGIC                     := '0';
  SIGNAL reg_a     : STD_LOGIC_VECTOR(4 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL reg_b     : STD_LOGIC_VECTOR(4 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL reg_input : STD_LOGIC_VECTOR(1 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL op_sel    : STD_LOGIC_VECTOR(3 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL we        : STD_LOGIC                     := '0';
  SIGNAL pc_input  : STD_LOGIC_VECTOR(1 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL pc_load   : STD_LOGIC                     := '0';
  SIGNAL dr_load   : STD_LOGIC                     := '0';
  SIGNAL ar_load   : STD_LOGIC                     := '0';
  SIGNAL aa_load   : STD_LOGIC                     := '0';
  SIGNAL ab_load   : STD_LOGIC                     := '0';
  SIGNAL addr_sel  : STD_LOGIC                     := '0';
  SIGNAL data_in   : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');

  SIGNAL l_dp_rst    : STD_LOGIC                     := '0';
  SIGNAL l_reg_a     : STD_LOGIC_VECTOR(4 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL l_reg_b     : STD_LOGIC_VECTOR(4 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL l_reg_input : STD_LOGIC_VECTOR(1 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL l_op_sel    : STD_LOGIC_VECTOR(3 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL l_we        : STD_LOGIC                     := '0';
  SIGNAL l_pc_input  : STD_LOGIC_VECTOR(1 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL l_pc_load   : STD_LOGIC                     := '0';
  SIGNAL l_dr_load   : STD_LOGIC                     := '0';
  SIGNAL l_ar_load   : STD_LOGIC                     := '0';
  SIGNAL l_aa_load   : STD_LOGIC                     := '0';
  SIGNAL l_ab_load   : STD_LOGIC                     := '0';
  SIGNAL l_addr_sel  : STD_LOGIC                     := '0';
  SIGNAL l_data_in   : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');

  --Outputs
  SIGNAL zero     : STD_LOGIC;
  SIGNAL n_zero   : STD_LOGIC;
  SIGNAL data_out : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL addr_out : STD_LOGIC_VECTOR(14 DOWNTO 0);

  -- Clock period definitions
  CONSTANT clock_period : TIME := 10 ns;

  SUBTYPE state_range IS NATURAL RANGE 0 TO 104;

  -- State machine definitions
  SIGNAL current : state_range := 0;
  SIGNAL next_s  : state_range := 0;
  
BEGIN

  -- Instantiate the Unit Under Test (UUT)
  uut : dp PORT MAP (
    reset     => dp_rst,
    clock     => clock,
    reg_a     => reg_a,
    reg_b     => reg_b,
    reg_input => reg_input,
    op_sel    => op_sel,
    we        => we,
    pc_input  => pc_input,
    pc_load   => pc_load,
    dr_load   => dr_load,
    ar_load   => ar_load,
    aa_load   => aa_load,
    ab_load   => ab_load,
    addr_sel  => addr_sel,
    zero      => zero,
    n_zero    => n_zero,
    data_in   => data_in,
    data_out  => data_out,
    addr_out  => addr_out
    );

  -- Clock process definitions
  clock_process : PROCESS
  BEGIN
    clock <= '0';
    WAIT FOR clock_period/2;
    clock <= '1';
    WAIT FOR clock_period/2;
  END PROCESS;


  -- Stimulus process
  stim_proc : PROCESS
  BEGIN
    -- hold reset state for 100 ns.
    WAIT FOR 100 ns;
    reset <= '1';
    WAIT FOR clock_period*10;

    -- insert stimulus here 

    IF current = 11 AND next_s = 11 THEN
      WAIT;
    END IF;
  END PROCESS;

  -- purpose: This is the microcontroller pipeline register
  -- type   : sequential
  -- inputs : clock, reset
  -- outputs: reg_a,reg_b,reg_input,op_sel
  pipeline_reg : PROCESS (clock, reset)
  BEGIN  -- PROCESS controller
    IF reset = '0' THEN                 -- asynchronous reset (active low)
      dp_rst    <= '0';
      reg_a     <= (OTHERS => '0');
      reg_b     <= (OTHERS => '0');
      reg_input <= (OTHERS => '0');
      op_sel    <= (OTHERS => '0');
      we        <= '0';
      pc_input  <= (OTHERS => '0');
      pc_load   <= '0';
      dr_load   <= '0';
      ar_load   <= '0';
      aa_load   <= '0';
      ab_load   <= '0';
      addr_sel  <= '0';
      data_in   <= (OTHERS => '0');
      current   <= 0;
    ELSIF rising_edge(clock) THEN       -- rising clock edge
      dp_rst    <= l_dp_rst;
      reg_a     <= l_reg_a;
      reg_b     <= l_reg_b;
      reg_input <= l_reg_input;
      op_sel    <= l_op_sel;
      we        <= l_we;
      pc_input  <= l_pc_input;
      pc_load   <= l_pc_load;
      dr_load   <= l_dr_load;
      ar_load   <= l_ar_load;
      aa_load   <= l_aa_load;
      ab_load   <= l_ab_load;
      addr_sel  <= l_addr_sel;
      data_in   <= l_data_in;
      current   <= next_s;
    END IF;
  END PROCESS pipeline_reg;

  -- purpose: Compute the next state based upon the current state and result zero state
  -- type   : combinational
  -- inputs : current, zero, n_zero
  -- outputs: l_*
  next_state_logic : PROCESS (current, zero, n_zero)
  BEGIN  -- PROCESS next_state_logic

    next_s      <= 0;
    l_dp_rst    <= '1';
    l_reg_a     <= (OTHERS => '0');
    l_reg_b     <= (OTHERS => '0');
    l_reg_input <= (OTHERS => '0');
    l_op_sel    <= (OTHERS => '0');
    l_we        <= '0';
    l_pc_input  <= (OTHERS => '0');
    l_pc_load   <= '0';
    l_dr_load   <= '0';
    l_ar_load   <= '0';
    l_aa_load   <= '0';
    l_ab_load   <= '0';
    l_addr_sel  <= '0';
    l_data_in   <= (OTHERS => '0');

    CASE current IS

      WHEN 0 =>
        next_s   <= 1;
        l_dp_rst <= '0';

      WHEN 1 =>
        next_s      <= 2;
        l_dp_rst    <= '1';
        l_reg_a     <= "00001";
        l_reg_input <= "00";
        l_we        <= '1';
        l_data_in   <= X"F0F0";

      WHEN 2 =>
        next_s     <= 3;
        l_reg_a    <= "00001";
        l_reg_b    <= "00001";
        l_pc_input <= "10";
        l_pc_load  <= '1';
        l_dr_load  <= '1';
        l_ar_load  <= '1';
        l_aa_load  <= '1';
        l_ab_load  <= '1';
        l_addr_sel <= '1';

      WHEN 3 =>
        next_s     <= 4;
        l_addr_sel <= '1';

      WHEN 4 =>
        next_s   <= 5;
        l_dp_rst <= '0';

      WHEN 5 =>
        next_s     <= 6;
        l_data_in  <= X"A1B2";
        l_pc_input <= "01";
        l_pc_load  <= '1';
        l_addr_sel <= '0';

      WHEN 6 =>
        next_s <= 7;

      WHEN 7 =>
        next_s   <= 8;
        l_dp_rst <= '0';

      WHEN 8 =>                         -- Reset state
        next_s      <= 9;
        l_data_in   <= X"DEAD";
        l_reg_input <= "00";
        l_reg_a     <= "00000";
        l_we        <= '1';

      WHEN 9 =>                         -- Present value to register file
        next_s     <= 10;
        l_reg_a    <= "00000";
        l_pc_input <= "10";
        l_pc_load  <= '1';

      WHEN 10 =>  -- Read value from register file into PC
        next_s <= 11;

      WHEN 11 =>
        next_s   <= 12;
        l_dp_rst <= '0';

      WHEN 12 =>                        -- Reset state
        next_s      <= 13;
        l_data_in   <= X"BEEF";
        l_reg_input <= "00";
        l_reg_a     <= "00010";
        l_we        <= '1';

      WHEN 13 =>                        -- Load into register 2
        next_s    <= 14;
        l_reg_a   <= "00010";
        l_dr_load <= '1';

      WHEN 14 =>                        -- Load from register into data out
        next_s <= 15;

      WHEN 15 =>
        next_s   <= 16;
        l_dp_rst <= '0';

      WHEN 16 =>
        next_s      <= 17;
        l_data_in   <= X"FEED";
        l_reg_input <= "00";
        l_reg_a     <= "00011";
        l_we        <= '1';
        
      WHEN 17 =>
        next_s      <= 18;
        l_reg_input <= "11";
        l_reg_a     <= "01111";
        l_reg_b     <= "00011";
        l_we        <= '1';
        
      WHEN 18 =>
        next_s    <= 19;
        l_reg_a   <= "01111";
        l_dr_load <= '1';
        
      WHEN 19 =>
        next_s <= 20;

      WHEN 20 =>                        -- Start AND cycle
        next_s   <= 21;
        l_dp_rst <= '0';
        
      WHEN 21 =>                        -- Reset cycle
        next_s      <= 22;
        l_data_in   <= X"0FA6";
        l_reg_input <= "00";
        l_reg_a     <= "00100";
        l_we        <= '1';

      WHEN 22 =>                        -- Present 0FA6 to register 00100
        next_s      <= 23;
        l_data_in   <= X"FA84";
        l_reg_input <= "00";
        l_reg_a     <= "00101";
        l_we        <= '1';

      WHEN 23 =>                        -- Present FA84 to register 00101
        next_s    <= 24;
        l_reg_a   <= "00100";
        l_reg_b   <= "00101";
        l_aa_load <= '1';
        l_ab_load <= '1';

      WHEN 24 =>                        -- Read reg a and b into A and B
        next_s      <= 25;
        l_reg_input <= "10";
        l_reg_a     <= "00110";
        l_we        <= '1';
        l_op_sel    <= "1010";

      WHEN 25 =>                        -- Perform AND operation, write result
                                        -- into reg 00110
        next_s    <= 26;
        l_reg_a   <= reg(6, 5);
        l_dr_load <= '1';

      WHEN 26 =>                        -- Load reg a into data out register
        next_s <= 27;

      WHEN 27 =>
        next_s   <= 28;
        l_dp_rst <= '0';

      WHEN 28 =>                        -- Reset cycle
        next_s      <= 29;
        l_data_in   <= X"0111";
        l_reg_input <= "00";
        l_reg_a     <= reg(7, 5);
        l_we        <= '1';

      WHEN 29 =>                        -- Present 0111 to register 00111
        next_s      <= 30;
        l_data_in   <= X"0F21";
        l_reg_input <= "00";
        l_reg_a     <= reg(8, 5);
        l_we        <= '1';

      WHEN 30 =>                        -- Present 0F21 to register 01000
        next_s    <= 31;
        l_reg_a   <= reg(7, 5);
        l_reg_b   <= reg(8, 5);
        l_aa_load <= '1';
        l_ab_load <= '1';

      WHEN 31 =>                        -- Read reg a and b into A and B
        next_s      <= 32;
        l_reg_input <= "10";
        l_reg_a     <= reg(9, 5);
        l_we        <= '1';
        l_op_sel    <= "0111";

      WHEN 32 =>                        -- Perform ADD operation, write result
                                        -- into reg 01001
        next_s    <= 33;
        l_reg_a   <= reg(9, 5);
        l_dr_load <= '1';

      WHEN 33 =>                        -- Load reg a into data out register
        next_s <= 34;

      WHEN 34 =>
        next_s   <= 35;
        l_dp_rst <= '0';
        
      WHEN 35 =>                        -- Reset cycle (1)
        next_s      <= 36;
        l_data_in   <= X"7321";
        l_reg_input <= "00";
        l_reg_a     <= reg(10, 5);
        l_we        <= '1';

      WHEN 36 =>                        -- Present X"7321" to register 10 (2)
        next_s      <= 37;
        l_data_in   <= X"6421";
        l_reg_input <= "00";
        l_reg_a     <= reg(11, 5);
        l_we        <= '1';

      WHEN 37 =>                        -- Present X"6421" to register 11 (3)
        next_s    <= 38;
        l_reg_a   <= reg(10, 5);
        l_reg_b   <= reg(11, 5);
        l_aa_load <= '1';
        l_ab_load <= '1';

      WHEN 38 =>                        -- Read reg a and b into A and B (4)
        next_s      <= 39;
        l_reg_input <= "10";
        l_reg_a     <= reg(12, 5);
        l_we        <= '1';
        l_op_sel    <= "1000";

      WHEN 39 =>                        -- Perform ADD operation, write result
                                        -- into reg 12 (5)
        next_s    <= 40;
        l_reg_a   <= reg(12, 5);
        l_dr_load <= '1';

      WHEN 40 =>  -- Load reg a into data out register (6)
        next_s <= 41;

      WHEN 41 =>
        next_s   <= 42;
        l_dp_rst <= '0';
        
      WHEN 42 =>                        -- Reset cycle (1)
        next_s      <= 43;
        l_data_in   <= X"0101";
        l_reg_input <= "00";
        l_reg_a     <= reg(13, 5);
        l_we        <= '1';

      WHEN 43 =>                        -- Present X"0101" to register 13 (2)
        next_s      <= 44;
        l_data_in   <= X"0011";
        l_reg_input <= "00";
        l_reg_a     <= reg(14, 5);
        l_we        <= '1';

      WHEN 44 =>                        -- Present X"0011" to register 14 (3)
        next_s    <= 45;
        l_reg_a   <= reg(13, 5);
        l_reg_b   <= reg(14, 5);
        l_aa_load <= '1';
        l_ab_load <= '1';

      WHEN 45 =>                        -- Read reg a and b into A and B (4)
        next_s      <= 46;
        l_reg_input <= "10";
        l_reg_a     <= reg(15, 5);
        l_we        <= '1';
        l_op_sel    <= "1011";

      WHEN 46 =>                        -- Perform OR operation, write result
                                        -- into reg 15 (5)
        next_s    <= 47;
        l_reg_a   <= reg(15, 5);
        l_dr_load <= '1';

      WHEN 47 =>  -- Load reg a into data out register (6)
        next_s <= 48;

      WHEN 48 =>
        next_s   <= 49;
        l_dp_rst <= '0';
        
      WHEN 49 =>                        -- Reset cycle (1)
        next_s      <= 50;
        l_data_in   <= X"0101";
        l_reg_input <= "00";
        l_reg_a     <= reg(0, 5);
        l_we        <= '1';

      WHEN 50 =>                        -- Present X"0101" to register 0 (2)
        next_s      <= 51;
        l_data_in   <= X"0011";
        l_reg_input <= "00";
        l_reg_a     <= reg(1, 5);
        l_we        <= '1';

      WHEN 51 =>                        -- Present X"0011" to register 1 (3)
        next_s    <= 52;
        l_reg_a   <= reg(0, 5);
        l_reg_b   <= reg(1, 5);
        l_aa_load <= '1';
        l_ab_load <= '1';

      WHEN 52 =>                        -- Read reg a and b into A and B (4)
        next_s      <= 53;
        l_reg_input <= "10";
        l_reg_a     <= reg(2, 5);
        l_we        <= '1';
        l_op_sel    <= "1100";

      WHEN 53 =>                        -- Perform XOR operation, write result
                                        -- into reg 2 (5)
        next_s    <= 54;
        l_reg_a   <= reg(2, 5);
        l_dr_load <= '1';

      WHEN 54 =>  -- Load reg a into data out register (6)
        next_s <= 55;

      WHEN 55 =>
        next_s   <= 56;
        l_dp_rst <= '0';
        
      WHEN 56 =>                        -- Reset cycle (1)
        next_s      <= 57;
        l_data_in   <= X"0A0C";
        l_reg_input <= "00";
        l_reg_a     <= reg(2, 5);
        l_we        <= '1';

      WHEN 57 =>                        -- Present X"0A0C" to register 2 (2)
        next_s    <= 58;
        l_reg_a   <= reg(2, 5);
        l_aa_load <= '1';

      WHEN 58 =>                        -- Read reg a into A (3)
        next_s      <= 59;
        l_reg_input <= "10";
        l_reg_a     <= reg(3, 5);
        l_we        <= '1';
        l_op_sel    <= "1101";

      WHEN 59 =>                        -- Perform NOT operation, write result
                                        -- into reg 3 (4)
        next_s    <= 60;
        l_reg_a   <= reg(3, 5);
        l_dr_load <= '1';

      WHEN 60 =>  -- Load reg a into data out register (5)
        next_s <= 61;

      WHEN 61 =>
        next_s   <= 62;
        l_dp_rst <= '0';

      WHEN 62 =>                        -- Reset cycle (1)
        next_s      <= 63;
        l_data_in   <= X"7310";
        l_reg_input <= "00";
        l_reg_a     <= reg(4, 5);
        l_we        <= '1';

      WHEN 63 =>                        -- Present X"7310" to register 4 (2)
        next_s    <= 64;
        l_reg_a   <= reg(4, 5);
        l_aa_load <= '1';

      WHEN 64 =>                        -- Read reg a into A (3)
        next_s      <= 65;
        l_reg_input <= "10";
        l_reg_a     <= reg(5, 5);
        l_we        <= '1';
        l_op_sel    <= "1110";

      WHEN 65 =>                        -- Perform SLL operation, write result
                                        -- into reg 5 (4)
        next_s    <= 66;
        l_reg_a   <= reg(5, 5);
        l_dr_load <= '1';

      WHEN 66 =>  -- Load reg a into data out register (5)
        next_s <= 67;

      WHEN 67 =>
        next_s   <= 68;
        l_dp_rst <= '0';

      WHEN 68 =>                        -- Reset cycle (1)
        next_s      <= 69;
        l_data_in   <= X"C426";
        l_reg_input <= "00";
        l_reg_a     <= reg(6, 5);
        l_we        <= '1';

      WHEN 69 =>                        -- Present X"C426" to register 6 (2)
        next_s    <= 70;
        l_reg_a   <= reg(6, 5);
        l_aa_load <= '1';

      WHEN 70 =>                        -- Read reg a into A (3)
        next_s      <= 71;
        l_reg_input <= "10";
        l_reg_a     <= reg(7, 5);
        l_we        <= '1';
        l_op_sel    <= "1111";

      WHEN 71 =>                        -- Perform SLL operation, write result
                                        -- into reg 5 (4)
        next_s    <= 72;
        l_reg_a   <= reg(7, 5);
        l_dr_load <= '1';

      WHEN 72 =>  -- Load reg a into data out register (5)
        next_s <= 73;

      WHEN 73 =>
        next_s   <= 74;
        l_dp_rst <= '0';

      WHEN 74 =>                        -- Reset cycle (1)
        next_s      <= 75;
        l_data_in   <= X"001F";
        l_reg_input <= "00";
        l_reg_a     <= reg(8, 5);
        l_we        <= '1';

      WHEN 75 =>                        -- Present X"C426" to register 6 (2)
        next_s    <= 76;
        l_reg_a   <= reg(8, 5);
        l_aa_load <= '1';

      WHEN 76 =>                        -- Read reg a into A (3)
        next_s      <= 77;
        l_reg_input <= "10";
        l_reg_a     <= reg(9, 5);
        l_we        <= '1';
        l_op_sel    <= "0000";

      WHEN 77 =>                        -- Perform INC operation, write result
                                        -- into reg 5 (4)
        next_s    <= 78;
        l_reg_a   <= reg(9, 5);
        l_dr_load <= '1';

      WHEN 78 =>  -- Load reg a into data out register (5)
        next_s <= 79;

      WHEN 79 =>
        next_s   <= 80;
        l_dp_rst <= '0';

      WHEN 80 =>                        -- Reset cycle (1)
        next_s      <= 81;
        l_data_in   <= X"1000";
        l_reg_input <= "00";
        l_reg_a     <= reg(9, 5);
        l_we        <= '1';

      WHEN 81 =>                        -- Present X"1000" to register 9 (2)
        next_s    <= 82;
        l_reg_a   <= reg(9, 5);
        l_aa_load <= '1';

      WHEN 82 =>                        -- Read reg a into A (3)
        next_s      <= 83;
        l_reg_input <= "10";
        l_reg_a     <= reg(10, 5);
        l_we        <= '1';
        l_op_sel    <= "0001";

      WHEN 83 =>                        -- Perform DEC operation, write result
                                        -- into reg 10 (4)
        next_s    <= 84;
        l_reg_a   <= reg(10, 5);
        l_dr_load <= '1';

      WHEN 84 =>  -- Load reg a into data out register (5)
        next_s <= 85;

      WHEN 85 =>
        next_s   <= 86;
        l_dp_rst <= '0';

      WHEN 86 =>                        -- Reset cycle (1)
        next_s     <= 87;
        l_data_in  <= X"1000";
        l_pc_input <= "01";
        l_pc_load  <= '1';

      WHEN 87 =>                        -- Present X"1000" to the program
                                        -- counter (2)
        next_s     <= 88;
        l_pc_input <= "00";
        l_pc_load  <= '1';

      WHEN 88 =>                        -- Reload the program counter
        next_s <= 89;

      WHEN 89 =>
        next_s   <= 90;
        l_dp_rst <= '0';
        
      WHEN 90 =>                        -- Reset cycle (1)
        next_s     <= 91;
        l_data_in  <= X"2000";
        l_pc_input <= "01";
        l_pc_load  <= '1';

      WHEN 91 =>                        -- Present X"2000" to the program
                                        -- counter (2)
        next_s      <= 92;
        l_reg_input <= "01";
        l_reg_a     <= reg(11, 5);
        l_we        <= '1';
        
      WHEN 92 =>                        -- Store PC in register 11
        next_s    <= 93;
        l_reg_a   <= reg(11, 5);
        l_dr_load <= '1';

      WHEN 93 =>                        -- Store reg 11 into data register
        next_s <= 94;

      WHEN 94 =>
        next_s   <= 95;
        l_dp_rst <= '0';

      WHEN 95 =>
        next_s      <= 96;
        l_data_in   <= X"0000";
        l_reg_input <= "00";
        l_reg_a     <= reg(12, 5);
        l_we        <= '1';

      WHEN 96 =>
        next_s  <= 97;
        l_reg_a <= reg(12, 5);

      WHEN 97 =>
        next_s <= 98;

      WHEN 98 =>
        next_s <= 99;

      WHEN 99 =>
        next_s <= 100;
        l_dp_rst <= '0';

      WHEN 100 =>
        next_s      <= 101;
        l_data_in   <= X"0001";
        l_reg_input <= "00";
        l_reg_a     <= reg(13, 5);
        l_we        <= '1';

      WHEN 101 =>
        next_s  <= 102;
        l_reg_a <= reg(13, 5);

      WHEN 102 =>
        next_s <= 103;

      WHEN 103 =>
        next_s <= 104;

      WHEN 104 =>
        next_s <= 104;

    END CASE;
    
  END PROCESS next_state_logic;

  -- purpose: This process checks the values of the data path for every state
  -- type   : sequential
  -- inputs : clock, reset
  -- outputs: 
  assert_tests : PROCESS (clock)
  BEGIN  -- PROCESS assert_tests
    IF rising_edge(clock) THEN          -- rising clock edge
      CASE current IS
        WHEN 1 =>
          ASSERT data_out = X"0000" REPORT "data out register not zero" SEVERITY failure;
          ASSERT addr_out = "111" & X"FF" & X"E" REPORT "address out register not zero" SEVERITY failure;
        WHEN 4 =>
          ASSERT data_out = X"F0F0" REPORT "data out register not F0F0" SEVERITY failure;
          ASSERT addr_out = "111" & X"0F" & X"0" REPORT "address out register not 70F0" SEVERITY failure;
        WHEN 7 =>
          ASSERT addr_out = "010" & X"1B" & X"2" REPORT "address out register not 21B2" SEVERITY failure;
        WHEN 11 =>
          ASSERT addr_out = "101" & X"EA" & X"D" REPORT "address out register not 5EAD" SEVERITY failure;
        WHEN 15 =>
          ASSERT data_out = X"BEEF" REPORT "data out register not BEEF" SEVERITY failure;
        WHEN 20 =>
          ASSERT data_out = X"FEED" REPORT "data out register not FEED" SEVERITY failure;
        WHEN 27 =>
          ASSERT data_out = X"0A84" REPORT "data out register not 0A84" SEVERITY failure;
        WHEN 34 =>
          ASSERT data_out = X"1032" REPORT "data out register not 1032" SEVERITY failure;
        WHEN 41 =>
          ASSERT data_out = X"0F00" REPORT "data out register not 0F00" SEVERITY failure;
        WHEN 48 =>
          ASSERT data_out = X"0111" REPORT "data out register not 0111" SEVERITY failure;
        WHEN 55 =>
          ASSERT data_out = X"0110" REPORT "XOR: data out register not 0110" SEVERITY failure;
        WHEN 61 =>
          ASSERT data_out = X"F5F3" REPORT "NOT: data out register not F5F3" SEVERITY failure;
        WHEN 67 =>
          ASSERT data_out = X"E620" REPORT "SLL: data out register not E620" SEVERITY failure;
        WHEN 73 =>
          ASSERT data_out = X"6213" REPORT "SLR: data out register not 6213" SEVERITY failure;
        WHEN 79 =>
          ASSERT data_out = X"0020" REPORT "INC: data out register not 0020" SEVERITY failure;
        WHEN 85 =>
          ASSERT data_out = X"0FFF" REPORT "DEC: data out register not 0FFF" SEVERITY failure;
        WHEN 89 =>
          ASSERT addr_out = "001000000000001" REPORT "PC-I: address out not 1001" SEVERITY failure;
        WHEN 94 =>
          ASSERT data_out = X"2000" REPORT "PC-II: data out register not 2000" SEVERITY failure;
        WHEN 98 =>
          ASSERT zero = '1' REPORT "TEST-I: zero result not correct" SEVERITY failure;
        WHEN OTHERS => NULL;
      END CASE;
    END IF;
  END PROCESS assert_tests;
END;
