-------------------------------------------------------------------------------
--
-- The Wishbone master module.
--
-- $Id: wb_master-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_wb_master_rtl_c0 of t48_wb_master is

  for rtl
  end for;

end t48_wb_master_rtl_c0;
