module ldpc_edgetable(
  input        clk,
  input        rst,
  input[12:0]  romaddr,
  output[16:0] romdata
);

reg[16:0] romdata_int;

assign romdata = romdata_int;

always @( posedge rst, posedge clk )
  if( rst )
    romdata_int <= 0;
  else
  case( romaddr )
    'h0   : romdata_int = 'h10015; // Pointer for 1_4
    'h1   : romdata_int = 'h101aa; // Pointer for 1_3
    'h2   : romdata_int = 'h1038a; // Pointer for 2_5
    'h3   : romdata_int = 'h105a6; // Pointer for 1_2
    'h4   : romdata_int = 'h107c2; // Pointer for 3_5
    'h5   : romdata_int = 'h10a92; // Pointer for 2_3
    'h6   : romdata_int = 'h10cae; // Pointer for 3_4
    'h7   : romdata_int = 'h10ef7; // Pointer for 4_5
    'h8   : romdata_int = 'h1115b; // Pointer for 5_6
    'h9   : romdata_int = 'h113d1; // Pointer for 8_9
    'ha   : romdata_int = 'h115d9; // Pointer for 9_10
    'hb   : romdata_int = 'h017e3; // Pointer for 1_5s
    'hc   : romdata_int = 'h01846; // Pointer for 1_3s
    'hd   : romdata_int = 'h018be; // Pointer for 2_5s
    'he   : romdata_int = 'h01945; // Pointer for 4_9s
    'hf   : romdata_int = 'h019b3; // Pointer for 3_5s
    'h10  : romdata_int = 'h01a67; // Pointer for 2_3s
    'h11  : romdata_int = 'h01aee; // Pointer for 11_15s
    'h12  : romdata_int = 'h01b66; // Pointer for 7_9s
    'h13  : romdata_int = 'h01bd9; // Pointer for 37_45s
    'h14  : romdata_int = 'h01c5a; // Pointer for 8_9s
    'h15  : romdata_int = 'h187; // Line descriptor for 1_4
    'h16  : romdata_int = 'h4;
    'h17  : romdata_int = 'h3645;
    'h18  : romdata_int = 'h187; // Line descriptor for 1_4
    'h19  : romdata_int = 'h390b;
    'h1a  : romdata_int = 'h58f3;
    'h1b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h1c  : romdata_int = 'hc0e;
    'h1d  : romdata_int = 'h1c14;
    'h1e  : romdata_int = 'h187; // Line descriptor for 1_4
    'h1f  : romdata_int = 'h1b4c;
    'h20  : romdata_int = 'h2945;
    'h21  : romdata_int = 'h187; // Line descriptor for 1_4
    'h22  : romdata_int = 'h27b;
    'h23  : romdata_int = 'h1763;
    'h24  : romdata_int = 'h187; // Line descriptor for 1_4
    'h25  : romdata_int = 'h8c9;
    'h26  : romdata_int = 'h3345;
    'h27  : romdata_int = 'h187; // Line descriptor for 1_4
    'h28  : romdata_int = 'ha67;
    'h29  : romdata_int = 'habd;
    'h2a  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h2b  : romdata_int = 'h1465;
    'h2c  : romdata_int = 'h1937;
    'h2d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h2e  : romdata_int = 'h311e;
    'h2f  : romdata_int = 'h46e2;
    'h30  : romdata_int = 'h187; // Line descriptor for 1_4
    'h31  : romdata_int = 'h222f;
    'h32  : romdata_int = 'h52db;
    'h33  : romdata_int = 'h187; // Line descriptor for 1_4
    'h34  : romdata_int = 'h1338;
    'h35  : romdata_int = 'h143f;
    'h36  : romdata_int = 'h187; // Line descriptor for 1_4
    'h37  : romdata_int = 'h461;
    'h38  : romdata_int = 'h183e;
    'h39  : romdata_int = 'h187; // Line descriptor for 1_4
    'h3a  : romdata_int = 'h10df;
    'h3b  : romdata_int = 'h1ea4;
    'h3c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h3d  : romdata_int = 'h1ced;
    'h3e  : romdata_int = 'h54f3;
    'h3f  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h40  : romdata_int = 'h1690;
    'h41  : romdata_int = 'h3a36;
    'h42  : romdata_int = 'h187; // Line descriptor for 1_4
    'h43  : romdata_int = 'h89;
    'h44  : romdata_int = 'h4e0;
    'h45  : romdata_int = 'h187; // Line descriptor for 1_4
    'h46  : romdata_int = 'h2e;
    'h47  : romdata_int = 'hf48;
    'h48  : romdata_int = 'h187; // Line descriptor for 1_4
    'h49  : romdata_int = 'h1144;
    'h4a  : romdata_int = 'h185c;
    'h4b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h4c  : romdata_int = 'h12ce;
    'h4d  : romdata_int = 'h507e;
    'h4e  : romdata_int = 'h187; // Line descriptor for 1_4
    'h4f  : romdata_int = 'h1135;
    'h50  : romdata_int = 'h18c3;
    'h51  : romdata_int = 'h187; // Line descriptor for 1_4
    'h52  : romdata_int = 'h1746;
    'h53  : romdata_int = 'h3c60;
    'h54  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h55  : romdata_int = 'h1ccb;
    'h56  : romdata_int = 'h2eb3;
    'h57  : romdata_int = 'h187; // Line descriptor for 1_4
    'h58  : romdata_int = 'h2b9;
    'h59  : romdata_int = 'h4711;
    'h5a  : romdata_int = 'h187; // Line descriptor for 1_4
    'h5b  : romdata_int = 'h14c0;
    'h5c  : romdata_int = 'h4838;
    'h5d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h5e  : romdata_int = 'hd4d;
    'h5f  : romdata_int = 'h10d6;
    'h60  : romdata_int = 'h187; // Line descriptor for 1_4
    'h61  : romdata_int = 'haa6;
    'h62  : romdata_int = 'h1b15;
    'h63  : romdata_int = 'h187; // Line descriptor for 1_4
    'h64  : romdata_int = 'h2303;
    'h65  : romdata_int = 'h44b5;
    'h66  : romdata_int = 'h187; // Line descriptor for 1_4
    'h67  : romdata_int = 'h642;
    'h68  : romdata_int = 'h8d5;
    'h69  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h6a  : romdata_int = 'hf2a;
    'h6b  : romdata_int = 'h1d1f;
    'h6c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h6d  : romdata_int = 'h137;
    'h6e  : romdata_int = 'h46b;
    'h6f  : romdata_int = 'h187; // Line descriptor for 1_4
    'h70  : romdata_int = 'hd38;
    'h71  : romdata_int = 'h3c7d;
    'h72  : romdata_int = 'h187; // Line descriptor for 1_4
    'h73  : romdata_int = 'h84a;
    'h74  : romdata_int = 'haf2;
    'h75  : romdata_int = 'h187; // Line descriptor for 1_4
    'h76  : romdata_int = 'h30e5;
    'h77  : romdata_int = 'h48b4;
    'h78  : romdata_int = 'h187; // Line descriptor for 1_4
    'h79  : romdata_int = 'h16b4;
    'h7a  : romdata_int = 'h3307;
    'h7b  : romdata_int = 'h187; // Line descriptor for 1_4
    'h7c  : romdata_int = 'h312;
    'h7d  : romdata_int = 'h10a0;
    'h7e  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h7f  : romdata_int = 'h14e5;
    'h80  : romdata_int = 'h5045;
    'h81  : romdata_int = 'h187; // Line descriptor for 1_4
    'h82  : romdata_int = 'h92b;
    'h83  : romdata_int = 'hcab;
    'h84  : romdata_int = 'h187; // Line descriptor for 1_4
    'h85  : romdata_int = 'h12fd;
    'h86  : romdata_int = 'h299;
    'h87  : romdata_int = 'h187; // Line descriptor for 1_4
    'h88  : romdata_int = 'h728;
    'h89  : romdata_int = 'h36a2;
    'h8a  : romdata_int = 'h187; // Line descriptor for 1_4
    'h8b  : romdata_int = 'h1221;
    'h8c  : romdata_int = 'h266a;
    'h8d  : romdata_int = 'h187; // Line descriptor for 1_4
    'h8e  : romdata_int = 'hb2c;
    'h8f  : romdata_int = 'h4241;
    'h90  : romdata_int = 'h187; // Line descriptor for 1_4
    'h91  : romdata_int = 'h1a64;
    'h92  : romdata_int = 'h1aad;
    'h93  : romdata_int = 'h4187; // Line descriptor for 1_4
    'h94  : romdata_int = 'hb0;
    'h95  : romdata_int = 'h208f;
    'h96  : romdata_int = 'h187; // Line descriptor for 1_4
    'h97  : romdata_int = 'h2a3f;
    'h98  : romdata_int = 'h4a03;
    'h99  : romdata_int = 'h187; // Line descriptor for 1_4
    'h9a  : romdata_int = 'h455;
    'h9b  : romdata_int = 'h121c;
    'h9c  : romdata_int = 'h187; // Line descriptor for 1_4
    'h9d  : romdata_int = 'ha88;
    'h9e  : romdata_int = 'h109b;
    'h9f  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha0  : romdata_int = 'hc25;
    'ha1  : romdata_int = 'h18ca;
    'ha2  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha3  : romdata_int = 'he66;
    'ha4  : romdata_int = 'h2767;
    'ha5  : romdata_int = 'h187; // Line descriptor for 1_4
    'ha6  : romdata_int = 'h167e;
    'ha7  : romdata_int = 'hc4c;
    'ha8  : romdata_int = 'h4187; // Line descriptor for 1_4
    'ha9  : romdata_int = 'h168f;
    'haa  : romdata_int = 'h1b58;
    'hab  : romdata_int = 'h187; // Line descriptor for 1_4
    'hac  : romdata_int = 'h864;
    'had  : romdata_int = 'h3ea6;
    'hae  : romdata_int = 'h187; // Line descriptor for 1_4
    'haf  : romdata_int = 'hf16;
    'hb0  : romdata_int = 'h1a17;
    'hb1  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb2  : romdata_int = 'h936;
    'hb3  : romdata_int = 'h1054;
    'hb4  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb5  : romdata_int = 'h10b;
    'hb6  : romdata_int = 'h1b06;
    'hb7  : romdata_int = 'h187; // Line descriptor for 1_4
    'hb8  : romdata_int = 'h1670;
    'hb9  : romdata_int = 'h2e97;
    'hba  : romdata_int = 'h187; // Line descriptor for 1_4
    'hbb  : romdata_int = 'h2cb1;
    'hbc  : romdata_int = 'h4e6;
    'hbd  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hbe  : romdata_int = 'h2cd5;
    'hbf  : romdata_int = 'h4ac8;
    'hc0  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc1  : romdata_int = 'hc41;
    'hc2  : romdata_int = 'h1319;
    'hc3  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc4  : romdata_int = 'h86;
    'hc5  : romdata_int = 'h4ce8;
    'hc6  : romdata_int = 'h187; // Line descriptor for 1_4
    'hc7  : romdata_int = 'h51e;
    'hc8  : romdata_int = 'h62d;
    'hc9  : romdata_int = 'h187; // Line descriptor for 1_4
    'hca  : romdata_int = 'h8;
    'hcb  : romdata_int = 'he58;
    'hcc  : romdata_int = 'h187; // Line descriptor for 1_4
    'hcd  : romdata_int = 'h161f;
    'hce  : romdata_int = 'h4e10;
    'hcf  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd0  : romdata_int = 'h33b;
    'hd1  : romdata_int = 'h1e3d;
    'hd2  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hd3  : romdata_int = 'h1d3d;
    'hd4  : romdata_int = 'h5280;
    'hd5  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd6  : romdata_int = 'h1a42;
    'hd7  : romdata_int = 'h72c;
    'hd8  : romdata_int = 'h187; // Line descriptor for 1_4
    'hd9  : romdata_int = 'hc75;
    'hda  : romdata_int = 'h173f;
    'hdb  : romdata_int = 'h187; // Line descriptor for 1_4
    'hdc  : romdata_int = 'h1a2b;
    'hdd  : romdata_int = 'h435e;
    'hde  : romdata_int = 'h187; // Line descriptor for 1_4
    'hdf  : romdata_int = 'h1030;
    'he0  : romdata_int = 'h1887;
    'he1  : romdata_int = 'h187; // Line descriptor for 1_4
    'he2  : romdata_int = 'h1623;
    'he3  : romdata_int = 'h4c59;
    'he4  : romdata_int = 'h187; // Line descriptor for 1_4
    'he5  : romdata_int = 'h122a;
    'he6  : romdata_int = 'h4606;
    'he7  : romdata_int = 'h4187; // Line descriptor for 1_4
    'he8  : romdata_int = 'h10d0;
    'he9  : romdata_int = 'h4ca0;
    'hea  : romdata_int = 'h187; // Line descriptor for 1_4
    'heb  : romdata_int = 'h4d5;
    'hec  : romdata_int = 'h3434;
    'hed  : romdata_int = 'h187; // Line descriptor for 1_4
    'hee  : romdata_int = 'h83b;
    'hef  : romdata_int = 'h446f;
    'hf0  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf1  : romdata_int = 'hb22;
    'hf2  : romdata_int = 'he4d;
    'hf3  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf4  : romdata_int = 'h48a;
    'hf5  : romdata_int = 'h862;
    'hf6  : romdata_int = 'h187; // Line descriptor for 1_4
    'hf7  : romdata_int = 'h12c9;
    'hf8  : romdata_int = 'h1522;
    'hf9  : romdata_int = 'h187; // Line descriptor for 1_4
    'hfa  : romdata_int = 'h1958;
    'hfb  : romdata_int = 'h4e85;
    'hfc  : romdata_int = 'h4187; // Line descriptor for 1_4
    'hfd  : romdata_int = 'h18db;
    'hfe  : romdata_int = 'ha5c;
    'hff  : romdata_int = 'h187; // Line descriptor for 1_4
    'h100 : romdata_int = 'h1d1d;
    'h101 : romdata_int = 'h346f;
    'h102 : romdata_int = 'h187; // Line descriptor for 1_4
    'h103 : romdata_int = 'h168c;
    'h104 : romdata_int = 'h4e08;
    'h105 : romdata_int = 'h187; // Line descriptor for 1_4
    'h106 : romdata_int = 'h954;
    'h107 : romdata_int = 'hd52;
    'h108 : romdata_int = 'h187; // Line descriptor for 1_4
    'h109 : romdata_int = 'h16da;
    'h10a : romdata_int = 'h22f8;
    'h10b : romdata_int = 'h187; // Line descriptor for 1_4
    'h10c : romdata_int = 'h24dc;
    'h10d : romdata_int = 'h4049;
    'h10e : romdata_int = 'h187; // Line descriptor for 1_4
    'h10f : romdata_int = 'h673;
    'h110 : romdata_int = 'hb49;
    'h111 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h112 : romdata_int = 'h279;
    'h113 : romdata_int = 'h3eaf;
    'h114 : romdata_int = 'h187; // Line descriptor for 1_4
    'h115 : romdata_int = 'h1006;
    'h116 : romdata_int = 'h4149;
    'h117 : romdata_int = 'h187; // Line descriptor for 1_4
    'h118 : romdata_int = 'h890;
    'h119 : romdata_int = 'h10be;
    'h11a : romdata_int = 'h187; // Line descriptor for 1_4
    'h11b : romdata_int = 'hef3;
    'h11c : romdata_int = 'h303c;
    'h11d : romdata_int = 'h187; // Line descriptor for 1_4
    'h11e : romdata_int = 'h2b8;
    'h11f : romdata_int = 'h4a5;
    'h120 : romdata_int = 'h187; // Line descriptor for 1_4
    'h121 : romdata_int = 'h187b;
    'h122 : romdata_int = 'h9a;
    'h123 : romdata_int = 'h187; // Line descriptor for 1_4
    'h124 : romdata_int = 'h1031;
    'h125 : romdata_int = 'h1845;
    'h126 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h127 : romdata_int = 'h302;
    'h128 : romdata_int = 'h3857;
    'h129 : romdata_int = 'h187; // Line descriptor for 1_4
    'h12a : romdata_int = 'h3b26;
    'h12b : romdata_int = 'h4a22;
    'h12c : romdata_int = 'h187; // Line descriptor for 1_4
    'h12d : romdata_int = 'h24da;
    'h12e : romdata_int = 'h5555;
    'h12f : romdata_int = 'h187; // Line descriptor for 1_4
    'h130 : romdata_int = 'h18ee;
    'h131 : romdata_int = 'h6e5;
    'h132 : romdata_int = 'h187; // Line descriptor for 1_4
    'h133 : romdata_int = 'h24e4;
    'h134 : romdata_int = 'h52b5;
    'h135 : romdata_int = 'h187; // Line descriptor for 1_4
    'h136 : romdata_int = 'h1906;
    'h137 : romdata_int = 'h1eb3;
    'h138 : romdata_int = 'h187; // Line descriptor for 1_4
    'h139 : romdata_int = 'h1c9a;
    'h13a : romdata_int = 'h2af5;
    'h13b : romdata_int = 'h4187; // Line descriptor for 1_4
    'h13c : romdata_int = 'hf58;
    'h13d : romdata_int = 'h2644;
    'h13e : romdata_int = 'h187; // Line descriptor for 1_4
    'h13f : romdata_int = 'h467;
    'h140 : romdata_int = 'h1308;
    'h141 : romdata_int = 'h187; // Line descriptor for 1_4
    'h142 : romdata_int = 'h6a7;
    'h143 : romdata_int = 'h1418;
    'h144 : romdata_int = 'h187; // Line descriptor for 1_4
    'h145 : romdata_int = 'he1a;
    'h146 : romdata_int = 'h3e52;
    'h147 : romdata_int = 'h187; // Line descriptor for 1_4
    'h148 : romdata_int = 'h1a35;
    'h149 : romdata_int = 'h5898;
    'h14a : romdata_int = 'h187; // Line descriptor for 1_4
    'h14b : romdata_int = 'h27f;
    'h14c : romdata_int = 'h14eb;
    'h14d : romdata_int = 'h187; // Line descriptor for 1_4
    'h14e : romdata_int = 'hd5;
    'h14f : romdata_int = 'hb27;
    'h150 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h151 : romdata_int = 'h3628;
    'h152 : romdata_int = 'h511e;
    'h153 : romdata_int = 'h187; // Line descriptor for 1_4
    'h154 : romdata_int = 'h14fd;
    'h155 : romdata_int = 'h3af9;
    'h156 : romdata_int = 'h187; // Line descriptor for 1_4
    'h157 : romdata_int = 'h1d31;
    'h158 : romdata_int = 'h1440;
    'h159 : romdata_int = 'h187; // Line descriptor for 1_4
    'h15a : romdata_int = 'h15c;
    'h15b : romdata_int = 'hd4f;
    'h15c : romdata_int = 'h187; // Line descriptor for 1_4
    'h15d : romdata_int = 'h8b6;
    'h15e : romdata_int = 'h38f3;
    'h15f : romdata_int = 'h187; // Line descriptor for 1_4
    'h160 : romdata_int = 'h1cc4;
    'h161 : romdata_int = 'h5959;
    'h162 : romdata_int = 'h187; // Line descriptor for 1_4
    'h163 : romdata_int = 'hc8f;
    'h164 : romdata_int = 'h1408;
    'h165 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h166 : romdata_int = 'h2e1d;
    'h167 : romdata_int = 'h5711;
    'h168 : romdata_int = 'h187; // Line descriptor for 1_4
    'h169 : romdata_int = 'h1233;
    'h16a : romdata_int = 'hc70;
    'h16b : romdata_int = 'h187; // Line descriptor for 1_4
    'h16c : romdata_int = 'h67c;
    'h16d : romdata_int = 'h6a4;
    'h16e : romdata_int = 'h187; // Line descriptor for 1_4
    'h16f : romdata_int = 'h1250;
    'h170 : romdata_int = 'h281e;
    'h171 : romdata_int = 'h187; // Line descriptor for 1_4
    'h172 : romdata_int = 'hae;
    'h173 : romdata_int = 'h40ff;
    'h174 : romdata_int = 'h187; // Line descriptor for 1_4
    'h175 : romdata_int = 'h29b;
    'h176 : romdata_int = 'h1a73;
    'h177 : romdata_int = 'h187; // Line descriptor for 1_4
    'h178 : romdata_int = 'h27c;
    'h179 : romdata_int = 'h145d;
    'h17a : romdata_int = 'h4187; // Line descriptor for 1_4
    'h17b : romdata_int = 'h40d;
    'h17c : romdata_int = 'h1c0a;
    'h17d : romdata_int = 'h187; // Line descriptor for 1_4
    'h17e : romdata_int = 'h2afe;
    'h17f : romdata_int = 'h5687;
    'h180 : romdata_int = 'h187; // Line descriptor for 1_4
    'h181 : romdata_int = 'h147b;
    'h182 : romdata_int = 'h3551;
    'h183 : romdata_int = 'h187; // Line descriptor for 1_4
    'h184 : romdata_int = 'h6a6;
    'h185 : romdata_int = 'h4550;
    'h186 : romdata_int = 'h187; // Line descriptor for 1_4
    'h187 : romdata_int = 'h2049;
    'h188 : romdata_int = 'h5696;
    'h189 : romdata_int = 'h187; // Line descriptor for 1_4
    'h18a : romdata_int = 'heee;
    'h18b : romdata_int = 'h54e5;
    'h18c : romdata_int = 'h187; // Line descriptor for 1_4
    'h18d : romdata_int = 'h1cc9;
    'h18e : romdata_int = 'h2ca6;
    'h18f : romdata_int = 'h4187; // Line descriptor for 1_4
    'h190 : romdata_int = 'h8f2;
    'h191 : romdata_int = 'h2919;
    'h192 : romdata_int = 'h187; // Line descriptor for 1_4
    'h193 : romdata_int = 'h20cd;
    'h194 : romdata_int = 'h3cdd;
    'h195 : romdata_int = 'h187; // Line descriptor for 1_4
    'h196 : romdata_int = 'hb01;
    'h197 : romdata_int = 'h1ac5;
    'h198 : romdata_int = 'h187; // Line descriptor for 1_4
    'h199 : romdata_int = 'h1d5b;
    'h19a : romdata_int = 'h329e;
    'h19b : romdata_int = 'h187; // Line descriptor for 1_4
    'h19c : romdata_int = 'he0a;
    'h19d : romdata_int = 'h4267;
    'h19e : romdata_int = 'h187; // Line descriptor for 1_4
    'h19f : romdata_int = 'h643;
    'h1a0 : romdata_int = 'ha48;
    'h1a1 : romdata_int = 'h187; // Line descriptor for 1_4
    'h1a2 : romdata_int = 'h6b0;
    'h1a3 : romdata_int = 'h12a2;
    'h1a4 : romdata_int = 'h4187; // Line descriptor for 1_4
    'h1a5 : romdata_int = 'h238;
    'h1a6 : romdata_int = 'he32;
    'h1a7 : romdata_int = 'h2187; // Line descriptor for 1_4
    'h1a8 : romdata_int = 'h528;
    'h1a9 : romdata_int = 'h4862;
    'h1aa : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ab : romdata_int = 'h2e;
    'h1ac : romdata_int = 'hb0;
    'h1ad : romdata_int = 'h5939;
    'h1ae : romdata_int = 'h278; // Line descriptor for 1_3
    'h1af : romdata_int = 'h46e4;
    'h1b0 : romdata_int = 'h5cb8;
    'h1b1 : romdata_int = 'h6cec;
    'h1b2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1b3 : romdata_int = 'hc8f;
    'h1b4 : romdata_int = 'h20f3;
    'h1b5 : romdata_int = 'h371c;
    'h1b6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1b7 : romdata_int = 'h27b;
    'h1b8 : romdata_int = 'h194c;
    'h1b9 : romdata_int = 'h5cd1;
    'h1ba : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1bb : romdata_int = 'h1563;
    'h1bc : romdata_int = 'h1a14;
    'h1bd : romdata_int = 'h2f59;
    'h1be : romdata_int = 'h278; // Line descriptor for 1_3
    'h1bf : romdata_int = 'h8c9;
    'h1c0 : romdata_int = 'h2256;
    'h1c1 : romdata_int = 'h2410;
    'h1c2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1c3 : romdata_int = 'ha67;
    'h1c4 : romdata_int = 'habd;
    'h1c5 : romdata_int = 'h1f07;
    'h1c6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1c7 : romdata_int = 'h1265;
    'h1c8 : romdata_int = 'h2480;
    'h1c9 : romdata_int = 'h5e43;
    'h1ca : romdata_int = 'h278; // Line descriptor for 1_3
    'h1cb : romdata_int = 'h2a91;
    'h1cc : romdata_int = 'h2c85;
    'h1cd : romdata_int = 'h454a;
    'h1ce : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1cf : romdata_int = 'h1321;
    'h1d0 : romdata_int = 'h2036;
    'h1d1 : romdata_int = 'h2ee3;
    'h1d2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1d3 : romdata_int = 'h461;
    'h1d4 : romdata_int = 'h26b1;
    'h1d5 : romdata_int = 'h5b07;
    'h1d6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1d7 : romdata_int = 'h206c;
    'h1d8 : romdata_int = 'h1138;
    'h1d9 : romdata_int = 'h123f;
    'h1da : romdata_int = 'h278; // Line descriptor for 1_3
    'h1db : romdata_int = 'h1c97;
    'h1dc : romdata_int = 'h6c29;
    'h1dd : romdata_int = 'h2137;
    'h1de : romdata_int = 'h278; // Line descriptor for 1_3
    'h1df : romdata_int = 'h86;
    'h1e0 : romdata_int = 'h163e;
    'h1e1 : romdata_int = 'h1490;
    'h1e2 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1e3 : romdata_int = 'h2d43;
    'h1e4 : romdata_int = 'h4e0;
    'h1e5 : romdata_int = 'h89;
    'h1e6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1e7 : romdata_int = 'hf48;
    'h1e8 : romdata_int = 'h165c;
    'h1e9 : romdata_int = 'h5877;
    'h1ea : romdata_int = 'h278; // Line descriptor for 1_3
    'h1eb : romdata_int = 'h2206;
    'h1ec : romdata_int = 'h680a;
    'h1ed : romdata_int = 'h7242;
    'h1ee : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ef : romdata_int = 'h1aed;
    'h1f0 : romdata_int = 'h44b0;
    'h1f1 : romdata_int = 'h46f5;
    'h1f2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h1f3 : romdata_int = 'hf05;
    'h1f4 : romdata_int = 'h10ce;
    'h1f5 : romdata_int = 'h7458;
    'h1f6 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h1f7 : romdata_int = 'h1546;
    'h1f8 : romdata_int = 'h2ced;
    'h1f9 : romdata_int = 'h5cd3;
    'h1fa : romdata_int = 'h278; // Line descriptor for 1_3
    'h1fb : romdata_int = 'h1c3f;
    'h1fc : romdata_int = 'h414c;
    'h1fd : romdata_int = 'h1461;
    'h1fe : romdata_int = 'h278; // Line descriptor for 1_3
    'h1ff : romdata_int = 'hb53;
    'h200 : romdata_int = 'h16c3;
    'h201 : romdata_int = 'h20ee;
    'h202 : romdata_int = 'h278; // Line descriptor for 1_3
    'h203 : romdata_int = 'h2b9;
    'h204 : romdata_int = 'hea1;
    'h205 : romdata_int = 'h1915;
    'h206 : romdata_int = 'h278; // Line descriptor for 1_3
    'h207 : romdata_int = 'h642;
    'h208 : romdata_int = 'h2249;
    'h209 : romdata_int = 'h3a94;
    'h20a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h20b : romdata_int = 'h12c0;
    'h20c : romdata_int = 'h4aa0;
    'h20d : romdata_int = 'h569b;
    'h20e : romdata_int = 'h278; // Line descriptor for 1_3
    'h20f : romdata_int = 'hc25;
    'h210 : romdata_int = 'h1e9e;
    'h211 : romdata_int = 'h24ee;
    'h212 : romdata_int = 'h278; // Line descriptor for 1_3
    'h213 : romdata_int = 'h4;
    'h214 : romdata_int = 'haa6;
    'h215 : romdata_int = 'h10fe;
    'h216 : romdata_int = 'h278; // Line descriptor for 1_3
    'h217 : romdata_int = 'h46b;
    'h218 : romdata_int = 'hf2a;
    'h219 : romdata_int = 'h6e22;
    'h21a : romdata_int = 'h278; // Line descriptor for 1_3
    'h21b : romdata_int = 'h8d5;
    'h21c : romdata_int = 'h2260;
    'h21d : romdata_int = 'h7343;
    'h21e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h21f : romdata_int = 'h1abb;
    'h220 : romdata_int = 'h28eb;
    'h221 : romdata_int = 'h52d6;
    'h222 : romdata_int = 'h278; // Line descriptor for 1_3
    'h223 : romdata_int = 'h312;
    'h224 : romdata_int = 'hd52;
    'h225 : romdata_int = 'h2091;
    'h226 : romdata_int = 'h278; // Line descriptor for 1_3
    'h227 : romdata_int = 'h92b;
    'h228 : romdata_int = 'h1b1f;
    'h229 : romdata_int = 'h774b;
    'h22a : romdata_int = 'h278; // Line descriptor for 1_3
    'h22b : romdata_int = 'haf2;
    'h22c : romdata_int = 'hc0e;
    'h22d : romdata_int = 'h273b;
    'h22e : romdata_int = 'h278; // Line descriptor for 1_3
    'h22f : romdata_int = 'h4205;
    'h230 : romdata_int = 'h608e;
    'h231 : romdata_int = 'h76d3;
    'h232 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h233 : romdata_int = 'h728;
    'h234 : romdata_int = 'h3167;
    'h235 : romdata_int = 'h6b66;
    'h236 : romdata_int = 'h278; // Line descriptor for 1_3
    'h237 : romdata_int = 'hb2c;
    'h238 : romdata_int = 'h1e39;
    'h239 : romdata_int = 'h1e8b;
    'h23a : romdata_int = 'h278; // Line descriptor for 1_3
    'h23b : romdata_int = 'h247e;
    'h23c : romdata_int = 'h5162;
    'h23d : romdata_int = 'h68d2;
    'h23e : romdata_int = 'h278; // Line descriptor for 1_3
    'h23f : romdata_int = 'h101c;
    'h240 : romdata_int = 'h10fd;
    'h241 : romdata_int = 'h3274;
    'h242 : romdata_int = 'h278; // Line descriptor for 1_3
    'h243 : romdata_int = 'h9a;
    'h244 : romdata_int = 'hd4f;
    'h245 : romdata_int = 'h12e5;
    'h246 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h247 : romdata_int = 'h16ca;
    'h248 : romdata_int = 'h1cfc;
    'h249 : romdata_int = 'h1cfe;
    'h24a : romdata_int = 'h278; // Line descriptor for 1_3
    'h24b : romdata_int = 'h147e;
    'h24c : romdata_int = 'h18ad;
    'h24d : romdata_int = 'h2430;
    'h24e : romdata_int = 'h278; // Line descriptor for 1_3
    'h24f : romdata_int = 'h455;
    'h250 : romdata_int = 'h200e;
    'h251 : romdata_int = 'h6a48;
    'h252 : romdata_int = 'h278; // Line descriptor for 1_3
    'h253 : romdata_int = 'he66;
    'h254 : romdata_int = 'h2458;
    'h255 : romdata_int = 'h7622;
    'h256 : romdata_int = 'h278; // Line descriptor for 1_3
    'h257 : romdata_int = 'h864;
    'h258 : romdata_int = 'h1817;
    'h259 : romdata_int = 'h1d38;
    'h25a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h25b : romdata_int = 'h24b5;
    'h25c : romdata_int = 'h3d4c;
    'h25d : romdata_int = 'h6052;
    'h25e : romdata_int = 'h278; // Line descriptor for 1_3
    'h25f : romdata_int = 'ha88;
    'h260 : romdata_int = 'h160b;
    'h261 : romdata_int = 'h5887;
    'h262 : romdata_int = 'h278; // Line descriptor for 1_3
    'h263 : romdata_int = 'h1470;
    'h264 : romdata_int = 'h1ee5;
    'h265 : romdata_int = 'h4e13;
    'h266 : romdata_int = 'h278; // Line descriptor for 1_3
    'h267 : romdata_int = 'hae;
    'h268 : romdata_int = 'h2238;
    'h269 : romdata_int = 'h647b;
    'h26a : romdata_int = 'h278; // Line descriptor for 1_3
    'h26b : romdata_int = 'h1958;
    'h26c : romdata_int = 'h24a8;
    'h26d : romdata_int = 'h7424;
    'h26e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h26f : romdata_int = 'h491;
    'h270 : romdata_int = 'hf16;
    'h271 : romdata_int = 'h6d1d;
    'h272 : romdata_int = 'h278; // Line descriptor for 1_3
    'h273 : romdata_int = 'h2057;
    'h274 : romdata_int = 'h1842;
    'h275 : romdata_int = 'h2465;
    'h276 : romdata_int = 'h278; // Line descriptor for 1_3
    'h277 : romdata_int = 'hd5;
    'h278 : romdata_int = 'h1b3d;
    'h279 : romdata_int = 'h20f4;
    'h27a : romdata_int = 'h278; // Line descriptor for 1_3
    'h27b : romdata_int = 'h51e;
    'h27c : romdata_int = 'h1e3c;
    'h27d : romdata_int = 'h3633;
    'h27e : romdata_int = 'h278; // Line descriptor for 1_3
    'h27f : romdata_int = 'h10b;
    'h280 : romdata_int = 'h936;
    'h281 : romdata_int = 'h26d4;
    'h282 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h283 : romdata_int = 'h3a54;
    'h284 : romdata_int = 'h4af2;
    'h285 : romdata_int = 'h6486;
    'h286 : romdata_int = 'h278; // Line descriptor for 1_3
    'h287 : romdata_int = 'h1119;
    'h288 : romdata_int = 'h1687;
    'h289 : romdata_int = 'h182b;
    'h28a : romdata_int = 'h278; // Line descriptor for 1_3
    'h28b : romdata_int = 'h72c;
    'h28c : romdata_int = 'h33b;
    'h28d : romdata_int = 'h5747;
    'h28e : romdata_int = 'h278; // Line descriptor for 1_3
    'h28f : romdata_int = 'hcab;
    'h290 : romdata_int = 'h1706;
    'h291 : romdata_int = 'h62d;
    'h292 : romdata_int = 'h278; // Line descriptor for 1_3
    'h293 : romdata_int = 'h141f;
    'h294 : romdata_int = 'h22d8;
    'h295 : romdata_int = 'h649b;
    'h296 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h297 : romdata_int = 'h28cf;
    'h298 : romdata_int = 'h3229;
    'h299 : romdata_int = 'h4818;
    'h29a : romdata_int = 'h278; // Line descriptor for 1_3
    'h29b : romdata_int = 'h1f66;
    'h29c : romdata_int = 'h1f4d;
    'h29d : romdata_int = 'h102a;
    'h29e : romdata_int = 'h278; // Line descriptor for 1_3
    'h29f : romdata_int = 'h1e81;
    'h2a0 : romdata_int = 'h391c;
    'h2a1 : romdata_int = 'he4d;
    'h2a2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2a3 : romdata_int = 'h4d5;
    'h2a4 : romdata_int = 'h223a;
    'h2a5 : romdata_int = 'h6ace;
    'h2a6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2a7 : romdata_int = 'h83b;
    'h2a8 : romdata_int = 'hb22;
    'h2a9 : romdata_int = 'h153f;
    'h2aa : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2ab : romdata_int = 'h48a;
    'h2ac : romdata_int = 'h4e70;
    'h2ad : romdata_int = 'h6712;
    'h2ae : romdata_int = 'h278; // Line descriptor for 1_3
    'h2af : romdata_int = 'h1423;
    'h2b0 : romdata_int = 'h2ee4;
    'h2b1 : romdata_int = 'h3a7a;
    'h2b2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2b3 : romdata_int = 'ha5c;
    'h2b4 : romdata_int = 'h1758;
    'h2b5 : romdata_int = 'h1f1e;
    'h2b6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2b7 : romdata_int = 'h862;
    'h2b8 : romdata_int = 'h148c;
    'h2b9 : romdata_int = 'h26f3;
    'h2ba : romdata_int = 'h278; // Line descriptor for 1_3
    'h2bb : romdata_int = 'h10c9;
    'h2bc : romdata_int = 'h167b;
    'h2bd : romdata_int = 'h7078;
    'h2be : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2bf : romdata_int = 'h14da;
    'h2c0 : romdata_int = 'h1f45;
    'h2c1 : romdata_int = 'h3157;
    'h2c2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2c3 : romdata_int = 'h954;
    'h2c4 : romdata_int = 'h16db;
    'h2c5 : romdata_int = 'h1d45;
    'h2c6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2c7 : romdata_int = 'h2203;
    'h2c8 : romdata_int = 'h2445;
    'h2c9 : romdata_int = 'h40f2;
    'h2ca : romdata_int = 'h278; // Line descriptor for 1_3
    'h2cb : romdata_int = 'h852;
    'h2cc : romdata_int = 'h3523;
    'h2cd : romdata_int = 'h4317;
    'h2ce : romdata_int = 'h278; // Line descriptor for 1_3
    'h2cf : romdata_int = 'h673;
    'h2d0 : romdata_int = 'h1c1e;
    'h2d1 : romdata_int = 'h246e;
    'h2d2 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2d3 : romdata_int = 'h279;
    'h2d4 : romdata_int = 'hd4d;
    'h2d5 : romdata_int = 'h1645;
    'h2d6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2d7 : romdata_int = 'h6f3;
    'h2d8 : romdata_int = 'h22b4;
    'h2d9 : romdata_int = 'h60a6;
    'h2da : romdata_int = 'h278; // Line descriptor for 1_3
    'h2db : romdata_int = 'h4ccb;
    'h2dc : romdata_int = 'hb49;
    'h2dd : romdata_int = 'hef3;
    'h2de : romdata_int = 'h278; // Line descriptor for 1_3
    'h2df : romdata_int = 'h70b8;
    'h2e0 : romdata_int = 'h4a2c;
    'h2e1 : romdata_int = 'h4cee;
    'h2e2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2e3 : romdata_int = 'h2b8;
    'h2e4 : romdata_int = 'h4a5;
    'h2e5 : romdata_int = 'h341c;
    'h2e6 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2e7 : romdata_int = 'h137;
    'h2e8 : romdata_int = 'h2687;
    'h2e9 : romdata_int = 'h5ab4;
    'h2ea : romdata_int = 'h278; // Line descriptor for 1_3
    'h2eb : romdata_int = 'h890;
    'h2ec : romdata_int = 'h1c78;
    'h2ed : romdata_int = 'h36ef;
    'h2ee : romdata_int = 'h278; // Line descriptor for 1_3
    'h2ef : romdata_int = 'h302;
    'h2f0 : romdata_int = 'h6665;
    'h2f1 : romdata_int = 'h72e1;
    'h2f2 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2f3 : romdata_int = 'h3032;
    'h2f4 : romdata_int = 'h3e0d;
    'h2f5 : romdata_int = 'h4c4f;
    'h2f6 : romdata_int = 'h278; // Line descriptor for 1_3
    'h2f7 : romdata_int = 'h16ee;
    'h2f8 : romdata_int = 'h1a2c;
    'h2f9 : romdata_int = 'h1a9a;
    'h2fa : romdata_int = 'h4278; // Line descriptor for 1_3
    'h2fb : romdata_int = 'h251e;
    'h2fc : romdata_int = 'h473e;
    'h2fd : romdata_int = 'h6f0b;
    'h2fe : romdata_int = 'h278; // Line descriptor for 1_3
    'h2ff : romdata_int = 'hc9f;
    'h300 : romdata_int = 'h22c8;
    'h301 : romdata_int = 'h6325;
    'h302 : romdata_int = 'h278; // Line descriptor for 1_3
    'h303 : romdata_int = 'h263d;
    'h304 : romdata_int = 'h12c0;
    'h305 : romdata_int = 'h1218;
    'h306 : romdata_int = 'h278; // Line descriptor for 1_3
    'h307 : romdata_int = 'h1835;
    'h308 : romdata_int = 'h1882;
    'h309 : romdata_int = 'h26d9;
    'h30a : romdata_int = 'h278; // Line descriptor for 1_3
    'h30b : romdata_int = 'h62df;
    'h30c : romdata_int = 'h2759;
    'h30d : romdata_int = 'h263a;
    'h30e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h30f : romdata_int = 'h467;
    'h310 : romdata_int = 'h6a7;
    'h311 : romdata_int = 'h12eb;
    'h312 : romdata_int = 'h278; // Line descriptor for 1_3
    'h313 : romdata_int = 'h5364;
    'h314 : romdata_int = 'h1ca6;
    'h315 : romdata_int = 'h395f;
    'h316 : romdata_int = 'h278; // Line descriptor for 1_3
    'h317 : romdata_int = 'he1a;
    'h318 : romdata_int = 'h12fd;
    'h319 : romdata_int = 'h5352;
    'h31a : romdata_int = 'h278; // Line descriptor for 1_3
    'h31b : romdata_int = 'h8;
    'h31c : romdata_int = 'h1ca8;
    'h31d : romdata_int = 'h4854;
    'h31e : romdata_int = 'h278; // Line descriptor for 1_3
    'h31f : romdata_int = 'h27f;
    'h320 : romdata_int = 'h3419;
    'h321 : romdata_int = 'h3cbd;
    'h322 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h323 : romdata_int = 'h147f;
    'h324 : romdata_int = 'h210b;
    'h325 : romdata_int = 'h3352;
    'h326 : romdata_int = 'h278; // Line descriptor for 1_3
    'h327 : romdata_int = 'hb27;
    'h328 : romdata_int = 'h1033;
    'h329 : romdata_int = 'h3e79;
    'h32a : romdata_int = 'h278; // Line descriptor for 1_3
    'h32b : romdata_int = 'h1b31;
    'h32c : romdata_int = 'hc70;
    'h32d : romdata_int = 'h8b6;
    'h32e : romdata_int = 'h278; // Line descriptor for 1_3
    'h32f : romdata_int = 'h4f4e;
    'h330 : romdata_int = 'h5e05;
    'h331 : romdata_int = 'h1a0a;
    'h332 : romdata_int = 'h278; // Line descriptor for 1_3
    'h333 : romdata_int = 'hc75;
    'h334 : romdata_int = 'h1208;
    'h335 : romdata_int = 'h550b;
    'h336 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h337 : romdata_int = 'h1050;
    'h338 : romdata_int = 'h1ac4;
    'h339 : romdata_int = 'h424f;
    'h33a : romdata_int = 'h278; // Line descriptor for 1_3
    'h33b : romdata_int = 'h67c;
    'h33c : romdata_int = 'h6a4;
    'h33d : romdata_int = 'hd38;
    'h33e : romdata_int = 'h278; // Line descriptor for 1_3
    'h33f : romdata_int = 'h3955;
    'h340 : romdata_int = 'h4134;
    'h341 : romdata_int = 'h5a38;
    'h342 : romdata_int = 'h278; // Line descriptor for 1_3
    'h343 : romdata_int = 'hc82;
    'h344 : romdata_int = 'h553d;
    'h345 : romdata_int = 'h6ef4;
    'h346 : romdata_int = 'h278; // Line descriptor for 1_3
    'h347 : romdata_int = 'h122;
    'h348 : romdata_int = 'h2126;
    'h349 : romdata_int = 'h50b3;
    'h34a : romdata_int = 'h4278; // Line descriptor for 1_3
    'h34b : romdata_int = 'h29b;
    'h34c : romdata_int = 'h105f;
    'h34d : romdata_int = 'h7015;
    'h34e : romdata_int = 'h278; // Line descriptor for 1_3
    'h34f : romdata_int = 'h125d;
    'h350 : romdata_int = 'h40d;
    'h351 : romdata_int = 'h27c;
    'h352 : romdata_int = 'h278; // Line descriptor for 1_3
    'h353 : romdata_int = 'h1873;
    'h354 : romdata_int = 'h2698;
    'h355 : romdata_int = 'h6944;
    'h356 : romdata_int = 'h278; // Line descriptor for 1_3
    'h357 : romdata_int = 'h127b;
    'h358 : romdata_int = 'h575c;
    'h359 : romdata_int = 'h1867;
    'h35a : romdata_int = 'h278; // Line descriptor for 1_3
    'h35b : romdata_int = 'h294c;
    'h35c : romdata_int = 'h5f25;
    'h35d : romdata_int = 'h74d9;
    'h35e : romdata_int = 'h4278; // Line descriptor for 1_3
    'h35f : romdata_int = 'h6a6;
    'h360 : romdata_int = 'h1ac9;
    'h361 : romdata_int = 'h2360;
    'h362 : romdata_int = 'h278; // Line descriptor for 1_3
    'h363 : romdata_int = 'heee;
    'h364 : romdata_int = 'h1e6b;
    'h365 : romdata_int = 'h6245;
    'h366 : romdata_int = 'h278; // Line descriptor for 1_3
    'h367 : romdata_int = 'h1d4b;
    'h368 : romdata_int = 'h2262;
    'h369 : romdata_int = 'h446b;
    'h36a : romdata_int = 'h278; // Line descriptor for 1_3
    'h36b : romdata_int = 'h8f2;
    'h36c : romdata_int = 'h271c;
    'h36d : romdata_int = 'h2721;
    'h36e : romdata_int = 'h278; // Line descriptor for 1_3
    'h36f : romdata_int = 'h2b44;
    'h370 : romdata_int = 'h3e81;
    'h371 : romdata_int = 'h214c;
    'h372 : romdata_int = 'h4278; // Line descriptor for 1_3
    'h373 : romdata_int = 'h1b5b;
    'h374 : romdata_int = 'h5038;
    'h375 : romdata_int = 'h2a76;
    'h376 : romdata_int = 'h278; // Line descriptor for 1_3
    'h377 : romdata_int = 'h18c5;
    'h378 : romdata_int = 'h3d5b;
    'h379 : romdata_int = 'h6629;
    'h37a : romdata_int = 'h278; // Line descriptor for 1_3
    'h37b : romdata_int = 'h260;
    'h37c : romdata_int = 'ha48;
    'h37d : romdata_int = 'he0a;
    'h37e : romdata_int = 'h278; // Line descriptor for 1_3
    'h37f : romdata_int = 'h643;
    'h380 : romdata_int = 'h6b0;
    'h381 : romdata_int = 'h5506;
    'h382 : romdata_int = 'h278; // Line descriptor for 1_3
    'h383 : romdata_int = 'h238;
    'h384 : romdata_int = 'he32;
    'h385 : romdata_int = 'h10a2;
    'h386 : romdata_int = 'h6278; // Line descriptor for 1_3
    'h387 : romdata_int = 'h528;
    'h388 : romdata_int = 'h1cf5;
    'h389 : romdata_int = 'h492f;
    'h38a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h38b : romdata_int = 'h2e;
    'h38c : romdata_int = 'hb0;
    'h38d : romdata_int = 'h4107;
    'h38e : romdata_int = 'h8f1c;
    'h38f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h390 : romdata_int = 'h22f3;
    'h391 : romdata_int = 'h2680;
    'h392 : romdata_int = 'h2ead;
    'h393 : romdata_int = 'h5a42;
    'h394 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h395 : romdata_int = 'hd38;
    'h396 : romdata_int = 'h1763;
    'h397 : romdata_int = 'h38d6;
    'h398 : romdata_int = 'h5089;
    'h399 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h39a : romdata_int = 'h27f;
    'h39b : romdata_int = 'h1937;
    'h39c : romdata_int = 'h2ed5;
    'h39d : romdata_int = 'h632a;
    'h39e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h39f : romdata_int = 'habd;
    'h3a0 : romdata_int = 'h1b4c;
    'h3a1 : romdata_int = 'h2107;
    'h3a2 : romdata_int = 'h8e89;
    'h3a3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3a4 : romdata_int = 'h8c9;
    'h3a5 : romdata_int = 'ha67;
    'h3a6 : romdata_int = 'h1c14;
    'h3a7 : romdata_int = 'h853a;
    'h3a8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3a9 : romdata_int = 'h14e5;
    'h3aa : romdata_int = 'h2236;
    'h3ab : romdata_int = 'h22f9;
    'h3ac : romdata_int = 'h5896;
    'h3ad : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3ae : romdata_int = 'h1338;
    'h3af : romdata_int = 'h30a0;
    'h3b0 : romdata_int = 'h403d;
    'h3b1 : romdata_int = 'h7b3d;
    'h3b2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3b3 : romdata_int = 'h10df;
    'h3b4 : romdata_int = 'h1887;
    'h3b5 : romdata_int = 'h28b1;
    'h3b6 : romdata_int = 'h5c58;
    'h3b7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3b8 : romdata_int = 'h461;
    'h3b9 : romdata_int = 'h1408;
    'h3ba : romdata_int = 'h26db;
    'h3bb : romdata_int = 'h5718;
    'h3bc : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3bd : romdata_int = 'h1690;
    'h3be : romdata_int = 'h24e2;
    'h3bf : romdata_int = 'h2ae6;
    'h3c0 : romdata_int = 'h8663;
    'h3c1 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3c2 : romdata_int = 'h183e;
    'h3c3 : romdata_int = 'h1ea6;
    'h3c4 : romdata_int = 'h226c;
    'h3c5 : romdata_int = 'h54a0;
    'h3c6 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3c7 : romdata_int = 'h86;
    'h3c8 : romdata_int = 'h4e0;
    'h3c9 : romdata_int = 'h2a26;
    'h3ca : romdata_int = 'h5ccb;
    'h3cb : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3cc : romdata_int = 'hf48;
    'h3cd : romdata_int = 'h89;
    'h3ce : romdata_int = 'h78cd;
    'h3cf : romdata_int = 'h1135;
    'h3d0 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3d1 : romdata_int = 'h1ced;
    'h3d2 : romdata_int = 'h3735;
    'h3d3 : romdata_int = 'h3521;
    'h3d4 : romdata_int = 'h5ed9;
    'h3d5 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3d6 : romdata_int = 'h727a;
    'h3d7 : romdata_int = 'h1ccb;
    'h3d8 : romdata_int = 'h2d08;
    'h3d9 : romdata_int = 'h2f62;
    'h3da : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3db : romdata_int = 'h1ef5;
    'h3dc : romdata_int = 'h22ee;
    'h3dd : romdata_int = 'h7661;
    'h3de : romdata_int = 'h2aba;
    'h3df : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3e0 : romdata_int = 'h877;
    'h3e1 : romdata_int = 'h1144;
    'h3e2 : romdata_int = 'h2ee4;
    'h3e3 : romdata_int = 'h760b;
    'h3e4 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3e5 : romdata_int = 'hea1;
    'h3e6 : romdata_int = 'h12ce;
    'h3e7 : romdata_int = 'h2a70;
    'h3e8 : romdata_int = 'h7ec4;
    'h3e9 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3ea : romdata_int = 'hd4f;
    'h3eb : romdata_int = 'h10d6;
    'h3ec : romdata_int = 'h1746;
    'h3ed : romdata_int = 'h887a;
    'h3ee : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3ef : romdata_int = 'h33b;
    'h3f0 : romdata_int = 'haa6;
    'h3f1 : romdata_int = 'h1b15;
    'h3f2 : romdata_int = 'h760e;
    'h3f3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3f4 : romdata_int = 'hf2a;
    'h3f5 : romdata_int = 'h1d1f;
    'h3f6 : romdata_int = 'h2c0d;
    'h3f7 : romdata_int = 'h60ad;
    'h3f8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h3f9 : romdata_int = 'h46b;
    'h3fa : romdata_int = 'h18c3;
    'h3fb : romdata_int = 'h2034;
    'h3fc : romdata_int = 'h7046;
    'h3fd : romdata_int = 'h436c; // Line descriptor for 2_5
    'h3fe : romdata_int = 'h4;
    'h3ff : romdata_int = 'h12fe;
    'h400 : romdata_int = 'h145d;
    'h401 : romdata_int = 'h82b8;
    'h402 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h403 : romdata_int = 'h642;
    'h404 : romdata_int = 'h84a;
    'h405 : romdata_int = 'haf2;
    'h406 : romdata_int = 'h62fe;
    'h407 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h408 : romdata_int = 'h209e;
    'h409 : romdata_int = 'h267e;
    'h40a : romdata_int = 'h30b0;
    'h40b : romdata_int = 'h7062;
    'h40c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h40d : romdata_int = 'h8d5;
    'h40e : romdata_int = 'h108d;
    'h40f : romdata_int = 'h2667;
    'h410 : romdata_int = 'h6b09;
    'h411 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h412 : romdata_int = 'h312;
    'h413 : romdata_int = 'h2039;
    'h414 : romdata_int = 'h2d1d;
    'h415 : romdata_int = 'h4eea;
    'h416 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h417 : romdata_int = 'hd4d;
    'h418 : romdata_int = 'h10a0;
    'h419 : romdata_int = 'h444b;
    'h41a : romdata_int = 'h6517;
    'h41b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h41c : romdata_int = 'h299;
    'h41d : romdata_int = 'h92b;
    'h41e : romdata_int = 'h2e18;
    'h41f : romdata_int = 'h8149;
    'h420 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h421 : romdata_int = 'hcab;
    'h422 : romdata_int = 'h6703;
    'h423 : romdata_int = 'h6b0;
    'h424 : romdata_int = 'h2549;
    'h425 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h426 : romdata_int = 'h3762;
    'h427 : romdata_int = 'hc8f;
    'h428 : romdata_int = 'h6ab6;
    'h429 : romdata_int = 'h16b4;
    'h42a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h42b : romdata_int = 'h1221;
    'h42c : romdata_int = 'h1e3f;
    'h42d : romdata_int = 'h2467;
    'h42e : romdata_int = 'h4c86;
    'h42f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h430 : romdata_int = 'h3ed1;
    'h431 : romdata_int = 'h8b20;
    'h432 : romdata_int = 'h12fd;
    'h433 : romdata_int = 'h2291;
    'h434 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h435 : romdata_int = 'h9a;
    'h436 : romdata_int = 'h14c0;
    'h437 : romdata_int = 'h1f38;
    'h438 : romdata_int = 'h72f8;
    'h439 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h43a : romdata_int = 'hc70;
    'h43b : romdata_int = 'h1a64;
    'h43c : romdata_int = 'h2ae3;
    'h43d : romdata_int = 'h8706;
    'h43e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h43f : romdata_int = 'h121c;
    'h440 : romdata_int = 'h1f4b;
    'h441 : romdata_int = 'h2257;
    'h442 : romdata_int = 'h6109;
    'h443 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h444 : romdata_int = 'h455;
    'h445 : romdata_int = 'h167e;
    'h446 : romdata_int = 'h430f;
    'h447 : romdata_int = 'h826b;
    'h448 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h449 : romdata_int = 'h109b;
    'h44a : romdata_int = 'h1b58;
    'h44b : romdata_int = 'h18ca;
    'h44c : romdata_int = 'h7c7b;
    'h44d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h44e : romdata_int = 'h864;
    'h44f : romdata_int = 'h168f;
    'h450 : romdata_int = 'h1aad;
    'h451 : romdata_int = 'h4a4e;
    'h452 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h453 : romdata_int = 'he66;
    'h454 : romdata_int = 'h208b;
    'h455 : romdata_int = 'h6525;
    'h456 : romdata_int = 'h2c79;
    'h457 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h458 : romdata_int = 'h936;
    'h459 : romdata_int = 'ha88;
    'h45a : romdata_int = 'h26b5;
    'h45b : romdata_int = 'h6505;
    'h45c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h45d : romdata_int = 'h2469;
    'h45e : romdata_int = 'hae;
    'h45f : romdata_int = 'h1b06;
    'h460 : romdata_int = 'h7553;
    'h461 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h462 : romdata_int = 'h1670;
    'h463 : romdata_int = 'h24ff;
    'h464 : romdata_int = 'h3326;
    'h465 : romdata_int = 'h88ca;
    'h466 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h467 : romdata_int = 'hf16;
    'h468 : romdata_int = 'h1ea1;
    'h469 : romdata_int = 'h2166;
    'h46a : romdata_int = 'h8a28;
    'h46b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h46c : romdata_int = 'h4e6;
    'h46d : romdata_int = 'h161f;
    'h46e : romdata_int = 'h1a17;
    'h46f : romdata_int = 'h4af0;
    'h470 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h471 : romdata_int = 'hd5;
    'h472 : romdata_int = 'h2f3e;
    'h473 : romdata_int = 'h4009;
    'h474 : romdata_int = 'h7493;
    'h475 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h476 : romdata_int = 'hc41;
    'h477 : romdata_int = 'h1d3d;
    'h478 : romdata_int = 'h2630;
    'h479 : romdata_int = 'h88c3;
    'h47a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h47b : romdata_int = 'h10b;
    'h47c : romdata_int = 'h51e;
    'h47d : romdata_int = 'h2b59;
    'h47e : romdata_int = 'h5248;
    'h47f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h480 : romdata_int = 'h643;
    'h481 : romdata_int = 'h173f;
    'h482 : romdata_int = 'h293b;
    'h483 : romdata_int = 'h4a7b;
    'h484 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h485 : romdata_int = 'h2e54;
    'h486 : romdata_int = 'h6a7;
    'h487 : romdata_int = 'h687b;
    'h488 : romdata_int = 'h27c;
    'h489 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h48a : romdata_int = 'h44bb;
    'h48b : romdata_int = 'h5813;
    'h48c : romdata_int = 'h1a2b;
    'h48d : romdata_int = 'h6c9;
    'h48e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h48f : romdata_int = 'h1319;
    'h490 : romdata_int = 'h1958;
    'h491 : romdata_int = 'h36e6;
    'h492 : romdata_int = 'h8a2c;
    'h493 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h494 : romdata_int = 'h22f4;
    'h495 : romdata_int = 'h2441;
    'h496 : romdata_int = 'h2c81;
    'h497 : romdata_int = 'h7d47;
    'h498 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h499 : romdata_int = 'hc0e;
    'h49a : romdata_int = 'h122a;
    'h49b : romdata_int = 'h1a42;
    'h49c : romdata_int = 'h4cb6;
    'h49d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h49e : romdata_int = 'h10d0;
    'h49f : romdata_int = 'h255e;
    'h4a0 : romdata_int = 'h26a8;
    'h4a1 : romdata_int = 'h7260;
    'h4a2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4a3 : romdata_int = 'he4d;
    'h4a4 : romdata_int = 'h1030;
    'h4a5 : romdata_int = 'h3270;
    'h4a6 : romdata_int = 'h6874;
    'h4a7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4a8 : romdata_int = 'h18db;
    'h4a9 : romdata_int = 'h2145;
    'h4aa : romdata_int = 'h2d4c;
    'h4ab : romdata_int = 'h80a1;
    'h4ac : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4ad : romdata_int = 'h48a;
    'h4ae : romdata_int = 'h4d5;
    'h4af : romdata_int = 'h1522;
    'h4b0 : romdata_int = 'h5f38;
    'h4b1 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4b2 : romdata_int = 'h12c9;
    'h4b3 : romdata_int = 'h1845;
    'h4b4 : romdata_int = 'h46f7;
    'h4b5 : romdata_int = 'h664e;
    'h4b6 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4b7 : romdata_int = 'h1623;
    'h4b8 : romdata_int = 'hb22;
    'h4b9 : romdata_int = 'h520b;
    'h4ba : romdata_int = 'h42b8;
    'h4bb : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4bc : romdata_int = 'h5d67;
    'h4bd : romdata_int = 'h28d4;
    'h4be : romdata_int = 'h168c;
    'h4bf : romdata_int = 'h1d1d;
    'h4c0 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4c1 : romdata_int = 'h862;
    'h4c2 : romdata_int = 'hc25;
    'h4c3 : romdata_int = 'h2ec7;
    'h4c4 : romdata_int = 'h50ec;
    'h4c5 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4c6 : romdata_int = 'h253f;
    'h4c7 : romdata_int = 'h266e;
    'h4c8 : romdata_int = 'h2d61;
    'h4c9 : romdata_int = 'h8537;
    'h4ca : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4cb : romdata_int = 'ha5c;
    'h4cc : romdata_int = 'h5ab5;
    'h4cd : romdata_int = 'h954;
    'h4ce : romdata_int = 'h2645;
    'h4cf : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4d0 : romdata_int = 'h668d;
    'h4d1 : romdata_int = 'h214d;
    'h4d2 : romdata_int = 'hb49;
    'h4d3 : romdata_int = 'h3b4f;
    'h4d4 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4d5 : romdata_int = 'h673;
    'h4d6 : romdata_int = 'h187b;
    'h4d7 : romdata_int = 'h2081;
    'h4d8 : romdata_int = 'h74c6;
    'h4d9 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4da : romdata_int = 'h2b8;
    'h4db : romdata_int = 'h10be;
    'h4dc : romdata_int = 'h3c01;
    'h4dd : romdata_int = 'h4913;
    'h4de : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4df : romdata_int = 'h890;
    'h4e0 : romdata_int = 'h2151;
    'h4e1 : romdata_int = 'h4220;
    'h4e2 : romdata_int = 'h551d;
    'h4e3 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4e4 : romdata_int = 'hef3;
    'h4e5 : romdata_int = 'h2665;
    'h4e6 : romdata_int = 'h4750;
    'h4e7 : romdata_int = 'h62d2;
    'h4e8 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4e9 : romdata_int = 'h27b;
    'h4ea : romdata_int = 'h1006;
    'h4eb : romdata_int = 'h2749;
    'h4ec : romdata_int = 'h5431;
    'h4ed : romdata_int = 'h436c; // Line descriptor for 2_5
    'h4ee : romdata_int = 'h137;
    'h4ef : romdata_int = 'h16da;
    'h4f0 : romdata_int = 'h2e36;
    'h4f1 : romdata_int = 'h6c29;
    'h4f2 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4f3 : romdata_int = 'h4a5;
    'h4f4 : romdata_int = 'h24a4;
    'h4f5 : romdata_int = 'h2aed;
    'h4f6 : romdata_int = 'h6e6e;
    'h4f7 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4f8 : romdata_int = 'h29b;
    'h4f9 : romdata_int = 'h1031;
    'h4fa : romdata_int = 'h28f3;
    'h4fb : romdata_int = 'h56fa;
    'h4fc : romdata_int = 'h36c; // Line descriptor for 2_5
    'h4fd : romdata_int = 'h185c;
    'h4fe : romdata_int = 'h18ee;
    'h4ff : romdata_int = 'h3e87;
    'h500 : romdata_int = 'h6a17;
    'h501 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h502 : romdata_int = 'h2449;
    'h503 : romdata_int = 'h3a61;
    'h504 : romdata_int = 'h3c42;
    'h505 : romdata_int = 'h60a7;
    'h506 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h507 : romdata_int = 'h6e5;
    'h508 : romdata_int = 'h1efc;
    'h509 : romdata_int = 'h30fc;
    'h50a : romdata_int = 'h4d54;
    'h50b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h50c : romdata_int = 'h2a85;
    'h50d : romdata_int = 'h2d2c;
    'h50e : romdata_int = 'h8c33;
    'h50f : romdata_int = 'h3f61;
    'h510 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h511 : romdata_int = 'h143f;
    'h512 : romdata_int = 'h1a35;
    'h513 : romdata_int = 'h1c9a;
    'h514 : romdata_int = 'h8c2c;
    'h515 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h516 : romdata_int = 'h6a6;
    'h517 : romdata_int = 'h1906;
    'h518 : romdata_int = 'h255d;
    'h519 : romdata_int = 'h8e9c;
    'h51a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h51b : romdata_int = 'h467;
    'h51c : romdata_int = 'he1a;
    'h51d : romdata_int = 'hf58;
    'h51e : romdata_int = 'h7a2f;
    'h51f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h520 : romdata_int = 'h1418;
    'h521 : romdata_int = 'h271e;
    'h522 : romdata_int = 'h2c4f;
    'h523 : romdata_int = 'h7e0d;
    'h524 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h525 : romdata_int = 'h283d;
    'h526 : romdata_int = 'h28d9;
    'h527 : romdata_int = 'h2f2f;
    'h528 : romdata_int = 'h4e43;
    'h529 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h52a : romdata_int = 'h8;
    'h52b : romdata_int = 'hb27;
    'h52c : romdata_int = 'h14eb;
    'h52d : romdata_int = 'h86b9;
    'h52e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h52f : romdata_int = 'h238;
    'h530 : romdata_int = 'h283a;
    'h531 : romdata_int = 'h2959;
    'h532 : romdata_int = 'h6889;
    'h533 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h534 : romdata_int = 'h14fd;
    'h535 : romdata_int = 'hc82;
    'h536 : romdata_int = 'h24c8;
    'h537 : romdata_int = 'h8332;
    'h538 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h539 : romdata_int = 'h7951;
    'h53a : romdata_int = 'h1440;
    'h53b : romdata_int = 'h1e97;
    'h53c : romdata_int = 'h1d31;
    'h53d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h53e : romdata_int = 'h230b;
    'h53f : romdata_int = 'h28ba;
    'h540 : romdata_int = 'h395f;
    'h541 : romdata_int = 'h8448;
    'h542 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h543 : romdata_int = 'h8b6;
    'h544 : romdata_int = 'h1233;
    'h545 : romdata_int = 'h3470;
    'h546 : romdata_int = 'h487d;
    'h547 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h548 : romdata_int = 'hc75;
    'h549 : romdata_int = 'h1465;
    'h54a : romdata_int = 'h6e4d;
    'h54b : romdata_int = 'h2efc;
    'h54c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h54d : romdata_int = 'h72c;
    'h54e : romdata_int = 'hd52;
    'h54f : romdata_int = 'h1ed5;
    'h550 : romdata_int = 'h6f06;
    'h551 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h552 : romdata_int = 'h3d47;
    'h553 : romdata_int = 'h4845;
    'h554 : romdata_int = 'h67c;
    'h555 : romdata_int = 'h1cc4;
    'h556 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h557 : romdata_int = 'hb34;
    'h558 : romdata_int = 'h1250;
    'h559 : romdata_int = 'h32ee;
    'h55a : romdata_int = 'h6cf3;
    'h55b : romdata_int = 'h36c; // Line descriptor for 2_5
    'h55c : romdata_int = 'h122;
    'h55d : romdata_int = 'h2099;
    'h55e : romdata_int = 'h2cc6;
    'h55f : romdata_int = 'h8c12;
    'h560 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h561 : romdata_int = 'h302;
    'h562 : romdata_int = 'h1a73;
    'h563 : romdata_int = 'h2898;
    'h564 : romdata_int = 'h5b28;
    'h565 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h566 : romdata_int = 'h40d;
    'h567 : romdata_int = 'h147b;
    'h568 : romdata_int = 'h1c0a;
    'h569 : romdata_int = 'h791a;
    'h56a : romdata_int = 'h36c; // Line descriptor for 2_5
    'h56b : romdata_int = 'h2ef5;
    'h56c : romdata_int = 'h3544;
    'h56d : romdata_int = 'h3913;
    'h56e : romdata_int = 'h570b;
    'h56f : romdata_int = 'h36c; // Line descriptor for 2_5
    'h570 : romdata_int = 'h62d;
    'h571 : romdata_int = 'h2851;
    'h572 : romdata_int = 'h2ac2;
    'h573 : romdata_int = 'h7008;
    'h574 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h575 : romdata_int = 'heee;
    'h576 : romdata_int = 'h224a;
    'h577 : romdata_int = 'h46a6;
    'h578 : romdata_int = 'h7a68;
    'h579 : romdata_int = 'h436c; // Line descriptor for 2_5
    'h57a : romdata_int = 'h1cc9;
    'h57b : romdata_int = 'h206b;
    'h57c : romdata_int = 'h2326;
    'h57d : romdata_int = 'h5144;
    'h57e : romdata_int = 'h36c; // Line descriptor for 2_5
    'h57f : romdata_int = 'h1eb1;
    'h580 : romdata_int = 'h8f2;
    'h581 : romdata_int = 'h3b3d;
    'h582 : romdata_int = 'h4e29;
    'h583 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h584 : romdata_int = 'h2b43;
    'h585 : romdata_int = 'h2356;
    'h586 : romdata_int = 'h5f4b;
    'h587 : romdata_int = 'h1ea8;
    'h588 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h589 : romdata_int = 'hb01;
    'h58a : romdata_int = 'h1d5b;
    'h58b : romdata_int = 'h291c;
    'h58c : romdata_int = 'h5878;
    'h58d : romdata_int = 'h436c; // Line descriptor for 2_5
    'h58e : romdata_int = 'h1ac5;
    'h58f : romdata_int = 'h2a1b;
    'h590 : romdata_int = 'h2ae4;
    'h591 : romdata_int = 'h6c39;
    'h592 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h593 : romdata_int = 'h2d34;
    'h594 : romdata_int = 'h279;
    'h595 : romdata_int = 'he0a;
    'h596 : romdata_int = 'h7d08;
    'h597 : romdata_int = 'h36c; // Line descriptor for 2_5
    'h598 : romdata_int = 'h728;
    'h599 : romdata_int = 'h2cf2;
    'h59a : romdata_int = 'h4525;
    'h59b : romdata_int = 'h80d9;
    'h59c : romdata_int = 'h36c; // Line descriptor for 2_5
    'h59d : romdata_int = 'h2b9;
    'h59e : romdata_int = 'ha48;
    'h59f : romdata_int = 'h12a2;
    'h5a0 : romdata_int = 'h7e52;
    'h5a1 : romdata_int = 'h636c; // Line descriptor for 2_5
    'h5a2 : romdata_int = 'h528;
    'h5a3 : romdata_int = 'he32;
    'h5a4 : romdata_int = 'h1efe;
    'h5a5 : romdata_int = 'h5201;
    'h5a6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5a7 : romdata_int = 'h352c;
    'h5a8 : romdata_int = 'h3703;
    'h5a9 : romdata_int = 'h3c43;
    'h5aa : romdata_int = 'h4800;
    'h5ab : romdata_int = 'h94b5;
    'h5ac : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5ad : romdata_int = 'h1432;
    'h5ae : romdata_int = 'h143d;
    'h5af : romdata_int = 'h291e;
    'h5b0 : romdata_int = 'h4a00;
    'h5b1 : romdata_int = 'h529a;
    'h5b2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5b3 : romdata_int = 'h81f;
    'h5b4 : romdata_int = 'h200e;
    'h5b5 : romdata_int = 'h373e;
    'h5b6 : romdata_int = 'h4c00;
    'h5b7 : romdata_int = 'h668a;
    'h5b8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5b9 : romdata_int = 'h506;
    'h5ba : romdata_int = 'hc45;
    'h5bb : romdata_int = 'h210b;
    'h5bc : romdata_int = 'h4e00;
    'h5bd : romdata_int = 'h8960;
    'h5be : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5bf : romdata_int = 'h133d;
    'h5c0 : romdata_int = 'h30ef;
    'h5c1 : romdata_int = 'h4224;
    'h5c2 : romdata_int = 'h5000;
    'h5c3 : romdata_int = 'ha516;
    'h5c4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5c5 : romdata_int = 'h698;
    'h5c6 : romdata_int = 'h1afe;
    'h5c7 : romdata_int = 'h3088;
    'h5c8 : romdata_int = 'h3cd1;
    'h5c9 : romdata_int = 'h5200;
    'h5ca : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5cb : romdata_int = 'h1d1e;
    'h5cc : romdata_int = 'h2a67;
    'h5cd : romdata_int = 'h40ec;
    'h5ce : romdata_int = 'h5400;
    'h5cf : romdata_int = 'h9952;
    'h5d0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5d1 : romdata_int = 'h87e;
    'h5d2 : romdata_int = 'h382c;
    'h5d3 : romdata_int = 'h4509;
    'h5d4 : romdata_int = 'h5600;
    'h5d5 : romdata_int = 'hb2d6;
    'h5d6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5d7 : romdata_int = 'h214c;
    'h5d8 : romdata_int = 'h240f;
    'h5d9 : romdata_int = 'h3d29;
    'h5da : romdata_int = 'h5800;
    'h5db : romdata_int = 'hae31;
    'h5dc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5dd : romdata_int = 'h2b55;
    'h5de : romdata_int = 'h3155;
    'h5df : romdata_int = 'h5a00;
    'h5e0 : romdata_int = 'h7528;
    'h5e1 : romdata_int = 'h9f61;
    'h5e2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5e3 : romdata_int = 'h21c;
    'h5e4 : romdata_int = 'h88c;
    'h5e5 : romdata_int = 'hab0;
    'h5e6 : romdata_int = 'h4a01;
    'h5e7 : romdata_int = 'h5c00;
    'h5e8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5e9 : romdata_int = 'h1115;
    'h5ea : romdata_int = 'h26c8;
    'h5eb : romdata_int = 'h2885;
    'h5ec : romdata_int = 'h40aa;
    'h5ed : romdata_int = 'h5e00;
    'h5ee : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5ef : romdata_int = 'h1f4d;
    'h5f0 : romdata_int = 'h344f;
    'h5f1 : romdata_int = 'h42b5;
    'h5f2 : romdata_int = 'h6000;
    'h5f3 : romdata_int = 'h9cc5;
    'h5f4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5f5 : romdata_int = 'h1064;
    'h5f6 : romdata_int = 'h2091;
    'h5f7 : romdata_int = 'h5d3b;
    'h5f8 : romdata_int = 'h6200;
    'h5f9 : romdata_int = 'h84e7;
    'h5fa : romdata_int = 'h45a; // Line descriptor for 1_2
    'h5fb : romdata_int = 'h1c;
    'h5fc : romdata_int = 'h24e2;
    'h5fd : romdata_int = 'h6400;
    'h5fe : romdata_int = 'h7e64;
    'h5ff : romdata_int = 'h8683;
    'h600 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h601 : romdata_int = 'h1aa6;
    'h602 : romdata_int = 'h2f4f;
    'h603 : romdata_int = 'h3cb8;
    'h604 : romdata_int = 'h6600;
    'h605 : romdata_int = 'h7f2b;
    'h606 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h607 : romdata_int = 'hc87;
    'h608 : romdata_int = 'h16ef;
    'h609 : romdata_int = 'h6800;
    'h60a : romdata_int = 'h767c;
    'h60b : romdata_int = 'h9255;
    'h60c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h60d : romdata_int = 'h10ad;
    'h60e : romdata_int = 'h3636;
    'h60f : romdata_int = 'h6279;
    'h610 : romdata_int = 'h6a00;
    'h611 : romdata_int = 'h712e;
    'h612 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h613 : romdata_int = 'h1c6e;
    'h614 : romdata_int = 'h2e33;
    'h615 : romdata_int = 'h3311;
    'h616 : romdata_int = 'h6c00;
    'h617 : romdata_int = 'ha2a1;
    'h618 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h619 : romdata_int = 'h4c0;
    'h61a : romdata_int = 'h1e8b;
    'h61b : romdata_int = 'h38a0;
    'h61c : romdata_int = 'h4c72;
    'h61d : romdata_int = 'h6e00;
    'h61e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h61f : romdata_int = 'h1632;
    'h620 : romdata_int = 'h2622;
    'h621 : romdata_int = 'h3f25;
    'h622 : romdata_int = 'h7000;
    'h623 : romdata_int = 'h945e;
    'h624 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h625 : romdata_int = 'h132;
    'h626 : romdata_int = 'h1017;
    'h627 : romdata_int = 'h16bc;
    'h628 : romdata_int = 'h7200;
    'h629 : romdata_int = 'h8718;
    'h62a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h62b : romdata_int = 'h2659;
    'h62c : romdata_int = 'h3f32;
    'h62d : romdata_int = 'h7400;
    'h62e : romdata_int = 'h8f22;
    'h62f : romdata_int = 'haa37;
    'h630 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h631 : romdata_int = 'h6cf;
    'h632 : romdata_int = 'h122c;
    'h633 : romdata_int = 'h26aa;
    'h634 : romdata_int = 'h5ab8;
    'h635 : romdata_int = 'h7600;
    'h636 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h637 : romdata_int = 'h823;
    'h638 : romdata_int = 'h2249;
    'h639 : romdata_int = 'h46cc;
    'h63a : romdata_int = 'h6861;
    'h63b : romdata_int = 'h7800;
    'h63c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h63d : romdata_int = 'h2603;
    'h63e : romdata_int = 'h3121;
    'h63f : romdata_int = 'h36e4;
    'h640 : romdata_int = 'h7a00;
    'h641 : romdata_int = 'h9c4c;
    'h642 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h643 : romdata_int = 'h521;
    'h644 : romdata_int = 'h3a75;
    'h645 : romdata_int = 'h6855;
    'h646 : romdata_int = 'h7c00;
    'h647 : romdata_int = 'ha6f3;
    'h648 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h649 : romdata_int = 'he82;
    'h64a : romdata_int = 'h1aa8;
    'h64b : romdata_int = 'h4445;
    'h64c : romdata_int = 'h7e00;
    'h64d : romdata_int = 'h8413;
    'h64e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h64f : romdata_int = 'h2511;
    'h650 : romdata_int = 'h334c;
    'h651 : romdata_int = 'h400a;
    'h652 : romdata_int = 'h5a7b;
    'h653 : romdata_int = 'h8000;
    'h654 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h655 : romdata_int = 'haee;
    'h656 : romdata_int = 'hcee;
    'h657 : romdata_int = 'h1c4a;
    'h658 : romdata_int = 'h468d;
    'h659 : romdata_int = 'h8200;
    'h65a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h65b : romdata_int = 'h287e;
    'h65c : romdata_int = 'h2c3d;
    'h65d : romdata_int = 'h5e9b;
    'h65e : romdata_int = 'h8400;
    'h65f : romdata_int = 'hac1e;
    'h660 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h661 : romdata_int = 'h680;
    'h662 : romdata_int = 'h946;
    'h663 : romdata_int = 'h5cb9;
    'h664 : romdata_int = 'h8600;
    'h665 : romdata_int = 'ha0e9;
    'h666 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h667 : romdata_int = 'hcca;
    'h668 : romdata_int = 'h2349;
    'h669 : romdata_int = 'h32bd;
    'h66a : romdata_int = 'h80d5;
    'h66b : romdata_int = 'h8800;
    'h66c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h66d : romdata_int = 'h1e6f;
    'h66e : romdata_int = 'h2057;
    'h66f : romdata_int = 'h4725;
    'h670 : romdata_int = 'h502e;
    'h671 : romdata_int = 'h8a00;
    'h672 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h673 : romdata_int = 'h162f;
    'h674 : romdata_int = 'h1920;
    'h675 : romdata_int = 'h8c00;
    'h676 : romdata_int = 'h9aab;
    'h677 : romdata_int = 'hb144;
    'h678 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h679 : romdata_int = 'h1ce5;
    'h67a : romdata_int = 'h2c98;
    'h67b : romdata_int = 'h38ad;
    'h67c : romdata_int = 'h4915;
    'h67d : romdata_int = 'h8e00;
    'h67e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h67f : romdata_int = 'ha23;
    'h680 : romdata_int = 'h2ae5;
    'h681 : romdata_int = 'h3315;
    'h682 : romdata_int = 'h6728;
    'h683 : romdata_int = 'h9000;
    'h684 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h685 : romdata_int = 'h890;
    'h686 : romdata_int = 'h151d;
    'h687 : romdata_int = 'h3e45;
    'h688 : romdata_int = 'h7ac4;
    'h689 : romdata_int = 'h9200;
    'h68a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h68b : romdata_int = 'he67;
    'h68c : romdata_int = 'h14a4;
    'h68d : romdata_int = 'h4a2b;
    'h68e : romdata_int = 'h642a;
    'h68f : romdata_int = 'h9400;
    'h690 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h691 : romdata_int = 'h2865;
    'h692 : romdata_int = 'h354c;
    'h693 : romdata_int = 'h6165;
    'h694 : romdata_int = 'h9600;
    'h695 : romdata_int = 'h6e5f;
    'h696 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h697 : romdata_int = 'h1f51;
    'h698 : romdata_int = 'h2858;
    'h699 : romdata_int = 'h8c88;
    'h69a : romdata_int = 'h9670;
    'h69b : romdata_int = 'h9800;
    'h69c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h69d : romdata_int = 'h235d;
    'h69e : romdata_int = 'h3f13;
    'h69f : romdata_int = 'h72a7;
    'h6a0 : romdata_int = 'h7443;
    'h6a1 : romdata_int = 'h9a00;
    'h6a2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6a3 : romdata_int = 'h2137;
    'h6a4 : romdata_int = 'h28ee;
    'h6a5 : romdata_int = 'h36f5;
    'h6a6 : romdata_int = 'h9c00;
    'h6a7 : romdata_int = 'hac49;
    'h6a8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6a9 : romdata_int = 'h1c3c;
    'h6aa : romdata_int = 'h2a32;
    'h6ab : romdata_int = 'h7673;
    'h6ac : romdata_int = 'h9e00;
    'h6ad : romdata_int = 'hb2df;
    'h6ae : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6af : romdata_int = 'h103c;
    'h6b0 : romdata_int = 'h2694;
    'h6b1 : romdata_int = 'h326b;
    'h6b2 : romdata_int = 'h4e08;
    'h6b3 : romdata_int = 'ha000;
    'h6b4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6b5 : romdata_int = 'h233;
    'h6b6 : romdata_int = 'ha44;
    'h6b7 : romdata_int = 'h243a;
    'h6b8 : romdata_int = 'h2cb1;
    'h6b9 : romdata_int = 'ha200;
    'h6ba : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6bb : romdata_int = 'he41;
    'h6bc : romdata_int = 'h2b49;
    'h6bd : romdata_int = 'h4219;
    'h6be : romdata_int = 'h8e48;
    'h6bf : romdata_int = 'ha400;
    'h6c0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6c1 : romdata_int = 'h5f;
    'h6c2 : romdata_int = 'h34a5;
    'h6c3 : romdata_int = 'h64ef;
    'h6c4 : romdata_int = 'h8354;
    'h6c5 : romdata_int = 'ha600;
    'h6c6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6c7 : romdata_int = 'h67;
    'h6c8 : romdata_int = 'h14b3;
    'h6c9 : romdata_int = 'h1ccc;
    'h6ca : romdata_int = 'h46d3;
    'h6cb : romdata_int = 'ha800;
    'h6cc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6cd : romdata_int = 'h71;
    'h6ce : romdata_int = 'haba;
    'h6cf : romdata_int = 'h3a13;
    'h6d0 : romdata_int = 'h4328;
    'h6d1 : romdata_int = 'haa00;
    'h6d2 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6d3 : romdata_int = 'h338;
    'h6d4 : romdata_int = 'h16f8;
    'h6d5 : romdata_int = 'h1874;
    'h6d6 : romdata_int = 'h7894;
    'h6d7 : romdata_int = 'hac00;
    'h6d8 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6d9 : romdata_int = 'h228;
    'h6da : romdata_int = 'h640;
    'h6db : romdata_int = 'h2af3;
    'h6dc : romdata_int = 'hae00;
    'h6dd : romdata_int = 'haae5;
    'h6de : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6df : romdata_int = 'haeb;
    'h6e0 : romdata_int = 'h235e;
    'h6e1 : romdata_int = 'h932b;
    'h6e2 : romdata_int = 'hae8d;
    'h6e3 : romdata_int = 'hb000;
    'h6e4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6e5 : romdata_int = 'h14f6;
    'h6e6 : romdata_int = 'h2e91;
    'h6e7 : romdata_int = 'h5089;
    'h6e8 : romdata_int = 'h88c5;
    'h6e9 : romdata_int = 'hb200;
    'h6ea : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6eb : romdata_int = 'h0;
    'h6ec : romdata_int = 'h722;
    'h6ed : romdata_int = 'hc5c;
    'h6ee : romdata_int = 'h1106;
    'h6ef : romdata_int = 'ha632;
    'h6f0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6f1 : romdata_int = 'h200;
    'h6f2 : romdata_int = 'h335b;
    'h6f3 : romdata_int = 'h3c05;
    'h6f4 : romdata_int = 'h6aa5;
    'h6f5 : romdata_int = 'hb006;
    'h6f6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6f7 : romdata_int = 'h400;
    'h6f8 : romdata_int = 'hd58;
    'h6f9 : romdata_int = 'h38b0;
    'h6fa : romdata_int = 'h3c20;
    'h6fb : romdata_int = 'h540b;
    'h6fc : romdata_int = 'h45a; // Line descriptor for 1_2
    'h6fd : romdata_int = 'h600;
    'h6fe : romdata_int = 'h6ab;
    'h6ff : romdata_int = 'h186a;
    'h700 : romdata_int = 'h3534;
    'h701 : romdata_int = 'h786a;
    'h702 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h703 : romdata_int = 'h800;
    'h704 : romdata_int = 'h93f;
    'h705 : romdata_int = 'h3a38;
    'h706 : romdata_int = 'h2ecf;
    'h707 : romdata_int = 'h4717;
    'h708 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h709 : romdata_int = 'ha00;
    'h70a : romdata_int = 'h2269;
    'h70b : romdata_int = 'h3a70;
    'h70c : romdata_int = 'h5859;
    'h70d : romdata_int = 'h6cae;
    'h70e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h70f : romdata_int = 'hc00;
    'h710 : romdata_int = 'h1967;
    'h711 : romdata_int = 'h2b37;
    'h712 : romdata_int = 'h4c02;
    'h713 : romdata_int = 'h732c;
    'h714 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h715 : romdata_int = 'he00;
    'h716 : romdata_int = 'h1956;
    'h717 : romdata_int = 'h3edf;
    'h718 : romdata_int = 'h7a4e;
    'h719 : romdata_int = 'h8d27;
    'h71a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h71b : romdata_int = 'h1000;
    'h71c : romdata_int = 'h181e;
    'h71d : romdata_int = 'h1844;
    'h71e : romdata_int = 'h4662;
    'h71f : romdata_int = 'h82c9;
    'h720 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h721 : romdata_int = 'h221;
    'h722 : romdata_int = 'h250;
    'h723 : romdata_int = 'h1200;
    'h724 : romdata_int = 'h3b44;
    'h725 : romdata_int = 'h4484;
    'h726 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h727 : romdata_int = 'h6b4;
    'h728 : romdata_int = 'h1400;
    'h729 : romdata_int = 'h2447;
    'h72a : romdata_int = 'h2f44;
    'h72b : romdata_int = 'h42e1;
    'h72c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h72d : romdata_int = 'h1600;
    'h72e : romdata_int = 'h1ad5;
    'h72f : romdata_int = 'h2267;
    'h730 : romdata_int = 'h5f12;
    'h731 : romdata_int = 'h9122;
    'h732 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h733 : romdata_int = 'hefd;
    'h734 : romdata_int = 'h1800;
    'h735 : romdata_int = 'h1e34;
    'h736 : romdata_int = 'h315f;
    'h737 : romdata_int = 'ha24d;
    'h738 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h739 : romdata_int = 'h12f6;
    'h73a : romdata_int = 'h1a00;
    'h73b : romdata_int = 'h3d0f;
    'h73c : romdata_int = 'h44e8;
    'h73d : romdata_int = 'h621e;
    'h73e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h73f : romdata_int = 'hcc3;
    'h740 : romdata_int = 'h1c00;
    'h741 : romdata_int = 'h3ef7;
    'h742 : romdata_int = 'h40ce;
    'h743 : romdata_int = 'h563a;
    'h744 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h745 : romdata_int = 'h1e00;
    'h746 : romdata_int = 'h2d59;
    'h747 : romdata_int = 'h347e;
    'h748 : romdata_int = 'h9e8a;
    'h749 : romdata_int = 'ha858;
    'h74a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h74b : romdata_int = 'h308;
    'h74c : romdata_int = 'h1af5;
    'h74d : romdata_int = 'h2000;
    'h74e : romdata_int = 'h2810;
    'h74f : romdata_int = 'h4089;
    'h750 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h751 : romdata_int = 'h512;
    'h752 : romdata_int = 'h2200;
    'h753 : romdata_int = 'h22a4;
    'h754 : romdata_int = 'h311c;
    'h755 : romdata_int = 'h383e;
    'h756 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h757 : romdata_int = 'h2400;
    'h758 : romdata_int = 'h408;
    'h759 : romdata_int = 'h44ad;
    'h75a : romdata_int = 'h4f0b;
    'h75b : romdata_int = 'h6ae0;
    'h75c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h75d : romdata_int = 'h24b8;
    'h75e : romdata_int = 'h2600;
    'h75f : romdata_int = 'h374a;
    'h760 : romdata_int = 'h464e;
    'h761 : romdata_int = 'h7cd8;
    'h762 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h763 : romdata_int = 'h2d1c;
    'h764 : romdata_int = 'h1331;
    'h765 : romdata_int = 'h12bb;
    'h766 : romdata_int = 'h2800;
    'h767 : romdata_int = 'h9682;
    'h768 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h769 : romdata_int = 'h2a00;
    'h76a : romdata_int = 'h2cd9;
    'h76b : romdata_int = 'h2f60;
    'h76c : romdata_int = 'h8a67;
    'h76d : romdata_int = 'h9a0e;
    'h76e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h76f : romdata_int = 'h1ccb;
    'h770 : romdata_int = 'h2c00;
    'h771 : romdata_int = 'h34f2;
    'h772 : romdata_int = 'h3b21;
    'h773 : romdata_int = 'h6d11;
    'h774 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h775 : romdata_int = 'he7d;
    'h776 : romdata_int = 'h2e00;
    'h777 : romdata_int = 'h3100;
    'h778 : romdata_int = 'h38fc;
    'h779 : romdata_int = 'h48a1;
    'h77a : romdata_int = 'h45a; // Line descriptor for 1_2
    'h77b : romdata_int = 'h1a97;
    'h77c : romdata_int = 'h1f13;
    'h77d : romdata_int = 'h3000;
    'h77e : romdata_int = 'h52b0;
    'h77f : romdata_int = 'h5938;
    'h780 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h781 : romdata_int = 'h465;
    'h782 : romdata_int = 'h2cf3;
    'h783 : romdata_int = 'h3200;
    'h784 : romdata_int = 'h60c7;
    'h785 : romdata_int = 'ha40a;
    'h786 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h787 : romdata_int = 'h43f;
    'h788 : romdata_int = 'h1b4b;
    'h789 : romdata_int = 'h3400;
    'h78a : romdata_int = 'h8062;
    'h78b : romdata_int = 'ha164;
    'h78c : romdata_int = 'h45a; // Line descriptor for 1_2
    'h78d : romdata_int = 'h20f3;
    'h78e : romdata_int = 'h3600;
    'h78f : romdata_int = 'h44fd;
    'h790 : romdata_int = 'h907c;
    'h791 : romdata_int = 'h994d;
    'h792 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h793 : romdata_int = 'h9f;
    'h794 : romdata_int = 'h131f;
    'h795 : romdata_int = 'h3800;
    'h796 : romdata_int = 'h44a7;
    'h797 : romdata_int = 'h6f62;
    'h798 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h799 : romdata_int = 'he9d;
    'h79a : romdata_int = 'h3602;
    'h79b : romdata_int = 'h3a00;
    'h79c : romdata_int = 'h42d9;
    'h79d : romdata_int = 'h7c0f;
    'h79e : romdata_int = 'h45a; // Line descriptor for 1_2
    'h79f : romdata_int = 'h16bd;
    'h7a0 : romdata_int = 'h2406;
    'h7a1 : romdata_int = 'h38f2;
    'h7a2 : romdata_int = 'h3c00;
    'h7a3 : romdata_int = 'h8b49;
    'h7a4 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7a5 : romdata_int = 'h12ed;
    'h7a6 : romdata_int = 'h14a2;
    'h7a7 : romdata_int = 'h3e00;
    'h7a8 : romdata_int = 'h3b4e;
    'h7a9 : romdata_int = 'h4242;
    'h7aa : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7ab : romdata_int = 'h114c;
    'h7ac : romdata_int = 'h2e76;
    'h7ad : romdata_int = 'h3f50;
    'h7ae : romdata_int = 'h4000;
    'h7af : romdata_int = 'h4144;
    'h7b0 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7b1 : romdata_int = 'h1703;
    'h7b2 : romdata_int = 'h3361;
    'h7b3 : romdata_int = 'h4200;
    'h7b4 : romdata_int = 'h54ec;
    'h7b5 : romdata_int = 'ha8f1;
    'h7b6 : romdata_int = 'h45a; // Line descriptor for 1_2
    'h7b7 : romdata_int = 'hab1;
    'h7b8 : romdata_int = 'he07;
    'h7b9 : romdata_int = 'h1e99;
    'h7ba : romdata_int = 'h4400;
    'h7bb : romdata_int = 'h70dd;
    'h7bc : romdata_int = 'h645a; // Line descriptor for 1_2
    'h7bd : romdata_int = 'h12a;
    'h7be : romdata_int = 'h26d8;
    'h7bf : romdata_int = 'h4166;
    'h7c0 : romdata_int = 'h4600;
    'h7c1 : romdata_int = 'h56a1;
    'h7c2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h7c3 : romdata_int = 'hed;
    'h7c4 : romdata_int = 'h1ec8;
    'h7c5 : romdata_int = 'h2d39;
    'h7c6 : romdata_int = 'h3086;
    'h7c7 : romdata_int = 'h4159;
    'h7c8 : romdata_int = 'h4272;
    'h7c9 : romdata_int = 'h4800;
    'h7ca : romdata_int = 'h50d1;
    'h7cb : romdata_int = 'hcacb;
    'h7cc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7cd : romdata_int = 'h9b;
    'h7ce : romdata_int = 'he8a;
    'h7cf : romdata_int = 'h121a;
    'h7d0 : romdata_int = 'h1706;
    'h7d1 : romdata_int = 'h3043;
    'h7d2 : romdata_int = 'h4286;
    'h7d3 : romdata_int = 'h4a00;
    'h7d4 : romdata_int = 'h584a;
    'h7d5 : romdata_int = 'hc35a;
    'h7d6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h7d7 : romdata_int = 'h565;
    'h7d8 : romdata_int = 'hd01;
    'h7d9 : romdata_int = 'h10b2;
    'h7da : romdata_int = 'h1c34;
    'h7db : romdata_int = 'h429c;
    'h7dc : romdata_int = 'h4423;
    'h7dd : romdata_int = 'h4c00;
    'h7de : romdata_int = 'h805e;
    'h7df : romdata_int = 'hb953;
    'h7e0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7e1 : romdata_int = 'h1947;
    'h7e2 : romdata_int = 'h22ba;
    'h7e3 : romdata_int = 'h22d9;
    'h7e4 : romdata_int = 'h2c91;
    'h7e5 : romdata_int = 'h3503;
    'h7e6 : romdata_int = 'h36f3;
    'h7e7 : romdata_int = 'h4e00;
    'h7e8 : romdata_int = 'h7367;
    'h7e9 : romdata_int = 'hd0d3;
    'h7ea : romdata_int = 'h848; // Line descriptor for 3_5
    'h7eb : romdata_int = 'hf61;
    'h7ec : romdata_int = 'h167d;
    'h7ed : romdata_int = 'h1c8b;
    'h7ee : romdata_int = 'h2432;
    'h7ef : romdata_int = 'h2479;
    'h7f0 : romdata_int = 'h3222;
    'h7f1 : romdata_int = 'h5000;
    'h7f2 : romdata_int = 'h6e17;
    'h7f3 : romdata_int = 'hc166;
    'h7f4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h7f5 : romdata_int = 'h2cd1;
    'h7f6 : romdata_int = 'h30d2;
    'h7f7 : romdata_int = 'h32a0;
    'h7f8 : romdata_int = 'h380b;
    'h7f9 : romdata_int = 'h3a35;
    'h7fa : romdata_int = 'h3e78;
    'h7fb : romdata_int = 'h5200;
    'h7fc : romdata_int = 'h60c9;
    'h7fd : romdata_int = 'hbc89;
    'h7fe : romdata_int = 'h848; // Line descriptor for 3_5
    'h7ff : romdata_int = 'hc55;
    'h800 : romdata_int = 'h14b4;
    'h801 : romdata_int = 'h1864;
    'h802 : romdata_int = 'h2360;
    'h803 : romdata_int = 'h28f5;
    'h804 : romdata_int = 'h331d;
    'h805 : romdata_int = 'h5400;
    'h806 : romdata_int = 'h64b8;
    'h807 : romdata_int = 'hc555;
    'h808 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h809 : romdata_int = 'h143e;
    'h80a : romdata_int = 'h24e4;
    'h80b : romdata_int = 'h32b8;
    'h80c : romdata_int = 'h372a;
    'h80d : romdata_int = 'h3c56;
    'h80e : romdata_int = 'h3e2c;
    'h80f : romdata_int = 'h5600;
    'h810 : romdata_int = 'h5b03;
    'h811 : romdata_int = 'hc31f;
    'h812 : romdata_int = 'h848; // Line descriptor for 3_5
    'h813 : romdata_int = 'h762;
    'h814 : romdata_int = 'h1062;
    'h815 : romdata_int = 'h1058;
    'h816 : romdata_int = 'h1079;
    'h817 : romdata_int = 'h2c38;
    'h818 : romdata_int = 'h46f6;
    'h819 : romdata_int = 'h4c82;
    'h81a : romdata_int = 'h5800;
    'h81b : romdata_int = 'h9f65;
    'h81c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h81d : romdata_int = 'h4e;
    'h81e : romdata_int = 'he75;
    'h81f : romdata_int = 'h169d;
    'h820 : romdata_int = 'h2c42;
    'h821 : romdata_int = 'h3d49;
    'h822 : romdata_int = 'h3ea9;
    'h823 : romdata_int = 'h5a00;
    'h824 : romdata_int = 'h8640;
    'h825 : romdata_int = 'h9b56;
    'h826 : romdata_int = 'h848; // Line descriptor for 3_5
    'h827 : romdata_int = 'h23a;
    'h828 : romdata_int = 'h1a3d;
    'h829 : romdata_int = 'h2251;
    'h82a : romdata_int = 'h2ebb;
    'h82b : romdata_int = 'h30ea;
    'h82c : romdata_int = 'h3c83;
    'h82d : romdata_int = 'h5c00;
    'h82e : romdata_int = 'h670b;
    'h82f : romdata_int = 'hce0d;
    'h830 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h831 : romdata_int = 'h86a;
    'h832 : romdata_int = 'h132c;
    'h833 : romdata_int = 'h165c;
    'h834 : romdata_int = 'h1688;
    'h835 : romdata_int = 'h1f50;
    'h836 : romdata_int = 'h20f3;
    'h837 : romdata_int = 'h5e00;
    'h838 : romdata_int = 'h703d;
    'h839 : romdata_int = 'ha520;
    'h83a : romdata_int = 'h848; // Line descriptor for 3_5
    'h83b : romdata_int = 'ha4a;
    'h83c : romdata_int = 'h16ca;
    'h83d : romdata_int = 'h1aa2;
    'h83e : romdata_int = 'h3318;
    'h83f : romdata_int = 'h435a;
    'h840 : romdata_int = 'h4667;
    'h841 : romdata_int = 'h5300;
    'h842 : romdata_int = 'h6000;
    'h843 : romdata_int = 'hbc72;
    'h844 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h845 : romdata_int = 'h65f;
    'h846 : romdata_int = 'h6dd;
    'h847 : romdata_int = 'he33;
    'h848 : romdata_int = 'h1f3f;
    'h849 : romdata_int = 'h3e28;
    'h84a : romdata_int = 'h44a3;
    'h84b : romdata_int = 'h4903;
    'h84c : romdata_int = 'h6200;
    'h84d : romdata_int = 'ha20e;
    'h84e : romdata_int = 'h848; // Line descriptor for 3_5
    'h84f : romdata_int = 'he41;
    'h850 : romdata_int = 'h1b1d;
    'h851 : romdata_int = 'h1e6f;
    'h852 : romdata_int = 'h234c;
    'h853 : romdata_int = 'h393e;
    'h854 : romdata_int = 'h3b60;
    'h855 : romdata_int = 'h6400;
    'h856 : romdata_int = 'h8a1c;
    'h857 : romdata_int = 'hb260;
    'h858 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h859 : romdata_int = 'h8c9;
    'h85a : romdata_int = 'h1e69;
    'h85b : romdata_int = 'h2f32;
    'h85c : romdata_int = 'h36e2;
    'h85d : romdata_int = 'h3e8f;
    'h85e : romdata_int = 'h4075;
    'h85f : romdata_int = 'h6600;
    'h860 : romdata_int = 'h78df;
    'h861 : romdata_int = 'ha0a7;
    'h862 : romdata_int = 'h848; // Line descriptor for 3_5
    'h863 : romdata_int = 'h1341;
    'h864 : romdata_int = 'h1af6;
    'h865 : romdata_int = 'h1e47;
    'h866 : romdata_int = 'h2700;
    'h867 : romdata_int = 'h3706;
    'h868 : romdata_int = 'h3a46;
    'h869 : romdata_int = 'h5356;
    'h86a : romdata_int = 'h6800;
    'h86b : romdata_int = 'hcc33;
    'h86c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h86d : romdata_int = 'h41e;
    'h86e : romdata_int = 'hb60;
    'h86f : romdata_int = 'h2e05;
    'h870 : romdata_int = 'h34cc;
    'h871 : romdata_int = 'h3b3f;
    'h872 : romdata_int = 'h4658;
    'h873 : romdata_int = 'h6a00;
    'h874 : romdata_int = 'h792c;
    'h875 : romdata_int = 'hb456;
    'h876 : romdata_int = 'h848; // Line descriptor for 3_5
    'h877 : romdata_int = 'h2e1;
    'h878 : romdata_int = 'h8f2;
    'h879 : romdata_int = 'h1c28;
    'h87a : romdata_int = 'h1c81;
    'h87b : romdata_int = 'h2854;
    'h87c : romdata_int = 'h2f50;
    'h87d : romdata_int = 'h6c00;
    'h87e : romdata_int = 'h753c;
    'h87f : romdata_int = 'hc6ac;
    'h880 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h881 : romdata_int = 'h4bc;
    'h882 : romdata_int = 'ha4e;
    'h883 : romdata_int = 'hf64;
    'h884 : romdata_int = 'h1268;
    'h885 : romdata_int = 'h3629;
    'h886 : romdata_int = 'h3e33;
    'h887 : romdata_int = 'h6e00;
    'h888 : romdata_int = 'h76c4;
    'h889 : romdata_int = 'hb6c1;
    'h88a : romdata_int = 'h848; // Line descriptor for 3_5
    'h88b : romdata_int = 'h479;
    'h88c : romdata_int = 'h1522;
    'h88d : romdata_int = 'h1733;
    'h88e : romdata_int = 'h267a;
    'h88f : romdata_int = 'h2ea6;
    'h890 : romdata_int = 'h4130;
    'h891 : romdata_int = 'h7000;
    'h892 : romdata_int = 'h7e70;
    'h893 : romdata_int = 'hb8b7;
    'h894 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h895 : romdata_int = 'h50b;
    'h896 : romdata_int = 'h6e6;
    'h897 : romdata_int = 'h950;
    'h898 : romdata_int = 'hc4b;
    'h899 : romdata_int = 'h1eb5;
    'h89a : romdata_int = 'h24e3;
    'h89b : romdata_int = 'h7200;
    'h89c : romdata_int = 'h7c08;
    'h89d : romdata_int = 'h9647;
    'h89e : romdata_int = 'h848; // Line descriptor for 3_5
    'h89f : romdata_int = 'h72e;
    'h8a0 : romdata_int = 'h223a;
    'h8a1 : romdata_int = 'h2ae6;
    'h8a2 : romdata_int = 'h348d;
    'h8a3 : romdata_int = 'h34d3;
    'h8a4 : romdata_int = 'h3b08;
    'h8a5 : romdata_int = 'h620a;
    'h8a6 : romdata_int = 'h7400;
    'h8a7 : romdata_int = 'hccec;
    'h8a8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8a9 : romdata_int = 'h2ec;
    'h8aa : romdata_int = 'h131d;
    'h8ab : romdata_int = 'h2721;
    'h8ac : romdata_int = 'h364d;
    'h8ad : romdata_int = 'h3639;
    'h8ae : romdata_int = 'h366e;
    'h8af : romdata_int = 'h550a;
    'h8b0 : romdata_int = 'h7600;
    'h8b1 : romdata_int = 'h9f30;
    'h8b2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h8b3 : romdata_int = 'h364;
    'h8b4 : romdata_int = 'hc7c;
    'h8b5 : romdata_int = 'h283e;
    'h8b6 : romdata_int = 'h2b52;
    'h8b7 : romdata_int = 'h3d32;
    'h8b8 : romdata_int = 'h4622;
    'h8b9 : romdata_int = 'h7800;
    'h8ba : romdata_int = 'h7d15;
    'h8bb : romdata_int = 'hac5a;
    'h8bc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8bd : romdata_int = 'h2f0;
    'h8be : romdata_int = 'h316;
    'h8bf : romdata_int = 'h16b0;
    'h8c0 : romdata_int = 'h22cf;
    'h8c1 : romdata_int = 'h3231;
    'h8c2 : romdata_int = 'h411c;
    'h8c3 : romdata_int = 'h66b8;
    'h8c4 : romdata_int = 'h7a00;
    'h8c5 : romdata_int = 'h993b;
    'h8c6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h8c7 : romdata_int = 'h2b;
    'h8c8 : romdata_int = 'h1d13;
    'h8c9 : romdata_int = 'h2030;
    'h8ca : romdata_int = 'h22d4;
    'h8cb : romdata_int = 'h391c;
    'h8cc : romdata_int = 'h4615;
    'h8cd : romdata_int = 'h6925;
    'h8ce : romdata_int = 'h7c00;
    'h8cf : romdata_int = 'h9860;
    'h8d0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8d1 : romdata_int = 'h1;
    'h8d2 : romdata_int = 'hcb5;
    'h8d3 : romdata_int = 'h14cf;
    'h8d4 : romdata_int = 'h20b5;
    'h8d5 : romdata_int = 'h4033;
    'h8d6 : romdata_int = 'h4632;
    'h8d7 : romdata_int = 'h5698;
    'h8d8 : romdata_int = 'h7e00;
    'h8d9 : romdata_int = 'ha6d3;
    'h8da : romdata_int = 'h848; // Line descriptor for 3_5
    'h8db : romdata_int = 'h44c;
    'h8dc : romdata_int = 'h1440;
    'h8dd : romdata_int = 'h14ab;
    'h8de : romdata_int = 'h2485;
    'h8df : romdata_int = 'h3d3a;
    'h8e0 : romdata_int = 'h40fd;
    'h8e1 : romdata_int = 'h5e65;
    'h8e2 : romdata_int = 'h8000;
    'h8e3 : romdata_int = 'h915b;
    'h8e4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8e5 : romdata_int = 'h53d;
    'h8e6 : romdata_int = 'hb18;
    'h8e7 : romdata_int = 'h14e4;
    'h8e8 : romdata_int = 'h1737;
    'h8e9 : romdata_int = 'h365e;
    'h8ea : romdata_int = 'h3ce4;
    'h8eb : romdata_int = 'h7695;
    'h8ec : romdata_int = 'h8200;
    'h8ed : romdata_int = 'h9726;
    'h8ee : romdata_int = 'h848; // Line descriptor for 3_5
    'h8ef : romdata_int = 'h137;
    'h8f0 : romdata_int = 'h1049;
    'h8f1 : romdata_int = 'h10f1;
    'h8f2 : romdata_int = 'h1acb;
    'h8f3 : romdata_int = 'h2d61;
    'h8f4 : romdata_int = 'h3b49;
    'h8f5 : romdata_int = 'h6b3c;
    'h8f6 : romdata_int = 'h8400;
    'h8f7 : romdata_int = 'hc633;
    'h8f8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h8f9 : romdata_int = 'h35c;
    'h8fa : romdata_int = 'h89a;
    'h8fb : romdata_int = 'h1480;
    'h8fc : romdata_int = 'h3517;
    'h8fd : romdata_int = 'h404b;
    'h8fe : romdata_int = 'h4296;
    'h8ff : romdata_int = 'h6854;
    'h900 : romdata_int = 'h8600;
    'h901 : romdata_int = 'haac7;
    'h902 : romdata_int = 'h848; // Line descriptor for 3_5
    'h903 : romdata_int = 'hd22;
    'h904 : romdata_int = 'hec5;
    'h905 : romdata_int = 'h2a13;
    'h906 : romdata_int = 'h2c87;
    'h907 : romdata_int = 'h2e8e;
    'h908 : romdata_int = 'h40df;
    'h909 : romdata_int = 'h84bc;
    'h90a : romdata_int = 'h8800;
    'h90b : romdata_int = 'hb07a;
    'h90c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h90d : romdata_int = 'h499;
    'h90e : romdata_int = 'h747;
    'h90f : romdata_int = 'h10c1;
    'h910 : romdata_int = 'h1d4d;
    'h911 : romdata_int = 'h2155;
    'h912 : romdata_int = 'h3d4f;
    'h913 : romdata_int = 'h4c95;
    'h914 : romdata_int = 'h8a00;
    'h915 : romdata_int = 'ha69c;
    'h916 : romdata_int = 'h848; // Line descriptor for 3_5
    'h917 : romdata_int = 'ha1;
    'h918 : romdata_int = 'h648;
    'h919 : romdata_int = 'hc5e;
    'h91a : romdata_int = 'h26b8;
    'h91b : romdata_int = 'h2e52;
    'h91c : romdata_int = 'h2eee;
    'h91d : romdata_int = 'h5707;
    'h91e : romdata_int = 'h8c00;
    'h91f : romdata_int = 'hc873;
    'h920 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h921 : romdata_int = 'h2;
    'h922 : romdata_int = 'h6a0;
    'h923 : romdata_int = 'h6ae;
    'h924 : romdata_int = 'h1aa4;
    'h925 : romdata_int = 'h314b;
    'h926 : romdata_int = 'h3744;
    'h927 : romdata_int = 'h4901;
    'h928 : romdata_int = 'h8e00;
    'h929 : romdata_int = 'hc0f1;
    'h92a : romdata_int = 'h848; // Line descriptor for 3_5
    'h92b : romdata_int = 'h20b;
    'h92c : romdata_int = 'h80f;
    'h92d : romdata_int = 'ha5a;
    'h92e : romdata_int = 'h1a0a;
    'h92f : romdata_int = 'h3029;
    'h930 : romdata_int = 'h3525;
    'h931 : romdata_int = 'h5f33;
    'h932 : romdata_int = 'h9000;
    'h933 : romdata_int = 'hd431;
    'h934 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h935 : romdata_int = 'h2a1;
    'h936 : romdata_int = 'had0;
    'h937 : romdata_int = 'h2067;
    'h938 : romdata_int = 'h234f;
    'h939 : romdata_int = 'h26ef;
    'h93a : romdata_int = 'h3065;
    'h93b : romdata_int = 'h823b;
    'h93c : romdata_int = 'h9200;
    'h93d : romdata_int = 'hcf13;
    'h93e : romdata_int = 'h848; // Line descriptor for 3_5
    'h93f : romdata_int = 'h133f;
    'h940 : romdata_int = 'h16fd;
    'h941 : romdata_int = 'h1915;
    'h942 : romdata_int = 'h3344;
    'h943 : romdata_int = 'h450a;
    'h944 : romdata_int = 'h46c0;
    'h945 : romdata_int = 'h5915;
    'h946 : romdata_int = 'h9400;
    'h947 : romdata_int = 'h9444;
    'h948 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h949 : romdata_int = 'h1e67;
    'h94a : romdata_int = 'h28e4;
    'h94b : romdata_int = 'h292f;
    'h94c : romdata_int = 'h2c77;
    'h94d : romdata_int = 'h3a7b;
    'h94e : romdata_int = 'h3c37;
    'h94f : romdata_int = 'h5520;
    'h950 : romdata_int = 'h9600;
    'h951 : romdata_int = 'hac21;
    'h952 : romdata_int = 'h848; // Line descriptor for 3_5
    'h953 : romdata_int = 'h166b;
    'h954 : romdata_int = 'h1e0f;
    'h955 : romdata_int = 'h28d5;
    'h956 : romdata_int = 'h2962;
    'h957 : romdata_int = 'h3215;
    'h958 : romdata_int = 'h3462;
    'h959 : romdata_int = 'h752e;
    'h95a : romdata_int = 'h9800;
    'h95b : romdata_int = 'hd0a8;
    'h95c : romdata_int = 'h4848; // Line descriptor for 3_5
    'h95d : romdata_int = 'h8e5;
    'h95e : romdata_int = 'h1228;
    'h95f : romdata_int = 'h330b;
    'h960 : romdata_int = 'h3355;
    'h961 : romdata_int = 'h3c48;
    'h962 : romdata_int = 'h455a;
    'h963 : romdata_int = 'h629a;
    'h964 : romdata_int = 'h9a00;
    'h965 : romdata_int = 'hbabb;
    'h966 : romdata_int = 'h848; // Line descriptor for 3_5
    'h967 : romdata_int = 'h28;
    'h968 : romdata_int = 'h49d;
    'h969 : romdata_int = 'h1418;
    'h96a : romdata_int = 'h2d47;
    'h96b : romdata_int = 'h3a8a;
    'h96c : romdata_int = 'h3f20;
    'h96d : romdata_int = 'h50b9;
    'h96e : romdata_int = 'h9c00;
    'h96f : romdata_int = 'ha351;
    'h970 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h971 : romdata_int = 'h8c4;
    'h972 : romdata_int = 'h1810;
    'h973 : romdata_int = 'h2470;
    'h974 : romdata_int = 'h30b5;
    'h975 : romdata_int = 'h4420;
    'h976 : romdata_int = 'h449c;
    'h977 : romdata_int = 'h8b10;
    'h978 : romdata_int = 'h9e00;
    'h979 : romdata_int = 'hb0c8;
    'h97a : romdata_int = 'h848; // Line descriptor for 3_5
    'h97b : romdata_int = 'h1037;
    'h97c : romdata_int = 'h112a;
    'h97d : romdata_int = 'h18ad;
    'h97e : romdata_int = 'h1f5e;
    'h97f : romdata_int = 'h28c7;
    'h980 : romdata_int = 'h3511;
    'h981 : romdata_int = 'h8084;
    'h982 : romdata_int = 'ha000;
    'h983 : romdata_int = 'ha4c2;
    'h984 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h985 : romdata_int = 'h42a;
    'h986 : romdata_int = 'h124e;
    'h987 : romdata_int = 'h2557;
    'h988 : romdata_int = 'h3c6b;
    'h989 : romdata_int = 'h3d37;
    'h98a : romdata_int = 'h4276;
    'h98b : romdata_int = 'h6f0d;
    'h98c : romdata_int = 'ha200;
    'h98d : romdata_int = 'hd428;
    'h98e : romdata_int = 'h848; // Line descriptor for 3_5
    'h98f : romdata_int = 'h101e;
    'h990 : romdata_int = 'h1158;
    'h991 : romdata_int = 'h30b6;
    'h992 : romdata_int = 'h314c;
    'h993 : romdata_int = 'h4259;
    'h994 : romdata_int = 'h4463;
    'h995 : romdata_int = 'h82f3;
    'h996 : romdata_int = 'h9a68;
    'h997 : romdata_int = 'ha400;
    'h998 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h999 : romdata_int = 'he7d;
    'h99a : romdata_int = 'h1a32;
    'h99b : romdata_int = 'h2b44;
    'h99c : romdata_int = 'h344e;
    'h99d : romdata_int = 'h3505;
    'h99e : romdata_int = 'h4627;
    'h99f : romdata_int = 'h6d12;
    'h9a0 : romdata_int = 'ha600;
    'h9a1 : romdata_int = 'hb638;
    'h9a2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9a3 : romdata_int = 'h923;
    'h9a4 : romdata_int = 'h1906;
    'h9a5 : romdata_int = 'h1b3e;
    'h9a6 : romdata_int = 'h2ab3;
    'h9a7 : romdata_int = 'h2b62;
    'h9a8 : romdata_int = 'h3736;
    'h9a9 : romdata_int = 'h8ef0;
    'h9aa : romdata_int = 'h90c1;
    'h9ab : romdata_int = 'ha800;
    'h9ac : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9ad : romdata_int = 'h734;
    'h9ae : romdata_int = 'h1312;
    'h9af : romdata_int = 'h1ab3;
    'h9b0 : romdata_int = 'h2818;
    'h9b1 : romdata_int = 'h2ef7;
    'h9b2 : romdata_int = 'h3838;
    'h9b3 : romdata_int = 'h7032;
    'h9b4 : romdata_int = 'h9338;
    'h9b5 : romdata_int = 'haa00;
    'h9b6 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9b7 : romdata_int = 'ha83;
    'h9b8 : romdata_int = 'hee9;
    'h9b9 : romdata_int = 'h1c0b;
    'h9ba : romdata_int = 'h28fc;
    'h9bb : romdata_int = 'h3b47;
    'h9bc : romdata_int = 'h4089;
    'h9bd : romdata_int = 'h4a29;
    'h9be : romdata_int = 'hac00;
    'h9bf : romdata_int = 'hd62f;
    'h9c0 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9c1 : romdata_int = 'h338;
    'h9c2 : romdata_int = 'h1916;
    'h9c3 : romdata_int = 'h1c45;
    'h9c4 : romdata_int = 'h2e4b;
    'h9c5 : romdata_int = 'h4308;
    'h9c6 : romdata_int = 'h4558;
    'h9c7 : romdata_int = 'h72b9;
    'h9c8 : romdata_int = 'ha8d7;
    'h9c9 : romdata_int = 'hae00;
    'h9ca : romdata_int = 'h848; // Line descriptor for 3_5
    'h9cb : romdata_int = 'he4c;
    'h9cc : romdata_int = 'h1c7a;
    'h9cd : romdata_int = 'h2a38;
    'h9ce : romdata_int = 'h2a75;
    'h9cf : romdata_int = 'h2edf;
    'h9d0 : romdata_int = 'h4291;
    'h9d1 : romdata_int = 'h4e6c;
    'h9d2 : romdata_int = 'haf5a;
    'h9d3 : romdata_int = 'hb000;
    'h9d4 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9d5 : romdata_int = 'h115;
    'h9d6 : romdata_int = 'hf4a;
    'h9d7 : romdata_int = 'h1221;
    'h9d8 : romdata_int = 'h1338;
    'h9d9 : romdata_int = 'h1a72;
    'h9da : romdata_int = 'h3844;
    'h9db : romdata_int = 'h7a33;
    'h9dc : romdata_int = 'h9cb1;
    'h9dd : romdata_int = 'hb200;
    'h9de : romdata_int = 'h848; // Line descriptor for 3_5
    'h9df : romdata_int = 'h20cb;
    'h9e0 : romdata_int = 'h2080;
    'h9e1 : romdata_int = 'h20e5;
    'h9e2 : romdata_int = 'h2233;
    'h9e3 : romdata_int = 'h275f;
    'h9e4 : romdata_int = 'h4023;
    'h9e5 : romdata_int = 'h8942;
    'h9e6 : romdata_int = 'hb400;
    'h9e7 : romdata_int = 'hd26b;
    'h9e8 : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9e9 : romdata_int = 'h259;
    'h9ea : romdata_int = 'h1923;
    'h9eb : romdata_int = 'h24e6;
    'h9ec : romdata_int = 'h366f;
    'h9ed : romdata_int = 'h3ab7;
    'h9ee : romdata_int = 'h3ea4;
    'h9ef : romdata_int = 'h7e4f;
    'h9f0 : romdata_int = 'hb600;
    'h9f1 : romdata_int = 'hcb16;
    'h9f2 : romdata_int = 'h848; // Line descriptor for 3_5
    'h9f3 : romdata_int = 'h1e41;
    'h9f4 : romdata_int = 'h2032;
    'h9f5 : romdata_int = 'h2559;
    'h9f6 : romdata_int = 'h2567;
    'h9f7 : romdata_int = 'h2c01;
    'h9f8 : romdata_int = 'h2c19;
    'h9f9 : romdata_int = 'h88a1;
    'h9fa : romdata_int = 'hb800;
    'h9fb : romdata_int = 'hd33c;
    'h9fc : romdata_int = 'h4848; // Line descriptor for 3_5
    'h9fd : romdata_int = 'h4ef;
    'h9fe : romdata_int = 'h1308;
    'h9ff : romdata_int = 'h1855;
    'ha00 : romdata_int = 'h20db;
    'ha01 : romdata_int = 'h2633;
    'ha02 : romdata_int = 'h4464;
    'ha03 : romdata_int = 'h7a58;
    'ha04 : romdata_int = 'haa82;
    'ha05 : romdata_int = 'hba00;
    'ha06 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha07 : romdata_int = 'h8e;
    'ha08 : romdata_int = 'ha0e;
    'ha09 : romdata_int = 'h32f4;
    'ha0a : romdata_int = 'h3864;
    'ha0b : romdata_int = 'h3e6e;
    'ha0c : romdata_int = 'h4428;
    'ha0d : romdata_int = 'h8618;
    'ha0e : romdata_int = 'hbc00;
    'ha0f : romdata_int = 'hbe15;
    'ha10 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha11 : romdata_int = 'h760;
    'ha12 : romdata_int = 'h894;
    'ha13 : romdata_int = 'hac5;
    'ha14 : romdata_int = 'h194c;
    'ha15 : romdata_int = 'h2149;
    'ha16 : romdata_int = 'h2646;
    'ha17 : romdata_int = 'h4eaa;
    'ha18 : romdata_int = 'h94ae;
    'ha19 : romdata_int = 'hbe00;
    'ha1a : romdata_int = 'h848; // Line descriptor for 3_5
    'ha1b : romdata_int = 'h4c7;
    'ha1c : romdata_int = 'hd34;
    'ha1d : romdata_int = 'h32fa;
    'ha1e : romdata_int = 'h3861;
    'ha1f : romdata_int = 'h429e;
    'ha20 : romdata_int = 'h46d0;
    'ha21 : romdata_int = 'h8ebe;
    'ha22 : romdata_int = 'ha00f;
    'ha23 : romdata_int = 'hc000;
    'ha24 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha25 : romdata_int = 'h711;
    'ha26 : romdata_int = 'hae7;
    'ha27 : romdata_int = 'h1d51;
    'ha28 : romdata_int = 'h251a;
    'ha29 : romdata_int = 'h28ad;
    'ha2a : romdata_int = 'h2b35;
    'ha2b : romdata_int = 'h64bf;
    'ha2c : romdata_int = 'hc200;
    'ha2d : romdata_int = 'hc812;
    'ha2e : romdata_int = 'h848; // Line descriptor for 3_5
    'ha2f : romdata_int = 'h72;
    'ha30 : romdata_int = 'h183c;
    'ha31 : romdata_int = 'h3b28;
    'ha32 : romdata_int = 'h3cb8;
    'ha33 : romdata_int = 'h409c;
    'ha34 : romdata_int = 'h42e3;
    'ha35 : romdata_int = 'h4a91;
    'ha36 : romdata_int = 'ha840;
    'ha37 : romdata_int = 'hc400;
    'ha38 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha39 : romdata_int = 'h339;
    'ha3a : romdata_int = 'h84e;
    'ha3b : romdata_int = 'h2d5c;
    'ha3c : romdata_int = 'h3953;
    'ha3d : romdata_int = 'h3f65;
    'ha3e : romdata_int = 'h413c;
    'ha3f : romdata_int = 'h8539;
    'ha40 : romdata_int = 'h925c;
    'ha41 : romdata_int = 'hc600;
    'ha42 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha43 : romdata_int = 'hc5f;
    'ha44 : romdata_int = 'h10e5;
    'ha45 : romdata_int = 'h1498;
    'ha46 : romdata_int = 'h2f25;
    'ha47 : romdata_int = 'h44e1;
    'ha48 : romdata_int = 'h4741;
    'ha49 : romdata_int = 'h5a9c;
    'ha4a : romdata_int = 'h9d52;
    'ha4b : romdata_int = 'hc800;
    'ha4c : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha4d : romdata_int = 'hf11;
    'ha4e : romdata_int = 'h1c99;
    'ha4f : romdata_int = 'h22eb;
    'ha50 : romdata_int = 'h34c2;
    'ha51 : romdata_int = 'h3eec;
    'ha52 : romdata_int = 'h4652;
    'ha53 : romdata_int = 'h8cbc;
    'ha54 : romdata_int = 'hca00;
    'ha55 : romdata_int = 'hd66b;
    'ha56 : romdata_int = 'h848; // Line descriptor for 3_5
    'ha57 : romdata_int = 'ha13;
    'ha58 : romdata_int = 'h2755;
    'ha59 : romdata_int = 'h28f2;
    'ha5a : romdata_int = 'h2a58;
    'ha5b : romdata_int = 'h3154;
    'ha5c : romdata_int = 'h3ac4;
    'ha5d : romdata_int = 'h8cba;
    'ha5e : romdata_int = 'haf56;
    'ha5f : romdata_int = 'hcc00;
    'ha60 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha61 : romdata_int = 'hcd9;
    'ha62 : romdata_int = 'hd2b;
    'ha63 : romdata_int = 'h1425;
    'ha64 : romdata_int = 'h3893;
    'ha65 : romdata_int = 'h424f;
    'ha66 : romdata_int = 'h44af;
    'ha67 : romdata_int = 'h5d1e;
    'ha68 : romdata_int = 'hb211;
    'ha69 : romdata_int = 'hce00;
    'ha6a : romdata_int = 'h848; // Line descriptor for 3_5
    'ha6b : romdata_int = 'h8d8;
    'ha6c : romdata_int = 'ha77;
    'ha6d : romdata_int = 'hc06;
    'ha6e : romdata_int = 'h1c6f;
    'ha6f : romdata_int = 'h233b;
    'ha70 : romdata_int = 'h34ad;
    'ha71 : romdata_int = 'h6a50;
    'ha72 : romdata_int = 'hbe53;
    'ha73 : romdata_int = 'hd000;
    'ha74 : romdata_int = 'h4848; // Line descriptor for 3_5
    'ha75 : romdata_int = 'h1761;
    'ha76 : romdata_int = 'h1958;
    'ha77 : romdata_int = 'h24ba;
    'ha78 : romdata_int = 'h271c;
    'ha79 : romdata_int = 'h38c6;
    'ha7a : romdata_int = 'h4607;
    'ha7b : romdata_int = 'h6131;
    'ha7c : romdata_int = 'hba54;
    'ha7d : romdata_int = 'hd200;
    'ha7e : romdata_int = 'h848; // Line descriptor for 3_5
    'ha7f : romdata_int = 'h1a9a;
    'ha80 : romdata_int = 'h2137;
    'ha81 : romdata_int = 'h2688;
    'ha82 : romdata_int = 'h3112;
    'ha83 : romdata_int = 'h380e;
    'ha84 : romdata_int = 'h383b;
    'ha85 : romdata_int = 'h5cd0;
    'ha86 : romdata_int = 'hb520;
    'ha87 : romdata_int = 'hd400;
    'ha88 : romdata_int = 'h6848; // Line descriptor for 3_5
    'ha89 : romdata_int = 'h140a;
    'ha8a : romdata_int = 'h1e4c;
    'ha8b : romdata_int = 'h26c4;
    'ha8c : romdata_int = 'h2a70;
    'ha8d : romdata_int = 'h2b21;
    'ha8e : romdata_int = 'h3f55;
    'ha8f : romdata_int = 'h6c3a;
    'ha90 : romdata_int = 'hc51d;
    'ha91 : romdata_int = 'hd600;
    'ha92 : romdata_int = 'h73c; // Line descriptor for 2_3
    'ha93 : romdata_int = 'h0;
    'ha94 : romdata_int = 'h4;
    'ha95 : romdata_int = 'h16ec;
    'ha96 : romdata_int = 'h18e6;
    'ha97 : romdata_int = 'h4f1c;
    'ha98 : romdata_int = 'h7800;
    'ha99 : romdata_int = 'h9ea5;
    'ha9a : romdata_int = 'h9ee8;
    'ha9b : romdata_int = 'h473c; // Line descriptor for 2_3
    'ha9c : romdata_int = 'h200;
    'ha9d : romdata_int = 'h6bd;
    'ha9e : romdata_int = 'hf37;
    'ha9f : romdata_int = 'h18ec;
    'haa0 : romdata_int = 'h22e1;
    'haa1 : romdata_int = 'h7a00;
    'haa2 : romdata_int = 'hde3d;
    'haa3 : romdata_int = 'he12e;
    'haa4 : romdata_int = 'h73c; // Line descriptor for 2_3
    'haa5 : romdata_int = 'h400;
    'haa6 : romdata_int = 'h1097;
    'haa7 : romdata_int = 'h1648;
    'haa8 : romdata_int = 'h4f3e;
    'haa9 : romdata_int = 'h5f5f;
    'haaa : romdata_int = 'h7c00;
    'haab : romdata_int = 'haa48;
    'haac : romdata_int = 'hea70;
    'haad : romdata_int = 'h473c; // Line descriptor for 2_3
    'haae : romdata_int = 'h334;
    'haaf : romdata_int = 'h600;
    'hab0 : romdata_int = 'h667;
    'hab1 : romdata_int = 'hce5;
    'hab2 : romdata_int = 'h2013;
    'hab3 : romdata_int = 'h7e00;
    'hab4 : romdata_int = 'hd50b;
    'hab5 : romdata_int = 'he52c;
    'hab6 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hab7 : romdata_int = 'h261;
    'hab8 : romdata_int = 'h4c9;
    'hab9 : romdata_int = 'h800;
    'haba : romdata_int = 'h3d53;
    'habb : romdata_int = 'h741f;
    'habc : romdata_int = 'h8000;
    'habd : romdata_int = 'h910a;
    'habe : romdata_int = 'h9c22;
    'habf : romdata_int = 'h473c; // Line descriptor for 2_3
    'hac0 : romdata_int = 'ha00;
    'hac1 : romdata_int = 'hb38;
    'hac2 : romdata_int = 'he5c;
    'hac3 : romdata_int = 'h129e;
    'hac4 : romdata_int = 'h72a4;
    'hac5 : romdata_int = 'h7c33;
    'hac6 : romdata_int = 'h8200;
    'hac7 : romdata_int = 'h84c1;
    'hac8 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hac9 : romdata_int = 'h89;
    'haca : romdata_int = 'hc00;
    'hacb : romdata_int = 'hc08;
    'hacc : romdata_int = 'h10d5;
    'hacd : romdata_int = 'h4660;
    'hace : romdata_int = 'h8400;
    'hacf : romdata_int = 'h8a14;
    'had0 : romdata_int = 'ha6a2;
    'had1 : romdata_int = 'h473c; // Line descriptor for 2_3
    'had2 : romdata_int = 'h2e;
    'had3 : romdata_int = 'h2e0;
    'had4 : romdata_int = 'he00;
    'had5 : romdata_int = 'hf58;
    'had6 : romdata_int = 'h1d0b;
    'had7 : romdata_int = 'h8600;
    'had8 : romdata_int = 'hb07b;
    'had9 : romdata_int = 'hc71e;
    'hada : romdata_int = 'h73c; // Line descriptor for 2_3
    'hadb : romdata_int = 'h1000;
    'hadc : romdata_int = 'h1406;
    'hadd : romdata_int = 'h16d2;
    'hade : romdata_int = 'h1a31;
    'hadf : romdata_int = 'h3ef3;
    'hae0 : romdata_int = 'h8800;
    'hae1 : romdata_int = 'hd654;
    'hae2 : romdata_int = 'hdd0d;
    'hae3 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hae4 : romdata_int = 'h948;
    'hae5 : romdata_int = 'hace;
    'hae6 : romdata_int = 'heb0;
    'hae7 : romdata_int = 'h1200;
    'hae8 : romdata_int = 'h5468;
    'hae9 : romdata_int = 'h8a00;
    'haea : romdata_int = 'hbc1a;
    'haeb : romdata_int = 'hcf33;
    'haec : romdata_int = 'h73c; // Line descriptor for 2_3
    'haed : romdata_int = 'hccf;
    'haee : romdata_int = 'he87;
    'haef : romdata_int = 'h1400;
    'haf0 : romdata_int = 'h4c44;
    'haf1 : romdata_int = 'h553d;
    'haf2 : romdata_int = 'h8c00;
    'haf3 : romdata_int = 'haa85;
    'haf4 : romdata_int = 'hbc7d;
    'haf5 : romdata_int = 'h473c; // Line descriptor for 2_3
    'haf6 : romdata_int = 'h477;
    'haf7 : romdata_int = 'hc5d;
    'haf8 : romdata_int = 'h103f;
    'haf9 : romdata_int = 'h1600;
    'hafa : romdata_int = 'h4344;
    'hafb : romdata_int = 'h8e00;
    'hafc : romdata_int = 'ha466;
    'hafd : romdata_int = 'hc203;
    'hafe : romdata_int = 'h73c; // Line descriptor for 2_3
    'haff : romdata_int = 'h6a6;
    'hb00 : romdata_int = 'h1351;
    'hb01 : romdata_int = 'h1800;
    'hb02 : romdata_int = 'h58c4;
    'hb03 : romdata_int = 'h7028;
    'hb04 : romdata_int = 'h7f30;
    'hb05 : romdata_int = 'h9000;
    'hb06 : romdata_int = 'hce8d;
    'hb07 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb08 : romdata_int = 'h137;
    'hb09 : romdata_int = 'h26b;
    'hb0a : romdata_int = 'h1643;
    'hb0b : romdata_int = 'h1a00;
    'hb0c : romdata_int = 'h5151;
    'hb0d : romdata_int = 'h82a9;
    'hb0e : romdata_int = 'h9200;
    'hb0f : romdata_int = 'h9804;
    'hb10 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb11 : romdata_int = 'h4d5;
    'hb12 : romdata_int = 'h92a;
    'hb13 : romdata_int = 'h1c00;
    'hb14 : romdata_int = 'h2ed2;
    'hb15 : romdata_int = 'h3711;
    'hb16 : romdata_int = 'h9400;
    'hb17 : romdata_int = 'h9a15;
    'hb18 : romdata_int = 'ha45a;
    'hb19 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb1a : romdata_int = 'h44a;
    'hb1b : romdata_int = 'h140f;
    'hb1c : romdata_int = 'h1e00;
    'hb1d : romdata_int = 'h3325;
    'hb1e : romdata_int = 'h7120;
    'hb1f : romdata_int = 'h8e9c;
    'hb20 : romdata_int = 'h9600;
    'hb21 : romdata_int = 'hd725;
    'hb22 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb23 : romdata_int = 'h6f2;
    'hb24 : romdata_int = 'h14e2;
    'hb25 : romdata_int = 'h2000;
    'hb26 : romdata_int = 'h2767;
    'hb27 : romdata_int = 'h4408;
    'hb28 : romdata_int = 'h9800;
    'hb29 : romdata_int = 'had04;
    'hb2a : romdata_int = 'hcc54;
    'hb2b : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb2c : romdata_int = 'h52b;
    'hb2d : romdata_int = 'ha21;
    'hb2e : romdata_int = 'hcc0;
    'hb2f : romdata_int = 'h2200;
    'hb30 : romdata_int = 'h4446;
    'hb31 : romdata_int = 'h9a00;
    'hb32 : romdata_int = 'h9cf6;
    'hb33 : romdata_int = 'hd850;
    'hb34 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb35 : romdata_int = 'hafd;
    'hb36 : romdata_int = 'h1313;
    'hb37 : romdata_int = 'h2400;
    'hb38 : romdata_int = 'h3a6f;
    'hb39 : romdata_int = 'h4c61;
    'hb3a : romdata_int = 'h8497;
    'hb3b : romdata_int = 'h9c00;
    'hb3c : romdata_int = 'hb159;
    'hb3d : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb3e : romdata_int = 'hb0;
    'hb3f : romdata_int = 'h134d;
    'hb40 : romdata_int = 'h2600;
    'hb41 : romdata_int = 'h5ec4;
    'hb42 : romdata_int = 'h6437;
    'hb43 : romdata_int = 'h8659;
    'hb44 : romdata_int = 'h9e00;
    'hb45 : romdata_int = 'ha85b;
    'hb46 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb47 : romdata_int = 'h255;
    'hb48 : romdata_int = 'ha1c;
    'hb49 : romdata_int = 'h2096;
    'hb4a : romdata_int = 'h2800;
    'hb4b : romdata_int = 'h5949;
    'hb4c : romdata_int = 'h7a9c;
    'hb4d : romdata_int = 'ha000;
    'hb4e : romdata_int = 'hb42b;
    'hb4f : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb50 : romdata_int = 'heca;
    'hb51 : romdata_int = 'hf33;
    'hb52 : romdata_int = 'h2a00;
    'hb53 : romdata_int = 'h3874;
    'hb54 : romdata_int = 'h48af;
    'hb55 : romdata_int = 'ha200;
    'hb56 : romdata_int = 'ha2a5;
    'hb57 : romdata_int = 'haf03;
    'hb58 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb59 : romdata_int = 'h688;
    'hb5a : romdata_int = 'h10a1;
    'hb5b : romdata_int = 'h2c00;
    'hb5c : romdata_int = 'h60a1;
    'hb5d : romdata_int = 'h6e56;
    'hb5e : romdata_int = 'h8c12;
    'hb5f : romdata_int = 'h9485;
    'hb60 : romdata_int = 'ha400;
    'hb61 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb62 : romdata_int = 'h10b;
    'hb63 : romdata_int = 'h866;
    'hb64 : romdata_int = 'h16aa;
    'hb65 : romdata_int = 'h2e00;
    'hb66 : romdata_int = 'h6a63;
    'hb67 : romdata_int = 'ha600;
    'hb68 : romdata_int = 'he633;
    'hb69 : romdata_int = 'he658;
    'hb6a : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb6b : romdata_int = 'h464;
    'hb6c : romdata_int = 'h10fe;
    'hb6d : romdata_int = 'h1766;
    'hb6e : romdata_int = 'h3000;
    'hb6f : romdata_int = 'h5b47;
    'hb70 : romdata_int = 'h8896;
    'hb71 : romdata_int = 'ha800;
    'hb72 : romdata_int = 'hb339;
    'hb73 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb74 : romdata_int = 'h86;
    'hb75 : romdata_int = 'h2e6;
    'hb76 : romdata_int = 'h1345;
    'hb77 : romdata_int = 'h3200;
    'hb78 : romdata_int = 'h4ac6;
    'hb79 : romdata_int = 'haa00;
    'hb7a : romdata_int = 'hc537;
    'hb7b : romdata_int = 'hd310;
    'hb7c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb7d : romdata_int = 'h8;
    'hb7e : romdata_int = 'h858;
    'hb7f : romdata_int = 'h3400;
    'hb80 : romdata_int = 'h6c7a;
    'hb81 : romdata_int = 'h6cc3;
    'hb82 : romdata_int = 'h9b41;
    'hb83 : romdata_int = 'ha32f;
    'hb84 : romdata_int = 'hac00;
    'hb85 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb86 : romdata_int = 'h31e;
    'hb87 : romdata_int = 'h916;
    'hb88 : romdata_int = 'h3600;
    'hb89 : romdata_int = 'h3cd8;
    'hb8a : romdata_int = 'h746f;
    'hb8b : romdata_int = 'h9064;
    'hb8c : romdata_int = 'hae00;
    'hb8d : romdata_int = 'hc098;
    'hb8e : romdata_int = 'h73c; // Line descriptor for 2_3
    'hb8f : romdata_int = 'h536;
    'hb90 : romdata_int = 'h143a;
    'hb91 : romdata_int = 'h144c;
    'hb92 : romdata_int = 'h2ca7;
    'hb93 : romdata_int = 'h3800;
    'hb94 : romdata_int = 'hb000;
    'hb95 : romdata_int = 'hd2d4;
    'hb96 : romdata_int = 'he295;
    'hb97 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hb98 : romdata_int = 'h1299;
    'hb99 : romdata_int = 'h1689;
    'hb9a : romdata_int = 'h387b;
    'hb9b : romdata_int = 'h3a00;
    'hb9c : romdata_int = 'h6e5d;
    'hb9d : romdata_int = 'h92f6;
    'hb9e : romdata_int = 'hb200;
    'hb9f : romdata_int = 'hb72a;
    'hba0 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hba1 : romdata_int = 'hb19;
    'hba2 : romdata_int = 'h126f;
    'hba3 : romdata_int = 'h2424;
    'hba4 : romdata_int = 'h3c00;
    'hba5 : romdata_int = 'h4679;
    'hba6 : romdata_int = 'hac5c;
    'hba7 : romdata_int = 'hb400;
    'hba8 : romdata_int = 'hc315;
    'hba9 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbaa : romdata_int = 'h84d;
    'hbab : romdata_int = 'hd22;
    'hbac : romdata_int = 'heee;
    'hbad : romdata_int = 'h160a;
    'hbae : romdata_int = 'h3e00;
    'hbaf : romdata_int = 'hb600;
    'hbb0 : romdata_int = 'hc838;
    'hbb1 : romdata_int = 'hea4f;
    'hbb2 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbb3 : romdata_int = 'h2d5;
    'hbb4 : romdata_int = 'ha2a;
    'hbb5 : romdata_int = 'he88;
    'hbb6 : romdata_int = 'h16ea;
    'hbb7 : romdata_int = 'h4000;
    'hbb8 : romdata_int = 'h926b;
    'hbb9 : romdata_int = 'ha007;
    'hbba : romdata_int = 'hb800;
    'hbbb : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbbc : romdata_int = 'h28a;
    'hbbd : romdata_int = 'h127a;
    'hbbe : romdata_int = 'h14b8;
    'hbbf : romdata_int = 'h3462;
    'hbc0 : romdata_int = 'h4200;
    'hbc1 : romdata_int = 'hba00;
    'hbc2 : romdata_int = 'hd0c9;
    'hbc3 : romdata_int = 'he2c4;
    'hbc4 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbc5 : romdata_int = 'h722;
    'hbc6 : romdata_int = 'hec3;
    'hbc7 : romdata_int = 'h4400;
    'hbc8 : romdata_int = 'h6883;
    'hbc9 : romdata_int = 'h7355;
    'hbca : romdata_int = 'h82b2;
    'hbcb : romdata_int = 'h8b10;
    'hbcc : romdata_int = 'hbc00;
    'hbcd : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbce : romdata_int = 'h462;
    'hbcf : romdata_int = 'h16ce;
    'hbd0 : romdata_int = 'h2e08;
    'hbd1 : romdata_int = 'h348d;
    'hbd2 : romdata_int = 'h4600;
    'hbd3 : romdata_int = 'h889e;
    'hbd4 : romdata_int = 'hbe00;
    'hbd5 : romdata_int = 'hd93c;
    'hbd6 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbd7 : romdata_int = 'h65c;
    'hbd8 : romdata_int = 'hac9;
    'hbd9 : romdata_int = 'h26cb;
    'hbda : romdata_int = 'h4800;
    'hbdb : romdata_int = 'h6648;
    'hbdc : romdata_int = 'h8f5a;
    'hbdd : romdata_int = 'hb66c;
    'hbde : romdata_int = 'hc000;
    'hbdf : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbe0 : romdata_int = 'h554;
    'hbe1 : romdata_int = 'h749;
    'hbe2 : romdata_int = 'h1281;
    'hbe3 : romdata_int = 'h294b;
    'hbe4 : romdata_int = 'h4a00;
    'hbe5 : romdata_int = 'hc200;
    'hbe6 : romdata_int = 'hc503;
    'hbe7 : romdata_int = 'hc75c;
    'hbe8 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbe9 : romdata_int = 'h8f3;
    'hbea : romdata_int = 'h128b;
    'hbeb : romdata_int = 'h2a84;
    'hbec : romdata_int = 'h412a;
    'hbed : romdata_int = 'h4c00;
    'hbee : romdata_int = 'hb801;
    'hbef : romdata_int = 'hc400;
    'hbf0 : romdata_int = 'hcc99;
    'hbf1 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hbf2 : romdata_int = 'h9a;
    'hbf3 : romdata_int = 'h174c;
    'hbf4 : romdata_int = 'h3b09;
    'hbf5 : romdata_int = 'h4b53;
    'hbf6 : romdata_int = 'h4e00;
    'hbf7 : romdata_int = 'hbb56;
    'hbf8 : romdata_int = 'hc600;
    'hbf9 : romdata_int = 'hde32;
    'hbfa : romdata_int = 'h73c; // Line descriptor for 2_3
    'hbfb : romdata_int = 'h2a5;
    'hbfc : romdata_int = 'he45;
    'hbfd : romdata_int = 'h2d09;
    'hbfe : romdata_int = 'h5000;
    'hbff : romdata_int = 'h6a48;
    'hc00 : romdata_int = 'hbf0a;
    'hc01 : romdata_int = 'hc800;
    'hc02 : romdata_int = 'hec84;
    'hc03 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc04 : romdata_int = 'h490;
    'hc05 : romdata_int = 'hf06;
    'hc06 : romdata_int = 'h308d;
    'hc07 : romdata_int = 'h5200;
    'hc08 : romdata_int = 'h5c3a;
    'hc09 : romdata_int = 'h8098;
    'hc0a : romdata_int = 'haeb1;
    'hc0b : romdata_int = 'hca00;
    'hc0c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc0d : romdata_int = 'hb08;
    'hc0e : romdata_int = 'h1550;
    'hc0f : romdata_int = 'h1eb8;
    'hc10 : romdata_int = 'h5400;
    'hc11 : romdata_int = 'h60d9;
    'hc12 : romdata_int = 'h8104;
    'hc13 : romdata_int = 'h96f5;
    'hc14 : romdata_int = 'hcc00;
    'hc15 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc16 : romdata_int = 'hc18;
    'hc17 : romdata_int = 'h1234;
    'hc18 : romdata_int = 'h36ad;
    'hc19 : romdata_int = 'h426f;
    'hc1a : romdata_int = 'h5600;
    'hc1b : romdata_int = 'hc0ab;
    'hc1c : romdata_int = 'hce00;
    'hc1d : romdata_int = 'hdb12;
    'hc1e : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc1f : romdata_int = 'h267;
    'hc20 : romdata_int = 'h958;
    'hc21 : romdata_int = 'h3317;
    'hc22 : romdata_int = 'h5800;
    'hc23 : romdata_int = 'h7756;
    'hc24 : romdata_int = 'hb495;
    'hc25 : romdata_int = 'hba3d;
    'hc26 : romdata_int = 'hd000;
    'hc27 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc28 : romdata_int = 'hceb;
    'hc29 : romdata_int = 'h14b5;
    'hc2a : romdata_int = 'h4894;
    'hc2b : romdata_int = 'h5342;
    'hc2c : romdata_int = 'h5a00;
    'hc2d : romdata_int = 'h9832;
    'hc2e : romdata_int = 'ha8c8;
    'hc2f : romdata_int = 'hd200;
    'hc30 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc31 : romdata_int = 'hd5;
    'hc32 : romdata_int = 'h1140;
    'hc33 : romdata_int = 'h1f55;
    'hc34 : romdata_int = 'h5345;
    'hc35 : romdata_int = 'h5c00;
    'hc36 : romdata_int = 'h792f;
    'hc37 : romdata_int = 'h7a89;
    'hc38 : romdata_int = 'hd400;
    'hc39 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc3a : romdata_int = 'hc40;
    'hc3b : romdata_int = 'hcfd;
    'hc3c : romdata_int = 'h1aa0;
    'hc3d : romdata_int = 'h5e00;
    'hc3e : romdata_int = 'h64b8;
    'hc3f : romdata_int = 'h791e;
    'hc40 : romdata_int = 'hd600;
    'hc41 : romdata_int = 'he4df;
    'hc42 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc43 : romdata_int = 'h15c;
    'hc44 : romdata_int = 'h81a;
    'hc45 : romdata_int = 'h2419;
    'hc46 : romdata_int = 'h5a7b;
    'hc47 : romdata_int = 'h6000;
    'hc48 : romdata_int = 'hb8b9;
    'hc49 : romdata_int = 'hd800;
    'hc4a : romdata_int = 'he915;
    'hc4b : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc4c : romdata_int = 'h727;
    'hc4d : romdata_int = 'ha33;
    'hc4e : romdata_int = 'h146f;
    'hc4f : romdata_int = 'h2a45;
    'hc50 : romdata_int = 'h6200;
    'hc51 : romdata_int = 'h96ea;
    'hc52 : romdata_int = 'hda00;
    'hc53 : romdata_int = 'hee3b;
    'hc54 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc55 : romdata_int = 'h4b6;
    'hc56 : romdata_int = 'h10a6;
    'hc57 : romdata_int = 'h308c;
    'hc58 : romdata_int = 'h3e29;
    'hc59 : romdata_int = 'h6400;
    'hc5a : romdata_int = 'hdc00;
    'hc5b : romdata_int = 'he13c;
    'hc5c : romdata_int = 'heef3;
    'hc5d : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc5e : romdata_int = 'hae;
    'hc5f : romdata_int = 'ha50;
    'hc60 : romdata_int = 'hc65;
    'hc61 : romdata_int = 'h1560;
    'hc62 : romdata_int = 'h6600;
    'hc63 : romdata_int = 'h9535;
    'hc64 : romdata_int = 'hde00;
    'hc65 : romdata_int = 'he808;
    'hc66 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc67 : romdata_int = 'h734;
    'hc68 : romdata_int = 'h10a8;
    'hc69 : romdata_int = 'h50cd;
    'hc6a : romdata_int = 'h673a;
    'hc6b : romdata_int = 'h6800;
    'hc6c : romdata_int = 'hbec2;
    'hc6d : romdata_int = 'hcb4e;
    'hc6e : romdata_int = 'he000;
    'hc6f : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc70 : romdata_int = 'hc7b;
    'hc71 : romdata_int = 'h1511;
    'hc72 : romdata_int = 'h1cf4;
    'hc73 : romdata_int = 'h573f;
    'hc74 : romdata_int = 'h6a00;
    'hc75 : romdata_int = 'h7c75;
    'hc76 : romdata_int = 'hd159;
    'hc77 : romdata_int = 'he200;
    'hc78 : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc79 : romdata_int = 'h105a;
    'hc7a : romdata_int = 'h1744;
    'hc7b : romdata_int = 'h2242;
    'hc7c : romdata_int = 'h6294;
    'hc7d : romdata_int = 'h6c00;
    'hc7e : romdata_int = 'h8cf9;
    'hc7f : romdata_int = 'ha07a;
    'hc80 : romdata_int = 'he400;
    'hc81 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc82 : romdata_int = 'h8ee;
    'hc83 : romdata_int = 'h10b1;
    'hc84 : romdata_int = 'h2822;
    'hc85 : romdata_int = 'h406e;
    'hc86 : romdata_int = 'h6e00;
    'hc87 : romdata_int = 'hd4b8;
    'hc88 : romdata_int = 'he600;
    'hc89 : romdata_int = 'hec5e;
    'hc8a : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc8b : romdata_int = 'h4f2;
    'hc8c : romdata_int = 'h120b;
    'hc8d : romdata_int = 'h5d0b;
    'hc8e : romdata_int = 'h7000;
    'hc8f : romdata_int = 'h7656;
    'hc90 : romdata_int = 'hc846;
    'hc91 : romdata_int = 'hda3a;
    'hc92 : romdata_int = 'he800;
    'hc93 : romdata_int = 'h473c; // Line descriptor for 2_3
    'hc94 : romdata_int = 'h701;
    'hc95 : romdata_int = 'h1447;
    'hc96 : romdata_int = 'h56b7;
    'hc97 : romdata_int = 'h6256;
    'hc98 : romdata_int = 'h7200;
    'hc99 : romdata_int = 'h7edf;
    'hc9a : romdata_int = 'ha6a7;
    'hc9b : romdata_int = 'hea00;
    'hc9c : romdata_int = 'h73c; // Line descriptor for 2_3
    'hc9d : romdata_int = 'h832;
    'hc9e : romdata_int = 'haa2;
    'hc9f : romdata_int = 'h114b;
    'hca0 : romdata_int = 'h6840;
    'hca1 : romdata_int = 'h7400;
    'hca2 : romdata_int = 'h869c;
    'hca3 : romdata_int = 'hb229;
    'hca4 : romdata_int = 'hec00;
    'hca5 : romdata_int = 'h673c; // Line descriptor for 2_3
    'hca6 : romdata_int = 'h328;
    'hca7 : romdata_int = 'h648;
    'hca8 : romdata_int = 'h80a;
    'hca9 : romdata_int = 'h10f5;
    'hcaa : romdata_int = 'h7600;
    'hcab : romdata_int = 'hcb1e;
    'hcac : romdata_int = 'hdc17;
    'hcad : romdata_int = 'hee00;
    'hcae : romdata_int = 'hb2d; // Line descriptor for 3_4
    'hcaf : romdata_int = 'h0;
    'hcb0 : romdata_int = 'h534;
    'hcb1 : romdata_int = 'h69b;
    'hcb2 : romdata_int = 'hcd7;
    'hcb3 : romdata_int = 'h14c4;
    'hcb4 : romdata_int = 'h3e61;
    'hcb5 : romdata_int = 'h5a00;
    'hcb6 : romdata_int = 'h76bb;
    'hcb7 : romdata_int = 'h8a3b;
    'hcb8 : romdata_int = 'hb400;
    'hcb9 : romdata_int = 'hbcad;
    'hcba : romdata_int = 'hfd1a;
    'hcbb : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcbc : romdata_int = 'h200;
    'hcbd : romdata_int = 'h651;
    'hcbe : romdata_int = 'he09;
    'hcbf : romdata_int = 'h122e;
    'hcc0 : romdata_int = 'h4f3e;
    'hcc1 : romdata_int = 'h50b5;
    'hcc2 : romdata_int = 'h5c00;
    'hcc3 : romdata_int = 'h7d0c;
    'hcc4 : romdata_int = 'ha4d1;
    'hcc5 : romdata_int = 'hb600;
    'hcc6 : romdata_int = 'he34b;
    'hcc7 : romdata_int = 'h102b4;
    'hcc8 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcc9 : romdata_int = 'h296;
    'hcca : romdata_int = 'h400;
    'hccb : romdata_int = 'h50f;
    'hccc : romdata_int = 'hf52;
    'hccd : romdata_int = 'h3c46;
    'hcce : romdata_int = 'h515b;
    'hccf : romdata_int = 'h5e00;
    'hcd0 : romdata_int = 'h66b0;
    'hcd1 : romdata_int = 'hab47;
    'hcd2 : romdata_int = 'hb49d;
    'hcd3 : romdata_int = 'hb800;
    'hcd4 : romdata_int = 'he54c;
    'hcd5 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcd6 : romdata_int = 'h600;
    'hcd7 : romdata_int = 'ha8c;
    'hcd8 : romdata_int = 'he58;
    'hcd9 : romdata_int = 'h100c;
    'hcda : romdata_int = 'h1135;
    'hcdb : romdata_int = 'h2323;
    'hcdc : romdata_int = 'h6000;
    'hcdd : romdata_int = 'h6106;
    'hcde : romdata_int = 'h649b;
    'hcdf : romdata_int = 'hba00;
    'hce0 : romdata_int = 'hf6a5;
    'hce1 : romdata_int = 'h10c40;
    'hce2 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hce3 : romdata_int = 'h541;
    'hce4 : romdata_int = 'h800;
    'hce5 : romdata_int = 'h149d;
    'hce6 : romdata_int = 'h175b;
    'hce7 : romdata_int = 'h3abf;
    'hce8 : romdata_int = 'h4829;
    'hce9 : romdata_int = 'h5a1c;
    'hcea : romdata_int = 'h5d18;
    'hceb : romdata_int = 'h6200;
    'hcec : romdata_int = 'hbc00;
    'hced : romdata_int = 'hc814;
    'hcee : romdata_int = 'hd6bd;
    'hcef : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcf0 : romdata_int = 'ha1f;
    'hcf1 : romdata_int = 'ha00;
    'hcf2 : romdata_int = 'hb16;
    'hcf3 : romdata_int = 'h12a1;
    'hcf4 : romdata_int = 'h3c4d;
    'hcf5 : romdata_int = 'h4131;
    'hcf6 : romdata_int = 'h6400;
    'hcf7 : romdata_int = 'h9364;
    'hcf8 : romdata_int = 'h9b0d;
    'hcf9 : romdata_int = 'hbc1f;
    'hcfa : romdata_int = 'hbe00;
    'hcfb : romdata_int = 'h10750;
    'hcfc : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hcfd : romdata_int = 'hb3b;
    'hcfe : romdata_int = 'hc00;
    'hcff : romdata_int = 'h10cc;
    'hd00 : romdata_int = 'h120c;
    'hd01 : romdata_int = 'h18c2;
    'hd02 : romdata_int = 'h212a;
    'hd03 : romdata_int = 'h6046;
    'hd04 : romdata_int = 'h6600;
    'hd05 : romdata_int = 'hb28a;
    'hd06 : romdata_int = 'hc000;
    'hd07 : romdata_int = 'hc46b;
    'hd08 : romdata_int = 'hd43d;
    'hd09 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd0a : romdata_int = 'he00;
    'hd0b : romdata_int = 'h1319;
    'hd0c : romdata_int = 'h1a96;
    'hd0d : romdata_int = 'h1cb5;
    'hd0e : romdata_int = 'h26a0;
    'hd0f : romdata_int = 'h433b;
    'hd10 : romdata_int = 'h5e3c;
    'hd11 : romdata_int = 'h6800;
    'hd12 : romdata_int = 'h8457;
    'hd13 : romdata_int = 'hc200;
    'hd14 : romdata_int = 'hd8c6;
    'hd15 : romdata_int = 'hf72b;
    'hd16 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd17 : romdata_int = 'h824;
    'hd18 : romdata_int = 'h1000;
    'hd19 : romdata_int = 'h104f;
    'hd1a : romdata_int = 'h14e0;
    'hd1b : romdata_int = 'h1948;
    'hd1c : romdata_int = 'h2a62;
    'hd1d : romdata_int = 'h6a00;
    'hd1e : romdata_int = 'h6e27;
    'hd1f : romdata_int = 'hb2ab;
    'hd20 : romdata_int = 'hc0ab;
    'hd21 : romdata_int = 'hc400;
    'hd22 : romdata_int = 'he892;
    'hd23 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd24 : romdata_int = 'h333;
    'hd25 : romdata_int = 'h48e;
    'hd26 : romdata_int = 'h8f0;
    'hd27 : romdata_int = 'hc5a;
    'hd28 : romdata_int = 'h1200;
    'hd29 : romdata_int = 'h3b1d;
    'hd2a : romdata_int = 'h6c00;
    'hd2b : romdata_int = 'h720c;
    'hd2c : romdata_int = 'hae1a;
    'hd2d : romdata_int = 'hc600;
    'hd2e : romdata_int = 'hd90f;
    'hd2f : romdata_int = 'hde59;
    'hd30 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd31 : romdata_int = 'h354;
    'hd32 : romdata_int = 'h86c;
    'hd33 : romdata_int = 'h1293;
    'hd34 : romdata_int = 'h1400;
    'hd35 : romdata_int = 'h1851;
    'hd36 : romdata_int = 'h1a0b;
    'hd37 : romdata_int = 'h6e00;
    'hd38 : romdata_int = 'h7eb3;
    'hd39 : romdata_int = 'h9d58;
    'hd3a : romdata_int = 'hc709;
    'hd3b : romdata_int = 'hc800;
    'hd3c : romdata_int = 'hc828;
    'hd3d : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd3e : romdata_int = 'h12;
    'hd3f : romdata_int = 'ha78;
    'hd40 : romdata_int = 'h1080;
    'hd41 : romdata_int = 'h1600;
    'hd42 : romdata_int = 'h1f0a;
    'hd43 : romdata_int = 'h2ea8;
    'hd44 : romdata_int = 'h7000;
    'hd45 : romdata_int = 'h7026;
    'hd46 : romdata_int = 'h7314;
    'hd47 : romdata_int = 'hc239;
    'hd48 : romdata_int = 'hca00;
    'hd49 : romdata_int = 'hf510;
    'hd4a : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd4b : romdata_int = 'h48;
    'hd4c : romdata_int = 'h4b1;
    'hd4d : romdata_int = 'h1800;
    'hd4e : romdata_int = 'h186d;
    'hd4f : romdata_int = 'h1a3a;
    'hd50 : romdata_int = 'h3f35;
    'hd51 : romdata_int = 'h694f;
    'hd52 : romdata_int = 'h7200;
    'hd53 : romdata_int = 'h98d5;
    'hd54 : romdata_int = 'hb44d;
    'hd55 : romdata_int = 'hcc00;
    'hd56 : romdata_int = 'hd0ae;
    'hd57 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd58 : romdata_int = 'h8ce;
    'hd59 : romdata_int = 'h14cd;
    'hd5a : romdata_int = 'h162a;
    'hd5b : romdata_int = 'h1a00;
    'hd5c : romdata_int = 'h1ac6;
    'hd5d : romdata_int = 'h52f9;
    'hd5e : romdata_int = 'h6a70;
    'hd5f : romdata_int = 'h7400;
    'hd60 : romdata_int = 'h8827;
    'hd61 : romdata_int = 'hce00;
    'hd62 : romdata_int = 'hd667;
    'hd63 : romdata_int = 'hdd18;
    'hd64 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd65 : romdata_int = 'h706;
    'hd66 : romdata_int = 'h8d7;
    'hd67 : romdata_int = 'h1962;
    'hd68 : romdata_int = 'h1b26;
    'hd69 : romdata_int = 'h1c00;
    'hd6a : romdata_int = 'h2c3b;
    'hd6b : romdata_int = 'h6765;
    'hd6c : romdata_int = 'h7600;
    'hd6d : romdata_int = 'h7c1f;
    'hd6e : romdata_int = 'hd000;
    'hd6f : romdata_int = 'hd287;
    'hd70 : romdata_int = 'he8be;
    'hd71 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd72 : romdata_int = 'h81b;
    'hd73 : romdata_int = 'hf0b;
    'hd74 : romdata_int = 'h1492;
    'hd75 : romdata_int = 'h1e00;
    'hd76 : romdata_int = 'h2541;
    'hd77 : romdata_int = 'h3488;
    'hd78 : romdata_int = 'h7800;
    'hd79 : romdata_int = 'h8882;
    'hd7a : romdata_int = 'had55;
    'hd7b : romdata_int = 'hcc4f;
    'hd7c : romdata_int = 'hd200;
    'hd7d : romdata_int = 'hfa38;
    'hd7e : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd7f : romdata_int = 'h6a2;
    'hd80 : romdata_int = 'hc67;
    'hd81 : romdata_int = 'hcc4;
    'hd82 : romdata_int = 'h12d9;
    'hd83 : romdata_int = 'h2000;
    'hd84 : romdata_int = 'h4675;
    'hd85 : romdata_int = 'h7a00;
    'hd86 : romdata_int = 'ha8bd;
    'hd87 : romdata_int = 'haabc;
    'hd88 : romdata_int = 'hb657;
    'hd89 : romdata_int = 'hd400;
    'hd8a : romdata_int = 'he49e;
    'hd8b : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd8c : romdata_int = 'h550;
    'hd8d : romdata_int = 'h727;
    'hd8e : romdata_int = 'h73e;
    'hd8f : romdata_int = 'h2200;
    'hd90 : romdata_int = 'h38c0;
    'hd91 : romdata_int = 'h4eaa;
    'hd92 : romdata_int = 'h7c00;
    'hd93 : romdata_int = 'h8b4c;
    'hd94 : romdata_int = 'hb034;
    'hd95 : romdata_int = 'hccfb;
    'hd96 : romdata_int = 'hd600;
    'hd97 : romdata_int = 'h102e2;
    'hd98 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hd99 : romdata_int = 'hce4;
    'hd9a : romdata_int = 'hce6;
    'hd9b : romdata_int = 'hecb;
    'hd9c : romdata_int = 'h16f0;
    'hd9d : romdata_int = 'h1d41;
    'hd9e : romdata_int = 'h2400;
    'hd9f : romdata_int = 'h6538;
    'hda0 : romdata_int = 'h78d9;
    'hda1 : romdata_int = 'h7e00;
    'hda2 : romdata_int = 'hd800;
    'hda3 : romdata_int = 'hef34;
    'hda4 : romdata_int = 'hf2ff;
    'hda5 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hda6 : romdata_int = 'h2fc;
    'hda7 : romdata_int = 'h944;
    'hda8 : romdata_int = 'h182f;
    'hda9 : romdata_int = 'h1b5a;
    'hdaa : romdata_int = 'h2600;
    'hdab : romdata_int = 'h474e;
    'hdac : romdata_int = 'h8000;
    'hdad : romdata_int = 'h9b56;
    'hdae : romdata_int = 'haeb0;
    'hdaf : romdata_int = 'hc037;
    'hdb0 : romdata_int = 'hda00;
    'hdb1 : romdata_int = 'hfecf;
    'hdb2 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdb3 : romdata_int = 'hb35;
    'hdb4 : romdata_int = 'h1013;
    'hdb5 : romdata_int = 'h14f6;
    'hdb6 : romdata_int = 'h2800;
    'hdb7 : romdata_int = 'h36a6;
    'hdb8 : romdata_int = 'h4c87;
    'hdb9 : romdata_int = 'h5cdd;
    'hdba : romdata_int = 'h8200;
    'hdbb : romdata_int = 'h9467;
    'hdbc : romdata_int = 'hdc00;
    'hdbd : romdata_int = 'he226;
    'hdbe : romdata_int = 'h10941;
    'hdbf : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdc0 : romdata_int = 'h22c;
    'hdc1 : romdata_int = 'h48c;
    'hdc2 : romdata_int = 'h8a9;
    'hdc3 : romdata_int = 'h16f5;
    'hdc4 : romdata_int = 'h2099;
    'hdc5 : romdata_int = 'h2a00;
    'hdc6 : romdata_int = 'h70b4;
    'hdc7 : romdata_int = 'h8400;
    'hdc8 : romdata_int = 'ha46a;
    'hdc9 : romdata_int = 'hcf4b;
    'hdca : romdata_int = 'hdc62;
    'hdcb : romdata_int = 'hde00;
    'hdcc : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdcd : romdata_int = 'h3c;
    'hdce : romdata_int = 'h52e;
    'hdcf : romdata_int = 'h8fd;
    'hdd0 : romdata_int = 'h1085;
    'hdd1 : romdata_int = 'h12a2;
    'hdd2 : romdata_int = 'h2c00;
    'hdd3 : romdata_int = 'h8600;
    'hdd4 : romdata_int = 'ha2b7;
    'hdd5 : romdata_int = 'ha83e;
    'hdd6 : romdata_int = 'hc55c;
    'hdd7 : romdata_int = 'he000;
    'hdd8 : romdata_int = 'hf107;
    'hdd9 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdda : romdata_int = 'h74;
    'hddb : romdata_int = 'haa3;
    'hddc : romdata_int = 'hcae;
    'hddd : romdata_int = 'h2e00;
    'hdde : romdata_int = 'h2ec8;
    'hddf : romdata_int = 'h4818;
    'hde0 : romdata_int = 'h6f57;
    'hde1 : romdata_int = 'h80bb;
    'hde2 : romdata_int = 'h8800;
    'hde3 : romdata_int = 'hd457;
    'hde4 : romdata_int = 'hdb14;
    'hde5 : romdata_int = 'he200;
    'hde6 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hde7 : romdata_int = 'h129;
    'hde8 : romdata_int = 'h124b;
    'hde9 : romdata_int = 'h1748;
    'hdea : romdata_int = 'h3000;
    'hdeb : romdata_int = 'h3743;
    'hdec : romdata_int = 'h4cd6;
    'hded : romdata_int = 'h8a00;
    'hdee : romdata_int = 'h9cc2;
    'hdef : romdata_int = 'ha159;
    'hdf0 : romdata_int = 'he400;
    'hdf1 : romdata_int = 'hf923;
    'hdf2 : romdata_int = 'h10af7;
    'hdf3 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hdf4 : romdata_int = 'h108a;
    'hdf5 : romdata_int = 'h126a;
    'hdf6 : romdata_int = 'h1700;
    'hdf7 : romdata_int = 'h2d36;
    'hdf8 : romdata_int = 'h3200;
    'hdf9 : romdata_int = 'h552f;
    'hdfa : romdata_int = 'h8c00;
    'hdfb : romdata_int = 'h9f54;
    'hdfc : romdata_int = 'ha242;
    'hdfd : romdata_int = 'hb8aa;
    'hdfe : romdata_int = 'he600;
    'hdff : romdata_int = 'hed1c;
    'he00 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he01 : romdata_int = 'haf;
    'he02 : romdata_int = 'hf0f;
    'he03 : romdata_int = 'h1c43;
    'he04 : romdata_int = 'h1c91;
    'he05 : romdata_int = 'h32a1;
    'he06 : romdata_int = 'h3400;
    'he07 : romdata_int = 'h749d;
    'he08 : romdata_int = 'h8655;
    'he09 : romdata_int = 'h8e00;
    'he0a : romdata_int = 'he800;
    'he0b : romdata_int = 'hf0f8;
    'he0c : romdata_int = 'h10155;
    'he0d : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he0e : romdata_int = 'hcb1;
    'he0f : romdata_int = 'h113b;
    'he10 : romdata_int = 'h126d;
    'he11 : romdata_int = 'h2849;
    'he12 : romdata_int = 'h3600;
    'he13 : romdata_int = 'h4524;
    'he14 : romdata_int = 'h5eb6;
    'he15 : romdata_int = 'h9000;
    'he16 : romdata_int = 'h92a9;
    'he17 : romdata_int = 'hc2af;
    'he18 : romdata_int = 'hea00;
    'he19 : romdata_int = 'hec06;
    'he1a : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he1b : romdata_int = 'h149f;
    'he1c : romdata_int = 'h1cc2;
    'he1d : romdata_int = 'h1d5d;
    'he1e : romdata_int = 'h329e;
    'he1f : romdata_int = 'h3800;
    'he20 : romdata_int = 'h56be;
    'he21 : romdata_int = 'h8e5f;
    'he22 : romdata_int = 'h9200;
    'he23 : romdata_int = 'h9723;
    'he24 : romdata_int = 'he0bc;
    'he25 : romdata_int = 'hec00;
    'he26 : romdata_int = 'h10137;
    'he27 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he28 : romdata_int = 'h37;
    'he29 : romdata_int = 'ha7e;
    'he2a : romdata_int = 'h1602;
    'he2b : romdata_int = 'h1820;
    'he2c : romdata_int = 'h242c;
    'he2d : romdata_int = 'h3a00;
    'he2e : romdata_int = 'h6221;
    'he2f : romdata_int = 'h9400;
    'he30 : romdata_int = 'ha040;
    'he31 : romdata_int = 'hb91e;
    'he32 : romdata_int = 'hd0aa;
    'he33 : romdata_int = 'hee00;
    'he34 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he35 : romdata_int = 'h622;
    'he36 : romdata_int = 'hc4b;
    'he37 : romdata_int = 'hc84;
    'he38 : romdata_int = 'h14a5;
    'he39 : romdata_int = 'h2857;
    'he3a : romdata_int = 'h3c00;
    'he3b : romdata_int = 'h8339;
    'he3c : romdata_int = 'h8c7b;
    'he3d : romdata_int = 'h9600;
    'he3e : romdata_int = 'hb733;
    'he3f : romdata_int = 'hf000;
    'he40 : romdata_int = 'hfc8f;
    'he41 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he42 : romdata_int = 'h144;
    'he43 : romdata_int = 'h952;
    'he44 : romdata_int = 'he62;
    'he45 : romdata_int = 'h1a5d;
    'he46 : romdata_int = 'h3e00;
    'he47 : romdata_int = 'h583b;
    'he48 : romdata_int = 'h761f;
    'he49 : romdata_int = 'h8f18;
    'he4a : romdata_int = 'h9800;
    'he4b : romdata_int = 'hc6e7;
    'he4c : romdata_int = 'hf200;
    'he4d : romdata_int = 'h10d42;
    'he4e : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he4f : romdata_int = 'h2fd;
    'he50 : romdata_int = 'h4ae;
    'he51 : romdata_int = 'h654;
    'he52 : romdata_int = 'h104d;
    'he53 : romdata_int = 'h2328;
    'he54 : romdata_int = 'h4000;
    'he55 : romdata_int = 'h5a16;
    'he56 : romdata_int = 'h8c8c;
    'he57 : romdata_int = 'h9a00;
    'he58 : romdata_int = 'hee94;
    'he59 : romdata_int = 'hf400;
    'he5a : romdata_int = 'hfe98;
    'he5b : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he5c : romdata_int = 'h14e1;
    'he5d : romdata_int = 'h1cf8;
    'he5e : romdata_int = 'h1d4f;
    'he5f : romdata_int = 'h4200;
    'he60 : romdata_int = 'h4a2d;
    'he61 : romdata_int = 'h548a;
    'he62 : romdata_int = 'h690d;
    'he63 : romdata_int = 'h821c;
    'he64 : romdata_int = 'h9c00;
    'he65 : romdata_int = 'hbecc;
    'he66 : romdata_int = 'hf600;
    'he67 : romdata_int = 'h1046b;
    'he68 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he69 : romdata_int = 'h52a;
    'he6a : romdata_int = 'hea5;
    'he6b : romdata_int = 'h1960;
    'he6c : romdata_int = 'h4400;
    'he6d : romdata_int = 'h4436;
    'he6e : romdata_int = 'h4a17;
    'he6f : romdata_int = 'h745b;
    'he70 : romdata_int = 'h7afb;
    'he71 : romdata_int = 'h9e00;
    'he72 : romdata_int = 'hd322;
    'he73 : romdata_int = 'hda7f;
    'he74 : romdata_int = 'hf800;
    'he75 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he76 : romdata_int = 'h680;
    'he77 : romdata_int = 'ha23;
    'he78 : romdata_int = 'h1604;
    'he79 : romdata_int = 'h1d1d;
    'he7a : romdata_int = 'h352f;
    'he7b : romdata_int = 'h4600;
    'he7c : romdata_int = 'h6a8f;
    'he7d : romdata_int = 'ha000;
    'he7e : romdata_int = 'hacad;
    'he7f : romdata_int = 'he133;
    'he80 : romdata_int = 'hf566;
    'he81 : romdata_int = 'hfa00;
    'he82 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he83 : romdata_int = 'h6ae;
    'he84 : romdata_int = 'hb60;
    'he85 : romdata_int = 'hd54;
    'he86 : romdata_int = 'h1ab8;
    'he87 : romdata_int = 'h3836;
    'he88 : romdata_int = 'h4800;
    'he89 : romdata_int = 'h8533;
    'he8a : romdata_int = 'h9ea4;
    'he8b : romdata_int = 'ha200;
    'he8c : romdata_int = 'hea08;
    'he8d : romdata_int = 'hf942;
    'he8e : romdata_int = 'hfc00;
    'he8f : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he90 : romdata_int = 'h31b;
    'he91 : romdata_int = 'h1247;
    'he92 : romdata_int = 'h183b;
    'he93 : romdata_int = 'h1ab0;
    'he94 : romdata_int = 'h1c6b;
    'he95 : romdata_int = 'h4a00;
    'he96 : romdata_int = 'h6d4b;
    'he97 : romdata_int = 'h9936;
    'he98 : romdata_int = 'ha400;
    'he99 : romdata_int = 'hcafb;
    'he9a : romdata_int = 'hfe00;
    'he9b : romdata_int = 'h10a72;
    'he9c : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'he9d : romdata_int = 'hf19;
    'he9e : romdata_int = 'h140a;
    'he9f : romdata_int = 'h1d2f;
    'hea0 : romdata_int = 'h2a8a;
    'hea1 : romdata_int = 'h42f3;
    'hea2 : romdata_int = 'h4c00;
    'hea3 : romdata_int = 'h8040;
    'hea4 : romdata_int = 'ha600;
    'hea5 : romdata_int = 'hb0c0;
    'hea6 : romdata_int = 'hfaf9;
    'hea7 : romdata_int = 'h10000;
    'hea8 : romdata_int = 'h10509;
    'hea9 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'heaa : romdata_int = 'ha3;
    'heab : romdata_int = 'he2e;
    'heac : romdata_int = 'h1523;
    'head : romdata_int = 'h265f;
    'heae : romdata_int = 'h4085;
    'heaf : romdata_int = 'h4e00;
    'heb0 : romdata_int = 'h6207;
    'heb1 : romdata_int = 'ha66b;
    'heb2 : romdata_int = 'ha800;
    'heb3 : romdata_int = 'hcacd;
    'heb4 : romdata_int = 'hde1d;
    'heb5 : romdata_int = 'h10200;
    'heb6 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'heb7 : romdata_int = 'h8d;
    'heb8 : romdata_int = 'hf8;
    'heb9 : romdata_int = 'h16eb;
    'heba : romdata_int = 'h189e;
    'hebb : romdata_int = 'h1a54;
    'hebc : romdata_int = 'h5000;
    'hebd : romdata_int = 'h7a8b;
    'hebe : romdata_int = 'h8658;
    'hebf : romdata_int = 'haa00;
    'hec0 : romdata_int = 'hce3a;
    'hec1 : romdata_int = 'hf33f;
    'hec2 : romdata_int = 'h10400;
    'hec3 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hec4 : romdata_int = 'had1;
    'hec5 : romdata_int = 'h10ba;
    'hec6 : romdata_int = 'h16b0;
    'hec7 : romdata_int = 'h1a11;
    'hec8 : romdata_int = 'h5200;
    'hec9 : romdata_int = 'h5904;
    'heca : romdata_int = 'h910f;
    'hecb : romdata_int = 'ha6f6;
    'hecc : romdata_int = 'hac00;
    'hecd : romdata_int = 'hbe82;
    'hece : romdata_int = 'h10600;
    'hecf : romdata_int = 'h108b2;
    'hed0 : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hed1 : romdata_int = 'h207;
    'hed2 : romdata_int = 'h212;
    'hed3 : romdata_int = 'h6c2;
    'hed4 : romdata_int = 'h3041;
    'hed5 : romdata_int = 'h313a;
    'hed6 : romdata_int = 'h5400;
    'hed7 : romdata_int = 'h6d19;
    'hed8 : romdata_int = 'h7ec9;
    'hed9 : romdata_int = 'hae00;
    'heda : romdata_int = 'hbab5;
    'hedb : romdata_int = 'hea6d;
    'hedc : romdata_int = 'h10800;
    'hedd : romdata_int = 'h4b2d; // Line descriptor for 3_4
    'hede : romdata_int = 'h23b;
    'hedf : romdata_int = 'h425;
    'hee0 : romdata_int = 'h82e;
    'hee1 : romdata_int = 'h16a7;
    'hee2 : romdata_int = 'h5265;
    'hee3 : romdata_int = 'h5600;
    'hee4 : romdata_int = 'h9102;
    'hee5 : romdata_int = 'h9539;
    'hee6 : romdata_int = 'hb000;
    'hee7 : romdata_int = 'he6c4;
    'hee8 : romdata_int = 'he74c;
    'hee9 : romdata_int = 'h10a00;
    'heea : romdata_int = 'h6b2d; // Line descriptor for 3_4
    'heeb : romdata_int = 'h2a0;
    'heec : romdata_int = 'he0d;
    'heed : romdata_int = 'h1871;
    'heee : romdata_int = 'h1e45;
    'heef : romdata_int = 'h56ae;
    'hef0 : romdata_int = 'h5800;
    'hef1 : romdata_int = 'h78a8;
    'hef2 : romdata_int = 'h96d4;
    'hef3 : romdata_int = 'hb200;
    'hef4 : romdata_int = 'hba26;
    'hef5 : romdata_int = 'h10687;
    'hef6 : romdata_int = 'h10c00;
    'hef7 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hef8 : romdata_int = 'h0;
    'hef9 : romdata_int = 'hc68;
    'hefa : romdata_int = 'h1945;
    'hefb : romdata_int = 'h1eb5;
    'hefc : romdata_int = 'h1f3f;
    'hefd : romdata_int = 'h22f3;
    'hefe : romdata_int = 'h3279;
    'heff : romdata_int = 'h4800;
    'hf00 : romdata_int = 'h4e3d;
    'hf01 : romdata_int = 'h6248;
    'hf02 : romdata_int = 'h9000;
    'hf03 : romdata_int = 'ha222;
    'hf04 : romdata_int = 'hacc8;
    'hf05 : romdata_int = 'hd800;
    'hf06 : romdata_int = 'hfae7;
    'hf07 : romdata_int = 'h11702;
    'hf08 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf09 : romdata_int = 'h200;
    'hf0a : romdata_int = 'h1207;
    'hf0b : romdata_int = 'h14f2;
    'hf0c : romdata_int = 'h1c60;
    'hf0d : romdata_int = 'h233b;
    'hf0e : romdata_int = 'h374a;
    'hf0f : romdata_int = 'h4321;
    'hf10 : romdata_int = 'h4a00;
    'hf11 : romdata_int = 'h5329;
    'hf12 : romdata_int = 'h7e61;
    'hf13 : romdata_int = 'h9200;
    'hf14 : romdata_int = 'hc017;
    'hf15 : romdata_int = 'hc567;
    'hf16 : romdata_int = 'hda00;
    'hf17 : romdata_int = 'hed58;
    'hf18 : romdata_int = 'hf2d3;
    'hf19 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf1a : romdata_int = 'h400;
    'hf1b : romdata_int = 'ha5f;
    'hf1c : romdata_int = 'he1f;
    'hf1d : romdata_int = 'h14da;
    'hf1e : romdata_int = 'h186b;
    'hf1f : romdata_int = 'h261c;
    'hf20 : romdata_int = 'h2b55;
    'hf21 : romdata_int = 'h4c00;
    'hf22 : romdata_int = 'h614c;
    'hf23 : romdata_int = 'h863a;
    'hf24 : romdata_int = 'h9400;
    'hf25 : romdata_int = 'h9c9c;
    'hf26 : romdata_int = 'hd4e2;
    'hf27 : romdata_int = 'hdc00;
    'hf28 : romdata_int = 'hed4d;
    'hf29 : romdata_int = 'hfab7;
    'hf2a : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf2b : romdata_int = 'h600;
    'hf2c : romdata_int = 'ha1c;
    'hf2d : romdata_int = 'ha3b;
    'hf2e : romdata_int = 'h1241;
    'hf2f : romdata_int = 'h16fe;
    'hf30 : romdata_int = 'h1e4c;
    'hf31 : romdata_int = 'h251a;
    'hf32 : romdata_int = 'h4e00;
    'hf33 : romdata_int = 'h50d1;
    'hf34 : romdata_int = 'h74d8;
    'hf35 : romdata_int = 'h9089;
    'hf36 : romdata_int = 'h9600;
    'hf37 : romdata_int = 'hbcb8;
    'hf38 : romdata_int = 'hde00;
    'hf39 : romdata_int = 'h10007;
    'hf3a : romdata_int = 'h102a2;
    'hf3b : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf3c : romdata_int = 'h800;
    'hf3d : romdata_int = 'h94d;
    'hf3e : romdata_int = 'hc1a;
    'hf3f : romdata_int = 'heb4;
    'hf40 : romdata_int = 'h1eb8;
    'hf41 : romdata_int = 'h3c3e;
    'hf42 : romdata_int = 'h3eb0;
    'hf43 : romdata_int = 'h5000;
    'hf44 : romdata_int = 'h62ce;
    'hf45 : romdata_int = 'h6ca7;
    'hf46 : romdata_int = 'h9800;
    'hf47 : romdata_int = 'ha85a;
    'hf48 : romdata_int = 'hd011;
    'hf49 : romdata_int = 'he000;
    'hf4a : romdata_int = 'hf403;
    'hf4b : romdata_int = 'h10d0e;
    'hf4c : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf4d : romdata_int = 'h4;
    'hf4e : romdata_int = 'ha00;
    'hf4f : romdata_int = 'ha71;
    'hf50 : romdata_int = 'h127d;
    'hf51 : romdata_int = 'h1b3e;
    'hf52 : romdata_int = 'h20e5;
    'hf53 : romdata_int = 'h2c7a;
    'hf54 : romdata_int = 'h5200;
    'hf55 : romdata_int = 'h58df;
    'hf56 : romdata_int = 'h6613;
    'hf57 : romdata_int = 'h9a00;
    'hf58 : romdata_int = 'hc23d;
    'hf59 : romdata_int = 'hd30f;
    'hf5a : romdata_int = 'he200;
    'hf5b : romdata_int = 'h10003;
    'hf5c : romdata_int = 'h102ac;
    'hf5d : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf5e : romdata_int = 'hc00;
    'hf5f : romdata_int = 'heda;
    'hf60 : romdata_int = 'h10ea;
    'hf61 : romdata_int = 'h163f;
    'hf62 : romdata_int = 'h16a8;
    'hf63 : romdata_int = 'h1a45;
    'hf64 : romdata_int = 'h3646;
    'hf65 : romdata_int = 'h5400;
    'hf66 : romdata_int = 'h544b;
    'hf67 : romdata_int = 'h726f;
    'hf68 : romdata_int = 'h9c00;
    'hf69 : romdata_int = 'hb03d;
    'hf6a : romdata_int = 'hb156;
    'hf6b : romdata_int = 'he400;
    'hf6c : romdata_int = 'h10898;
    'hf6d : romdata_int = 'h10f40;
    'hf6e : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf6f : romdata_int = 'h94f;
    'hf70 : romdata_int = 'hc4e;
    'hf71 : romdata_int = 'he00;
    'hf72 : romdata_int = 'h14bc;
    'hf73 : romdata_int = 'h14e3;
    'hf74 : romdata_int = 'h1caf;
    'hf75 : romdata_int = 'h2723;
    'hf76 : romdata_int = 'h5600;
    'hf77 : romdata_int = 'h5a7b;
    'hf78 : romdata_int = 'h7e44;
    'hf79 : romdata_int = 'h9275;
    'hf7a : romdata_int = 'h9e00;
    'hf7b : romdata_int = 'hac5b;
    'hf7c : romdata_int = 'he600;
    'hf7d : romdata_int = 'he8ce;
    'hf7e : romdata_int = 'h11108;
    'hf7f : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf80 : romdata_int = 'he1;
    'hf81 : romdata_int = 'h1000;
    'hf82 : romdata_int = 'h1106;
    'hf83 : romdata_int = 'h122b;
    'hf84 : romdata_int = 'h14f8;
    'hf85 : romdata_int = 'h1c69;
    'hf86 : romdata_int = 'h28f7;
    'hf87 : romdata_int = 'h5800;
    'hf88 : romdata_int = 'h6824;
    'hf89 : romdata_int = 'h8cec;
    'hf8a : romdata_int = 'h9af9;
    'hf8b : romdata_int = 'ha000;
    'hf8c : romdata_int = 'hc8a5;
    'hf8d : romdata_int = 'he060;
    'hf8e : romdata_int = 'he800;
    'hf8f : romdata_int = 'h10a3b;
    'hf90 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hf91 : romdata_int = 'hec;
    'hf92 : romdata_int = 'h31e;
    'hf93 : romdata_int = 'h49a;
    'hf94 : romdata_int = 'h523;
    'hf95 : romdata_int = 'h1200;
    'hf96 : romdata_int = 'h1aa2;
    'hf97 : romdata_int = 'h34c6;
    'hf98 : romdata_int = 'h490b;
    'hf99 : romdata_int = 'h5a00;
    'hf9a : romdata_int = 'h786e;
    'hf9b : romdata_int = 'ha200;
    'hf9c : romdata_int = 'hc6f3;
    'hf9d : romdata_int = 'hd520;
    'hf9e : romdata_int = 'hea00;
    'hf9f : romdata_int = 'hf6dd;
    'hfa0 : romdata_int = 'h11e9a;
    'hfa1 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfa2 : romdata_int = 'h65a;
    'hfa3 : romdata_int = 'h8ab;
    'hfa4 : romdata_int = 'h1400;
    'hfa5 : romdata_int = 'h183c;
    'hfa6 : romdata_int = 'h186e;
    'hfa7 : romdata_int = 'h1b4c;
    'hfa8 : romdata_int = 'h3308;
    'hfa9 : romdata_int = 'h5c00;
    'hfaa : romdata_int = 'h5eb6;
    'hfab : romdata_int = 'h82b7;
    'hfac : romdata_int = 'ha2f6;
    'hfad : romdata_int = 'ha400;
    'hfae : romdata_int = 'hb91e;
    'hfaf : romdata_int = 'hec00;
    'hfb0 : romdata_int = 'hf11a;
    'hfb1 : romdata_int = 'hf428;
    'hfb2 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfb3 : romdata_int = 'h1072;
    'hfb4 : romdata_int = 'h10ee;
    'hfb5 : romdata_int = 'h1600;
    'hfb6 : romdata_int = 'h1966;
    'hfb7 : romdata_int = 'h1e0f;
    'hfb8 : romdata_int = 'h1f50;
    'hfb9 : romdata_int = 'h4344;
    'hfba : romdata_int = 'h5e00;
    'hfbb : romdata_int = 'h707b;
    'hfbc : romdata_int = 'h833f;
    'hfbd : romdata_int = 'h9697;
    'hfbe : romdata_int = 'ha600;
    'hfbf : romdata_int = 'hb50a;
    'hfc0 : romdata_int = 'hee00;
    'hfc1 : romdata_int = 'hfcfa;
    'hfc2 : romdata_int = 'h11156;
    'hfc3 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfc4 : romdata_int = 'hb;
    'hfc5 : romdata_int = 'h164;
    'hfc6 : romdata_int = 'h44e;
    'hfc7 : romdata_int = 'h142f;
    'hfc8 : romdata_int = 'h16f5;
    'hfc9 : romdata_int = 'h1800;
    'hfca : romdata_int = 'h3cf2;
    'hfcb : romdata_int = 'h5d00;
    'hfcc : romdata_int = 'h6000;
    'hfcd : romdata_int = 'h7a79;
    'hfce : romdata_int = 'ha0f6;
    'hfcf : romdata_int = 'ha800;
    'hfd0 : romdata_int = 'haaa2;
    'hfd1 : romdata_int = 'he2c1;
    'hfd2 : romdata_int = 'hf000;
    'hfd3 : romdata_int = 'h10c26;
    'hfd4 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfd5 : romdata_int = 'h60e;
    'hfd6 : romdata_int = 'h88f;
    'hfd7 : romdata_int = 'he7e;
    'hfd8 : romdata_int = 'h129d;
    'hfd9 : romdata_int = 'h1a00;
    'hfda : romdata_int = 'h2032;
    'hfdb : romdata_int = 'h3b2f;
    'hfdc : romdata_int = 'h6200;
    'hfdd : romdata_int = 'h870b;
    'hfde : romdata_int = 'h8c33;
    'hfdf : romdata_int = 'h9859;
    'hfe0 : romdata_int = 'ha67a;
    'hfe1 : romdata_int = 'haa00;
    'hfe2 : romdata_int = 'hd8ca;
    'hfe3 : romdata_int = 'hf200;
    'hfe4 : romdata_int = 'h10661;
    'hfe5 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hfe6 : romdata_int = 'he23;
    'hfe7 : romdata_int = 'h174b;
    'hfe8 : romdata_int = 'h1c00;
    'hfe9 : romdata_int = 'h1ee2;
    'hfea : romdata_int = 'h223a;
    'hfeb : romdata_int = 'h2cc4;
    'hfec : romdata_int = 'h40ee;
    'hfed : romdata_int = 'h6400;
    'hfee : romdata_int = 'h7c94;
    'hfef : romdata_int = 'h8a63;
    'hff0 : romdata_int = 'ha607;
    'hff1 : romdata_int = 'hac00;
    'hff2 : romdata_int = 'haf39;
    'hff3 : romdata_int = 'hf400;
    'hff4 : romdata_int = 'hff05;
    'hff5 : romdata_int = 'h10566;
    'hff6 : romdata_int = 'h4f24; // Line descriptor for 4_5
    'hff7 : romdata_int = 'h683;
    'hff8 : romdata_int = 'hac5;
    'hff9 : romdata_int = 'he70;
    'hffa : romdata_int = 'hf46;
    'hffb : romdata_int = 'h16fc;
    'hffc : romdata_int = 'h18cb;
    'hffd : romdata_int = 'h1e00;
    'hffe : romdata_int = 'h6600;
    'hfff : romdata_int = 'h7309;
    'h1000: romdata_int = 'h8883;
    'h1001: romdata_int = 'hae00;
    'h1002: romdata_int = 'hc63b;
    'h1003: romdata_int = 'hd6a1;
    'h1004: romdata_int = 'hdee7;
    'h1005: romdata_int = 'hf225;
    'h1006: romdata_int = 'hf600;
    'h1007: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1008: romdata_int = 'h137;
    'h1009: romdata_int = 'ha67;
    'h100a: romdata_int = 'hd2c;
    'h100b: romdata_int = 'h1745;
    'h100c: romdata_int = 'h1e47;
    'h100d: romdata_int = 'h2000;
    'h100e: romdata_int = 'h22ba;
    'h100f: romdata_int = 'h6800;
    'h1010: romdata_int = 'h7caf;
    'h1011: romdata_int = 'h8a48;
    'h1012: romdata_int = 'h9d5a;
    'h1013: romdata_int = 'hb000;
    'h1014: romdata_int = 'hc94d;
    'h1015: romdata_int = 'hf800;
    'h1016: romdata_int = 'h11a07;
    'h1017: romdata_int = 'h11ec5;
    'h1018: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1019: romdata_int = 'h26b;
    'h101a: romdata_int = 'h261;
    'h101b: romdata_int = 'h291;
    'h101c: romdata_int = 'hd41;
    'h101d: romdata_int = 'h100b;
    'h101e: romdata_int = 'h2200;
    'h101f: romdata_int = 'h2298;
    'h1020: romdata_int = 'h5c73;
    'h1021: romdata_int = 'h6a00;
    'h1022: romdata_int = 'h8840;
    'h1023: romdata_int = 'h9e28;
    'h1024: romdata_int = 'hb200;
    'h1025: romdata_int = 'hc10d;
    'h1026: romdata_int = 'hf8cd;
    'h1027: romdata_int = 'hf8f8;
    'h1028: romdata_int = 'hfa00;
    'h1029: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h102a: romdata_int = 'h116;
    'h102b: romdata_int = 'h1158;
    'h102c: romdata_int = 'h12fd;
    'h102d: romdata_int = 'h18e5;
    'h102e: romdata_int = 'h20b5;
    'h102f: romdata_int = 'h2400;
    'h1030: romdata_int = 'h4658;
    'h1031: romdata_int = 'h6b4b;
    'h1032: romdata_int = 'h6c00;
    'h1033: romdata_int = 'h7629;
    'h1034: romdata_int = 'hb400;
    'h1035: romdata_int = 'hbb33;
    'h1036: romdata_int = 'hd0c6;
    'h1037: romdata_int = 'hf6eb;
    'h1038: romdata_int = 'hfc00;
    'h1039: romdata_int = 'hfeab;
    'h103a: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h103b: romdata_int = 'h4d8;
    'h103c: romdata_int = 'h825;
    'h103d: romdata_int = 'ha9f;
    'h103e: romdata_int = 'h1697;
    'h103f: romdata_int = 'h2080;
    'h1040: romdata_int = 'h2600;
    'h1041: romdata_int = 'h2b1c;
    'h1042: romdata_int = 'h4c87;
    'h1043: romdata_int = 'h6d09;
    'h1044: romdata_int = 'h6e00;
    'h1045: romdata_int = 'ha4e8;
    'h1046: romdata_int = 'hb600;
    'h1047: romdata_int = 'hc232;
    'h1048: romdata_int = 'hdcfa;
    'h1049: romdata_int = 'hef0e;
    'h104a: romdata_int = 'hfe00;
    'h104b: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h104c: romdata_int = 'h452;
    'h104d: romdata_int = 'h550;
    'h104e: romdata_int = 'h677;
    'h104f: romdata_int = 'h1cdd;
    'h1050: romdata_int = 'h2251;
    'h1051: romdata_int = 'h2800;
    'h1052: romdata_int = 'h3a54;
    'h1053: romdata_int = 'h4e09;
    'h1054: romdata_int = 'h6819;
    'h1055: romdata_int = 'h7000;
    'h1056: romdata_int = 'h9e23;
    'h1057: romdata_int = 'hb800;
    'h1058: romdata_int = 'hd6d3;
    'h1059: romdata_int = 'heae1;
    'h105a: romdata_int = 'h10000;
    'h105b: romdata_int = 'h11655;
    'h105c: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h105d: romdata_int = 'h328;
    'h105e: romdata_int = 'h1b37;
    'h105f: romdata_int = 'h1ca6;
    'h1060: romdata_int = 'h1cd6;
    'h1061: romdata_int = 'h2359;
    'h1062: romdata_int = 'h2a00;
    'h1063: romdata_int = 'h351d;
    'h1064: romdata_int = 'h7074;
    'h1065: romdata_int = 'h7200;
    'h1066: romdata_int = 'h792a;
    'h1067: romdata_int = 'h9a12;
    'h1068: romdata_int = 'hb94e;
    'h1069: romdata_int = 'hba00;
    'h106a: romdata_int = 'he89b;
    'h106b: romdata_int = 'h10200;
    'h106c: romdata_int = 'h10679;
    'h106d: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h106e: romdata_int = 'h20d;
    'h106f: romdata_int = 'hd08;
    'h1070: romdata_int = 'hd3f;
    'h1071: romdata_int = 'h20a8;
    'h1072: romdata_int = 'h2067;
    'h1073: romdata_int = 'h2149;
    'h1074: romdata_int = 'h2c00;
    'h1075: romdata_int = 'h56a6;
    'h1076: romdata_int = 'h5a86;
    'h1077: romdata_int = 'h7400;
    'h1078: romdata_int = 'h96c1;
    'h1079: romdata_int = 'h989c;
    'h107a: romdata_int = 'hbc00;
    'h107b: romdata_int = 'hde7a;
    'h107c: romdata_int = 'h10400;
    'h107d: romdata_int = 'h114fa;
    'h107e: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h107f: romdata_int = 'h841;
    'h1080: romdata_int = 'h952;
    'h1081: romdata_int = 'hf3f;
    'h1082: romdata_int = 'he90;
    'h1083: romdata_int = 'hf63;
    'h1084: romdata_int = 'h2e00;
    'h1085: romdata_int = 'h44b3;
    'h1086: romdata_int = 'h54bb;
    'h1087: romdata_int = 'h7600;
    'h1088: romdata_int = 'h7a60;
    'h1089: romdata_int = 'hb27d;
    'h108a: romdata_int = 'hbe00;
    'h108b: romdata_int = 'hca58;
    'h108c: romdata_int = 'he238;
    'h108d: romdata_int = 'h10600;
    'h108e: romdata_int = 'h112e4;
    'h108f: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1090: romdata_int = 'hb0;
    'h1091: romdata_int = 'h40f;
    'h1092: romdata_int = 'habd;
    'h1093: romdata_int = 'hb32;
    'h1094: romdata_int = 'h1678;
    'h1095: romdata_int = 'h1f11;
    'h1096: romdata_int = 'h3000;
    'h1097: romdata_int = 'h650b;
    'h1098: romdata_int = 'h6e08;
    'h1099: romdata_int = 'h7800;
    'h109a: romdata_int = 'h9530;
    'h109b: romdata_int = 'hc000;
    'h109c: romdata_int = 'hcec5;
    'h109d: romdata_int = 'hdad7;
    'h109e: romdata_int = 'h10800;
    'h109f: romdata_int = 'h11230;
    'h10a0: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10a1: romdata_int = 'h718;
    'h10a2: romdata_int = 'h1a16;
    'h10a3: romdata_int = 'h1c7d;
    'h10a4: romdata_int = 'h22d9;
    'h10a5: romdata_int = 'h234c;
    'h10a6: romdata_int = 'h3200;
    'h10a7: romdata_int = 'h3836;
    'h10a8: romdata_int = 'h7a00;
    'h10a9: romdata_int = 'h80cd;
    'h10aa: romdata_int = 'h8151;
    'h10ab: romdata_int = 'hbf12;
    'h10ac: romdata_int = 'hc200;
    'h10ad: romdata_int = 'hcd2f;
    'h10ae: romdata_int = 'hea87;
    'h10af: romdata_int = 'h10a00;
    'h10b0: romdata_int = 'h10a7b;
    'h10b1: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10b2: romdata_int = 'h267;
    'h10b3: romdata_int = 'hc28;
    'h10b4: romdata_int = 'h1273;
    'h10b5: romdata_int = 'h14e4;
    'h10b6: romdata_int = 'h1a7a;
    'h10b7: romdata_int = 'h291c;
    'h10b8: romdata_int = 'h3400;
    'h10b9: romdata_int = 'h50b8;
    'h10ba: romdata_int = 'h64f4;
    'h10bb: romdata_int = 'h7c00;
    'h10bc: romdata_int = 'h94df;
    'h10bd: romdata_int = 'hae29;
    'h10be: romdata_int = 'hc400;
    'h10bf: romdata_int = 'he613;
    'h10c0: romdata_int = 'hef16;
    'h10c1: romdata_int = 'h10c00;
    'h10c2: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10c3: romdata_int = 'hd38;
    'h10c4: romdata_int = 'h107b;
    'h10c5: romdata_int = 'h1282;
    'h10c6: romdata_int = 'h14f6;
    'h10c7: romdata_int = 'h1a28;
    'h10c8: romdata_int = 'h1e6f;
    'h10c9: romdata_int = 'h3600;
    'h10ca: romdata_int = 'h5932;
    'h10cb: romdata_int = 'h7e00;
    'h10cc: romdata_int = 'h847b;
    'h10cd: romdata_int = 'haaa7;
    'h10ce: romdata_int = 'hb4c2;
    'h10cf: romdata_int = 'hc600;
    'h10d0: romdata_int = 'h10e00;
    'h10d1: romdata_int = 'h118d0;
    'h10d2: romdata_int = 'h11c6f;
    'h10d3: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10d4: romdata_int = 'h613;
    'h10d5: romdata_int = 'h6d0;
    'h10d6: romdata_int = 'hb2a;
    'h10d7: romdata_int = 'hc21;
    'h10d8: romdata_int = 'h22d4;
    'h10d9: romdata_int = 'h314c;
    'h10da: romdata_int = 'h3800;
    'h10db: romdata_int = 'h5243;
    'h10dc: romdata_int = 'h7553;
    'h10dd: romdata_int = 'h8000;
    'h10de: romdata_int = 'hba8d;
    'h10df: romdata_int = 'hc800;
    'h10e0: romdata_int = 'hcaf1;
    'h10e1: romdata_int = 'hf00b;
    'h10e2: romdata_int = 'h1046a;
    'h10e3: romdata_int = 'h11000;
    'h10e4: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10e5: romdata_int = 'h4c4;
    'h10e6: romdata_int = 'h1907;
    'h10e7: romdata_int = 'h1a0e;
    'h10e8: romdata_int = 'h1c2a;
    'h10e9: romdata_int = 'h20db;
    'h10ea: romdata_int = 'h393e;
    'h10eb: romdata_int = 'h3a00;
    'h10ec: romdata_int = 'h6a22;
    'h10ed: romdata_int = 'h6ed2;
    'h10ee: romdata_int = 'h8200;
    'h10ef: romdata_int = 'hb21a;
    'h10f0: romdata_int = 'hc4b9;
    'h10f1: romdata_int = 'hca00;
    'h10f2: romdata_int = 'h11200;
    'h10f3: romdata_int = 'h1140d;
    'h10f4: romdata_int = 'h11d56;
    'h10f5: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h10f6: romdata_int = 'h28a;
    'h10f7: romdata_int = 'h4f2;
    'h10f8: romdata_int = 'h103e;
    'h10f9: romdata_int = 'h1c52;
    'h10fa: romdata_int = 'h2155;
    'h10fb: romdata_int = 'h3c00;
    'h10fc: romdata_int = 'h4752;
    'h10fd: romdata_int = 'h5f54;
    'h10fe: romdata_int = 'h6696;
    'h10ff: romdata_int = 'h8400;
    'h1100: romdata_int = 'hbcbf;
    'h1101: romdata_int = 'hcc00;
    'h1102: romdata_int = 'hd28e;
    'h1103: romdata_int = 'he011;
    'h1104: romdata_int = 'he415;
    'h1105: romdata_int = 'h11400;
    'h1106: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1107: romdata_int = 'h9a;
    'h1108: romdata_int = 'h15c;
    'h1109: romdata_int = 'h10db;
    'h110a: romdata_int = 'h1a91;
    'h110b: romdata_int = 'h2f54;
    'h110c: romdata_int = 'h3e00;
    'h110d: romdata_int = 'h4562;
    'h110e: romdata_int = 'h4a9b;
    'h110f: romdata_int = 'h8600;
    'h1110: romdata_int = 'h8e6f;
    'h1111: romdata_int = 'h909c;
    'h1112: romdata_int = 'ha06b;
    'h1113: romdata_int = 'hce00;
    'h1114: romdata_int = 'hdb2d;
    'h1115: romdata_int = 'hdd56;
    'h1116: romdata_int = 'h11600;
    'h1117: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1118: romdata_int = 'h255;
    'h1119: romdata_int = 'h10c3;
    'h111a: romdata_int = 'h1738;
    'h111b: romdata_int = 'h1d08;
    'h111c: romdata_int = 'h30bd;
    'h111d: romdata_int = 'h3efc;
    'h111e: romdata_int = 'h4000;
    'h111f: romdata_int = 'h568e;
    'h1120: romdata_int = 'h60d2;
    'h1121: romdata_int = 'h8800;
    'h1122: romdata_int = 'ha4a5;
    'h1123: romdata_int = 'hb646;
    'h1124: romdata_int = 'hd000;
    'h1125: romdata_int = 'h108f0;
    'h1126: romdata_int = 'h11800;
    'h1127: romdata_int = 'h11a4a;
    'h1128: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h1129: romdata_int = 'h43b;
    'h112a: romdata_int = 'h64e;
    'h112b: romdata_int = 'h80e;
    'h112c: romdata_int = 'h126b;
    'h112d: romdata_int = 'h191e;
    'h112e: romdata_int = 'h2030;
    'h112f: romdata_int = 'h4200;
    'h1130: romdata_int = 'h493d;
    'h1131: romdata_int = 'h8547;
    'h1132: romdata_int = 'h8a00;
    'h1133: romdata_int = 'hbe3a;
    'h1134: romdata_int = 'hceae;
    'h1135: romdata_int = 'hd200;
    'h1136: romdata_int = 'he453;
    'h1137: romdata_int = 'h11844;
    'h1138: romdata_int = 'h11a00;
    'h1139: romdata_int = 'h4f24; // Line descriptor for 4_5
    'h113a: romdata_int = 'h6e7;
    'h113b: romdata_int = 'h875;
    'h113c: romdata_int = 'h1267;
    'h113d: romdata_int = 'h14dc;
    'h113e: romdata_int = 'h2474;
    'h113f: romdata_int = 'h40cb;
    'h1140: romdata_int = 'h4400;
    'h1141: romdata_int = 'h4acf;
    'h1142: romdata_int = 'h76f3;
    'h1143: romdata_int = 'h8c00;
    'h1144: romdata_int = 'h9233;
    'h1145: romdata_int = 'ha866;
    'h1146: romdata_int = 'hd400;
    'h1147: romdata_int = 'he639;
    'h1148: romdata_int = 'hfcbd;
    'h1149: romdata_int = 'h11c00;
    'h114a: romdata_int = 'h6f24; // Line descriptor for 4_5
    'h114b: romdata_int = 'h2d5;
    'h114c: romdata_int = 'h64a;
    'h114d: romdata_int = 'h938;
    'h114e: romdata_int = 'h14ef;
    'h114f: romdata_int = 'h1839;
    'h1150: romdata_int = 'h2e6b;
    'h1151: romdata_int = 'h4600;
    'h1152: romdata_int = 'h4c77;
    'h1153: romdata_int = 'h8e00;
    'h1154: romdata_int = 'h8e1f;
    'h1155: romdata_int = 'hb638;
    'h1156: romdata_int = 'hcce2;
    'h1157: romdata_int = 'hd600;
    'h1158: romdata_int = 'hd911;
    'h1159: romdata_int = 'h10f50;
    'h115a: romdata_int = 'h11e00;
    'h115b: romdata_int = 'h531e; // Line descriptor for 5_6
    'h115c: romdata_int = 'h0;
    'h115d: romdata_int = 'h738;
    'h115e: romdata_int = 'hd4c;
    'h115f: romdata_int = 'h1056;
    'h1160: romdata_int = 'h1280;
    'h1161: romdata_int = 'h1a8e;
    'h1162: romdata_int = 'h1c13;
    'h1163: romdata_int = 'h1c78;
    'h1164: romdata_int = 'h3c00;
    'h1165: romdata_int = 'h5058;
    'h1166: romdata_int = 'h6d18;
    'h1167: romdata_int = 'h7800;
    'h1168: romdata_int = 'h9118;
    'h1169: romdata_int = 'h9c15;
    'h116a: romdata_int = 'hb400;
    'h116b: romdata_int = 'hc26c;
    'h116c: romdata_int = 'heca1;
    'h116d: romdata_int = 'hf000;
    'h116e: romdata_int = 'h1106f;
    'h116f: romdata_int = 'h11897;
    'h1170: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1171: romdata_int = 'h200;
    'h1172: romdata_int = 'h2c9;
    'h1173: romdata_int = 'h467;
    'h1174: romdata_int = 'h4bd;
    'h1175: romdata_int = 'hf07;
    'h1176: romdata_int = 'h1adf;
    'h1177: romdata_int = 'h1efe;
    'h1178: romdata_int = 'h271c;
    'h1179: romdata_int = 'h3e00;
    'h117a: romdata_int = 'h3e58;
    'h117b: romdata_int = 'h5d11;
    'h117c: romdata_int = 'h7a00;
    'h117d: romdata_int = 'h86ab;
    'h117e: romdata_int = 'h8ad3;
    'h117f: romdata_int = 'hb600;
    'h1180: romdata_int = 'hc8bf;
    'h1181: romdata_int = 'hcacc;
    'h1182: romdata_int = 'hf200;
    'h1183: romdata_int = 'h1062b;
    'h1184: romdata_int = 'h12847;
    'h1185: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1186: romdata_int = 'h61;
    'h1187: romdata_int = 'h400;
    'h1188: romdata_int = 'ha87;
    'h1189: romdata_int = 'h12db;
    'h118a: romdata_int = 'h18f5;
    'h118b: romdata_int = 'h193e;
    'h118c: romdata_int = 'h36a9;
    'h118d: romdata_int = 'h3876;
    'h118e: romdata_int = 'h4000;
    'h118f: romdata_int = 'h54ba;
    'h1190: romdata_int = 'h70a8;
    'h1191: romdata_int = 'h7c00;
    'h1192: romdata_int = 'h829b;
    'h1193: romdata_int = 'h8cde;
    'h1194: romdata_int = 'hb678;
    'h1195: romdata_int = 'hb800;
    'h1196: romdata_int = 'he80c;
    'h1197: romdata_int = 'hf400;
    'h1198: romdata_int = 'h104cc;
    'h1199: romdata_int = 'h10961;
    'h119a: romdata_int = 'h531e; // Line descriptor for 5_6
    'h119b: romdata_int = 'he0;
    'h119c: romdata_int = 'h600;
    'h119d: romdata_int = 'h948;
    'h119e: romdata_int = 'ha7b;
    'h119f: romdata_int = 'h1060;
    'h11a0: romdata_int = 'h1761;
    'h11a1: romdata_int = 'h1962;
    'h11a2: romdata_int = 'h22f3;
    'h11a3: romdata_int = 'h4200;
    'h11a4: romdata_int = 'h44fa;
    'h11a5: romdata_int = 'h74f0;
    'h11a6: romdata_int = 'h7e00;
    'h11a7: romdata_int = 'h80d9;
    'h11a8: romdata_int = 'h9e0c;
    'h11a9: romdata_int = 'hb469;
    'h11aa: romdata_int = 'hba00;
    'h11ab: romdata_int = 'hde19;
    'h11ac: romdata_int = 'hf600;
    'h11ad: romdata_int = 'h11360;
    'h11ae: romdata_int = 'h1289c;
    'h11af: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11b0: romdata_int = 'h800;
    'h11b1: romdata_int = 'h905;
    'h11b2: romdata_int = 'haee;
    'h11b3: romdata_int = 'h1022;
    'h11b4: romdata_int = 'h1245;
    'h11b5: romdata_int = 'h1267;
    'h11b6: romdata_int = 'h160d;
    'h11b7: romdata_int = 'h1ed2;
    'h11b8: romdata_int = 'h4400;
    'h11b9: romdata_int = 'h4e84;
    'h11ba: romdata_int = 'h6e0d;
    'h11bb: romdata_int = 'h8000;
    'h11bc: romdata_int = 'h9a5f;
    'h11bd: romdata_int = 'haeca;
    'h11be: romdata_int = 'hbc00;
    'h11bf: romdata_int = 'hdb2e;
    'h11c0: romdata_int = 'he257;
    'h11c1: romdata_int = 'hf800;
    'h11c2: romdata_int = 'h1128e;
    'h11c3: romdata_int = 'h124d6;
    'h11c4: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11c5: romdata_int = 'h4a6;
    'h11c6: romdata_int = 'h553;
    'h11c7: romdata_int = 'h8a1;
    'h11c8: romdata_int = 'ha00;
    'h11c9: romdata_int = 'he9e;
    'h11ca: romdata_int = 'h1049;
    'h11cb: romdata_int = 'h1818;
    'h11cc: romdata_int = 'h1a7d;
    'h11cd: romdata_int = 'h4600;
    'h11ce: romdata_int = 'h606e;
    'h11cf: romdata_int = 'h6f13;
    'h11d0: romdata_int = 'h7f61;
    'h11d1: romdata_int = 'h8200;
    'h11d2: romdata_int = 'hb260;
    'h11d3: romdata_int = 'hb687;
    'h11d4: romdata_int = 'hbe00;
    'h11d5: romdata_int = 'he645;
    'h11d6: romdata_int = 'hfa00;
    'h11d7: romdata_int = 'h1092a;
    'h11d8: romdata_int = 'h1267d;
    'h11d9: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11da: romdata_int = 'h6b;
    'h11db: romdata_int = 'h74d;
    'h11dc: romdata_int = 'hc00;
    'h11dd: romdata_int = 'hd15;
    'h11de: romdata_int = 'he8b;
    'h11df: romdata_int = 'h127e;
    'h11e0: romdata_int = 'h1679;
    'h11e1: romdata_int = 'h22e2;
    'h11e2: romdata_int = 'h4800;
    'h11e3: romdata_int = 'h4b35;
    'h11e4: romdata_int = 'h5a96;
    'h11e5: romdata_int = 'h8400;
    'h11e6: romdata_int = 'h9331;
    'h11e7: romdata_int = 'hac97;
    'h11e8: romdata_int = 'hc000;
    'h11e9: romdata_int = 'hd70b;
    'h11ea: romdata_int = 'hdef4;
    'h11eb: romdata_int = 'hfc00;
    'h11ec: romdata_int = 'h10342;
    'h11ed: romdata_int = 'h11e46;
    'h11ee: romdata_int = 'h531e; // Line descriptor for 5_6
    'h11ef: romdata_int = 'h2d5;
    'h11f0: romdata_int = 'h4f2;
    'h11f1: romdata_int = 'h68f;
    'h11f2: romdata_int = 'he34;
    'h11f3: romdata_int = 'he00;
    'h11f4: romdata_int = 'he39;
    'h11f5: romdata_int = 'h2d3d;
    'h11f6: romdata_int = 'h3623;
    'h11f7: romdata_int = 'h4a00;
    'h11f8: romdata_int = 'h5ecd;
    'h11f9: romdata_int = 'h6825;
    'h11fa: romdata_int = 'h7c02;
    'h11fb: romdata_int = 'h8600;
    'h11fc: romdata_int = 'ha6c0;
    'h11fd: romdata_int = 'hb839;
    'h11fe: romdata_int = 'hc200;
    'h11ff: romdata_int = 'he89c;
    'h1200: romdata_int = 'hf105;
    'h1201: romdata_int = 'hf67a;
    'h1202: romdata_int = 'hfe00;
    'h1203: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1204: romdata_int = 'h32b;
    'h1205: romdata_int = 'h6ab;
    'h1206: romdata_int = 'h74f;
    'h1207: romdata_int = 'h1000;
    'h1208: romdata_int = 'h18fc;
    'h1209: romdata_int = 'h1b25;
    'h120a: romdata_int = 'h2d56;
    'h120b: romdata_int = 'h3908;
    'h120c: romdata_int = 'h4c00;
    'h120d: romdata_int = 'h4e0b;
    'h120e: romdata_int = 'h70d3;
    'h120f: romdata_int = 'h7cf1;
    'h1210: romdata_int = 'h8800;
    'h1211: romdata_int = 'h8f55;
    'h1212: romdata_int = 'hbd07;
    'h1213: romdata_int = 'hc400;
    'h1214: romdata_int = 'hc906;
    'h1215: romdata_int = 'h10000;
    'h1216: romdata_int = 'h104ec;
    'h1217: romdata_int = 'h11ae3;
    'h1218: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1219: romdata_int = 'h52c;
    'h121a: romdata_int = 'h84f;
    'h121b: romdata_int = 'hc17;
    'h121c: romdata_int = 'hcad;
    'h121d: romdata_int = 'h1038;
    'h121e: romdata_int = 'h1094;
    'h121f: romdata_int = 'h1200;
    'h1220: romdata_int = 'h1af7;
    'h1221: romdata_int = 'h4e00;
    'h1222: romdata_int = 'h6abb;
    'h1223: romdata_int = 'h7442;
    'h1224: romdata_int = 'h8a00;
    'h1225: romdata_int = 'h9b1a;
    'h1226: romdata_int = 'ha52e;
    'h1227: romdata_int = 'hc53c;
    'h1228: romdata_int = 'hc600;
    'h1229: romdata_int = 'hd264;
    'h122a: romdata_int = 'hf238;
    'h122b: romdata_int = 'h10200;
    'h122c: romdata_int = 'h10a78;
    'h122d: romdata_int = 'h531e; // Line descriptor for 5_6
    'h122e: romdata_int = 'h55;
    'h122f: romdata_int = 'h670;
    'h1230: romdata_int = 'h866;
    'h1231: romdata_int = 'h1230;
    'h1232: romdata_int = 'h1400;
    'h1233: romdata_int = 'h1cd9;
    'h1234: romdata_int = 'h24c6;
    'h1235: romdata_int = 'h30b9;
    'h1236: romdata_int = 'h4539;
    'h1237: romdata_int = 'h5000;
    'h1238: romdata_int = 'h6233;
    'h1239: romdata_int = 'h8c00;
    'h123a: romdata_int = 'h9838;
    'h123b: romdata_int = 'ha687;
    'h123c: romdata_int = 'hc800;
    'h123d: romdata_int = 'hce13;
    'h123e: romdata_int = 'heb4b;
    'h123f: romdata_int = 'h1006e;
    'h1240: romdata_int = 'h10400;
    'h1241: romdata_int = 'h10aed;
    'h1242: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1243: romdata_int = 'h264;
    'h1244: romdata_int = 'hb06;
    'h1245: romdata_int = 'hc42;
    'h1246: romdata_int = 'hd58;
    'h1247: romdata_int = 'h1600;
    'h1248: romdata_int = 'h171d;
    'h1249: romdata_int = 'h1854;
    'h124a: romdata_int = 'h1aee;
    'h124b: romdata_int = 'h5200;
    'h124c: romdata_int = 'h5a74;
    'h124d: romdata_int = 'h763b;
    'h124e: romdata_int = 'h7f26;
    'h124f: romdata_int = 'h8e00;
    'h1250: romdata_int = 'hb244;
    'h1251: romdata_int = 'hb564;
    'h1252: romdata_int = 'hca00;
    'h1253: romdata_int = 'he614;
    'h1254: romdata_int = 'h10600;
    'h1255: romdata_int = 'h120e5;
    'h1256: romdata_int = 'h12248;
    'h1257: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1258: romdata_int = 'h91;
    'h1259: romdata_int = 'h488;
    'h125a: romdata_int = 'hf66;
    'h125b: romdata_int = 'h1232;
    'h125c: romdata_int = 'h153b;
    'h125d: romdata_int = 'h1681;
    'h125e: romdata_int = 'h1800;
    'h125f: romdata_int = 'h3a7d;
    'h1260: romdata_int = 'h4a38;
    'h1261: romdata_int = 'h5400;
    'h1262: romdata_int = 'h5c8b;
    'h1263: romdata_int = 'h9000;
    'h1264: romdata_int = 'ha2df;
    'h1265: romdata_int = 'had28;
    'h1266: romdata_int = 'hc4de;
    'h1267: romdata_int = 'hcc00;
    'h1268: romdata_int = 'hcd30;
    'h1269: romdata_int = 'h10800;
    'h126a: romdata_int = 'h10f0c;
    'h126b: romdata_int = 'h12487;
    'h126c: romdata_int = 'h531e; // Line descriptor for 5_6
    'h126d: romdata_int = 'h11e;
    'h126e: romdata_int = 'h336;
    'h126f: romdata_int = 'h916;
    'h1270: romdata_int = 'hee5;
    'h1271: romdata_int = 'h131e;
    'h1272: romdata_int = 'h1836;
    'h1273: romdata_int = 'h1a00;
    'h1274: romdata_int = 'h1b13;
    'h1275: romdata_int = 'h54bd;
    'h1276: romdata_int = 'h5600;
    'h1277: romdata_int = 'h573d;
    'h1278: romdata_int = 'h9200;
    'h1279: romdata_int = 'hae1c;
    'h127a: romdata_int = 'hb0c4;
    'h127b: romdata_int = 'hcca1;
    'h127c: romdata_int = 'hce00;
    'h127d: romdata_int = 'hee2d;
    'h127e: romdata_int = 'h10a00;
    'h127f: romdata_int = 'h11c71;
    'h1280: romdata_int = 'h12081;
    'h1281: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1282: romdata_int = 'h60e;
    'h1283: romdata_int = 'ha45;
    'h1284: romdata_int = 'hc2b;
    'h1285: romdata_int = 'hf45;
    'h1286: romdata_int = 'h12b5;
    'h1287: romdata_int = 'h1711;
    'h1288: romdata_int = 'h1802;
    'h1289: romdata_int = 'h1c00;
    'h128a: romdata_int = 'h405c;
    'h128b: romdata_int = 'h5800;
    'h128c: romdata_int = 'h76ac;
    'h128d: romdata_int = 'h7a8c;
    'h128e: romdata_int = 'h8f40;
    'h128f: romdata_int = 'h9400;
    'h1290: romdata_int = 'hd000;
    'h1291: romdata_int = 'he305;
    'h1292: romdata_int = 'heb21;
    'h1293: romdata_int = 'hfa8d;
    'h1294: romdata_int = 'hfe83;
    'h1295: romdata_int = 'h10c00;
    'h1296: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1297: romdata_int = 'hd5;
    'h1298: romdata_int = 'ha72;
    'h1299: romdata_int = 'hadb;
    'h129a: romdata_int = 'h154c;
    'h129b: romdata_int = 'h1708;
    'h129c: romdata_int = 'h1c42;
    'h129d: romdata_int = 'h1e00;
    'h129e: romdata_int = 'h3212;
    'h129f: romdata_int = 'h3f41;
    'h12a0: romdata_int = 'h5a00;
    'h12a1: romdata_int = 'h66de;
    'h12a2: romdata_int = 'h910b;
    'h12a3: romdata_int = 'h9600;
    'h12a4: romdata_int = 'ha089;
    'h12a5: romdata_int = 'hd200;
    'h12a6: romdata_int = 'hd406;
    'h12a7: romdata_int = 'hd932;
    'h12a8: romdata_int = 'hfd55;
    'h12a9: romdata_int = 'h10e00;
    'h12aa: romdata_int = 'h11060;
    'h12ab: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12ac: romdata_int = 'h8a;
    'h12ad: romdata_int = 'h23b;
    'h12ae: romdata_int = 'h522;
    'h12af: romdata_int = 'ha3e;
    'h12b0: romdata_int = 'h10d8;
    'h12b1: romdata_int = 'h1cb5;
    'h12b2: romdata_int = 'h2000;
    'h12b3: romdata_int = 'h3a6b;
    'h12b4: romdata_int = 'h495c;
    'h12b5: romdata_int = 'h561e;
    'h12b6: romdata_int = 'h5c00;
    'h12b7: romdata_int = 'h7a70;
    'h12b8: romdata_int = 'h9800;
    'h12b9: romdata_int = 'ha533;
    'h12ba: romdata_int = 'hd400;
    'h12bb: romdata_int = 'hd832;
    'h12bc: romdata_int = 'he415;
    'h12bd: romdata_int = 'h102d3;
    'h12be: romdata_int = 'h11000;
    'h12bf: romdata_int = 'h114d8;
    'h12c0: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12c1: romdata_int = 'h262;
    'h12c2: romdata_int = 'h354;
    'h12c3: romdata_int = 'h45c;
    'h12c4: romdata_int = 'h84d;
    'h12c5: romdata_int = 'hc82;
    'h12c6: romdata_int = 'h12a8;
    'h12c7: romdata_int = 'h2200;
    'h12c8: romdata_int = 'h347f;
    'h12c9: romdata_int = 'h4d4e;
    'h12ca: romdata_int = 'h50a9;
    'h12cb: romdata_int = 'h5e00;
    'h12cc: romdata_int = 'h8ab7;
    'h12cd: romdata_int = 'h94eb;
    'h12ce: romdata_int = 'h9a00;
    'h12cf: romdata_int = 'hbe14;
    'h12d0: romdata_int = 'hc6f8;
    'h12d1: romdata_int = 'hd600;
    'h12d2: romdata_int = 'h11200;
    'h12d3: romdata_int = 'h11725;
    'h12d4: romdata_int = 'h12b0b;
    'h12d5: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12d6: romdata_int = 'h625;
    'h12d7: romdata_int = 'ha0b;
    'h12d8: romdata_int = 'he81;
    'h12d9: romdata_int = 'h143d;
    'h12da: romdata_int = 'h174c;
    'h12db: romdata_int = 'h1c19;
    'h12dc: romdata_int = 'h20d8;
    'h12dd: romdata_int = 'h2400;
    'h12de: romdata_int = 'h4c86;
    'h12df: romdata_int = 'h521c;
    'h12e0: romdata_int = 'h6000;
    'h12e1: romdata_int = 'h8706;
    'h12e2: romdata_int = 'h9c00;
    'h12e3: romdata_int = 'ha0e9;
    'h12e4: romdata_int = 'hd24b;
    'h12e5: romdata_int = 'hd800;
    'h12e6: romdata_int = 'heeea;
    'h12e7: romdata_int = 'hf74a;
    'h12e8: romdata_int = 'h10d31;
    'h12e9: romdata_int = 'h11400;
    'h12ea: romdata_int = 'h531e; // Line descriptor for 5_6
    'h12eb: romdata_int = 'ha5;
    'h12ec: romdata_int = 'h252;
    'h12ed: romdata_int = 'h290;
    'h12ee: romdata_int = 'h549;
    'h12ef: romdata_int = 'hf4d;
    'h12f0: romdata_int = 'h14d4;
    'h12f1: romdata_int = 'h2600;
    'h12f2: romdata_int = 'h2f37;
    'h12f3: romdata_int = 'h6200;
    'h12f4: romdata_int = 'h6687;
    'h12f5: romdata_int = 'h72aa;
    'h12f6: romdata_int = 'h7876;
    'h12f7: romdata_int = 'h842f;
    'h12f8: romdata_int = 'h9e00;
    'h12f9: romdata_int = 'hbc40;
    'h12fa: romdata_int = 'hd450;
    'h12fb: romdata_int = 'hda00;
    'h12fc: romdata_int = 'hf44e;
    'h12fd: romdata_int = 'h11600;
    'h12fe: romdata_int = 'h11842;
    'h12ff: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1300: romdata_int = 'hac3;
    'h1301: romdata_int = 'ha5c;
    'h1302: romdata_int = 'hb58;
    'h1303: romdata_int = 'h10b4;
    'h1304: romdata_int = 'h1c06;
    'h1305: romdata_int = 'h2800;
    'h1306: romdata_int = 'h2a27;
    'h1307: romdata_int = 'h351e;
    'h1308: romdata_int = 'h3c50;
    'h1309: romdata_int = 'h463d;
    'h130a: romdata_int = 'h6400;
    'h130b: romdata_int = 'h82b0;
    'h130c: romdata_int = 'h92bb;
    'h130d: romdata_int = 'ha000;
    'h130e: romdata_int = 'hc669;
    'h130f: romdata_int = 'hd135;
    'h1310: romdata_int = 'hdc00;
    'h1311: romdata_int = 'hf54f;
    'h1312: romdata_int = 'hf8e6;
    'h1313: romdata_int = 'h11800;
    'h1314: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1315: romdata_int = 'h8f3;
    'h1316: romdata_int = 'hc35;
    'h1317: romdata_int = 'hc67;
    'h1318: romdata_int = 'h1003;
    'h1319: romdata_int = 'h126e;
    'h131a: romdata_int = 'h1ce1;
    'h131b: romdata_int = 'h2a00;
    'h131c: romdata_int = 'h2e48;
    'h131d: romdata_int = 'h4243;
    'h131e: romdata_int = 'h42b1;
    'h131f: romdata_int = 'h6600;
    'h1320: romdata_int = 'h8028;
    'h1321: romdata_int = 'h8ca4;
    'h1322: romdata_int = 'ha200;
    'h1323: romdata_int = 'hcf3f;
    'h1324: romdata_int = 'hde00;
    'h1325: romdata_int = 'he0d1;
    'h1326: romdata_int = 'hf27e;
    'h1327: romdata_int = 'hfd04;
    'h1328: romdata_int = 'h11a00;
    'h1329: romdata_int = 'h531e; // Line descriptor for 5_6
    'h132a: romdata_int = 'h67;
    'h132b: romdata_int = 'h72d;
    'h132c: romdata_int = 'h1349;
    'h132d: romdata_int = 'h1559;
    'h132e: romdata_int = 'h1a45;
    'h132f: romdata_int = 'h1a52;
    'h1330: romdata_int = 'h1d28;
    'h1331: romdata_int = 'h2c00;
    'h1332: romdata_int = 'h4051;
    'h1333: romdata_int = 'h5f53;
    'h1334: romdata_int = 'h6800;
    'h1335: romdata_int = 'ha235;
    'h1336: romdata_int = 'ha400;
    'h1337: romdata_int = 'haab9;
    'h1338: romdata_int = 'hcb65;
    'h1339: romdata_int = 'hdb0c;
    'h133a: romdata_int = 'he000;
    'h133b: romdata_int = 'h10d2f;
    'h133c: romdata_int = 'h11b32;
    'h133d: romdata_int = 'h11c00;
    'h133e: romdata_int = 'h531e; // Line descriptor for 5_6
    'h133f: romdata_int = 'h10c8;
    'h1340: romdata_int = 'h14f3;
    'h1341: romdata_int = 'h1aa6;
    'h1342: romdata_int = 'h1b32;
    'h1343: romdata_int = 'h1c24;
    'h1344: romdata_int = 'h263b;
    'h1345: romdata_int = 'h2b45;
    'h1346: romdata_int = 'h2e00;
    'h1347: romdata_int = 'h5273;
    'h1348: romdata_int = 'h6a00;
    'h1349: romdata_int = 'h6d1a;
    'h134a: romdata_int = 'h9eb5;
    'h134b: romdata_int = 'ha600;
    'h134c: romdata_int = 'ha87c;
    'h134d: romdata_int = 'he07f;
    'h134e: romdata_int = 'he200;
    'h134f: romdata_int = 'he44c;
    'h1350: romdata_int = 'h10ece;
    'h1351: romdata_int = 'h11e00;
    'h1352: romdata_int = 'h11f2c;
    'h1353: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1354: romdata_int = 'h2b6;
    'h1355: romdata_int = 'h527;
    'h1356: romdata_int = 'h682;
    'h1357: romdata_int = 'h81a;
    'h1358: romdata_int = 'he99;
    'h1359: romdata_int = 'h28cd;
    'h135a: romdata_int = 'h2905;
    'h135b: romdata_int = 'h3000;
    'h135c: romdata_int = 'h4945;
    'h135d: romdata_int = 'h6c00;
    'h135e: romdata_int = 'h72cd;
    'h135f: romdata_int = 'h7830;
    'h1360: romdata_int = 'h8956;
    'h1361: romdata_int = 'ha800;
    'h1362: romdata_int = 'hc02d;
    'h1363: romdata_int = 'hc11c;
    'h1364: romdata_int = 'he400;
    'h1365: romdata_int = 'hf83f;
    'h1366: romdata_int = 'h11c39;
    'h1367: romdata_int = 'h12000;
    'h1368: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1369: romdata_int = 'h69f;
    'h136a: romdata_int = 'h752;
    'h136b: romdata_int = 'h1498;
    'h136c: romdata_int = 'h164f;
    'h136d: romdata_int = 'h1903;
    'h136e: romdata_int = 'h192f;
    'h136f: romdata_int = 'h1b50;
    'h1370: romdata_int = 'h3200;
    'h1371: romdata_int = 'h3cea;
    'h1372: romdata_int = 'h6a66;
    'h1373: romdata_int = 'h6e00;
    'h1374: romdata_int = 'h8893;
    'h1375: romdata_int = 'h9671;
    'h1376: romdata_int = 'haa00;
    'h1377: romdata_int = 'hdc45;
    'h1378: romdata_int = 'he600;
    'h1379: romdata_int = 'hec44;
    'h137a: romdata_int = 'h116fe;
    'h137b: romdata_int = 'h12200;
    'h137c: romdata_int = 'h12281;
    'h137d: romdata_int = 'h531e; // Line descriptor for 5_6
    'h137e: romdata_int = 'hd;
    'h137f: romdata_int = 'hc73;
    'h1380: romdata_int = 'h143a;
    'h1381: romdata_int = 'h14ba;
    'h1382: romdata_int = 'h1451;
    'h1383: romdata_int = 'h14d9;
    'h1384: romdata_int = 'h3233;
    'h1385: romdata_int = 'h3400;
    'h1386: romdata_int = 'h649e;
    'h1387: romdata_int = 'h6821;
    'h1388: romdata_int = 'h7000;
    'h1389: romdata_int = 'h9880;
    'h138a: romdata_int = 'h9cce;
    'h138b: romdata_int = 'hac00;
    'h138c: romdata_int = 'hbe06;
    'h138d: romdata_int = 'hc363;
    'h138e: romdata_int = 'he800;
    'h138f: romdata_int = 'h1155f;
    'h1390: romdata_int = 'h12400;
    'h1391: romdata_int = 'h1273d;
    'h1392: romdata_int = 'h531e; // Line descriptor for 5_6
    'h1393: romdata_int = 'h8ee;
    'h1394: romdata_int = 'he6b;
    'h1395: romdata_int = 'h1160;
    'h1396: romdata_int = 'h1734;
    'h1397: romdata_int = 'h18d5;
    'h1398: romdata_int = 'h18e4;
    'h1399: romdata_int = 'h1c96;
    'h139a: romdata_int = 'h3600;
    'h139b: romdata_int = 'h5888;
    'h139c: romdata_int = 'h6459;
    'h139d: romdata_int = 'h7200;
    'h139e: romdata_int = 'h972c;
    'h139f: romdata_int = 'ha933;
    'h13a0: romdata_int = 'hae00;
    'h13a1: romdata_int = 'hd0d0;
    'h13a2: romdata_int = 'hd633;
    'h13a3: romdata_int = 'hea00;
    'h13a4: romdata_int = 'h10704;
    'h13a5: romdata_int = 'h12600;
    'h13a6: romdata_int = 'h12af4;
    'h13a7: romdata_int = 'h531e; // Line descriptor for 5_6
    'h13a8: romdata_int = 'h2f2;
    'h13a9: romdata_int = 'h832;
    'h13aa: romdata_int = 'h1062;
    'h13ab: romdata_int = 'h151c;
    'h13ac: romdata_int = 'h16c6;
    'h13ad: romdata_int = 'h1d43;
    'h13ae: romdata_int = 'h2438;
    'h13af: romdata_int = 'h3800;
    'h13b0: romdata_int = 'h464d;
    'h13b1: romdata_int = 'h60bc;
    'h13b2: romdata_int = 'h7400;
    'h13b3: romdata_int = 'h9527;
    'h13b4: romdata_int = 'haae9;
    'h13b5: romdata_int = 'hb000;
    'h13b6: romdata_int = 'hb80a;
    'h13b7: romdata_int = 'hdd2a;
    'h13b8: romdata_int = 'hec00;
    'h13b9: romdata_int = 'hfefe;
    'h13ba: romdata_int = 'h100b6;
    'h13bb: romdata_int = 'h12800;
    'h13bc: romdata_int = 'h731e; // Line descriptor for 5_6
    'h13bd: romdata_int = 'h128;
    'h13be: romdata_int = 'h448;
    'h13bf: romdata_int = 'h80a;
    'h13c0: romdata_int = 'hcc5;
    'h13c1: romdata_int = 'h16f2;
    'h13c2: romdata_int = 'h2132;
    'h13c3: romdata_int = 'h3040;
    'h13c4: romdata_int = 'h3a00;
    'h13c5: romdata_int = 'h5833;
    'h13c6: romdata_int = 'h6272;
    'h13c7: romdata_int = 'h7600;
    'h13c8: romdata_int = 'h8544;
    'h13c9: romdata_int = 'hb10c;
    'h13ca: romdata_int = 'hb200;
    'h13cb: romdata_int = 'hba49;
    'h13cc: romdata_int = 'hbb35;
    'h13cd: romdata_int = 'hee00;
    'h13ce: romdata_int = 'hf03a;
    'h13cf: romdata_int = 'hfabc;
    'h13d0: romdata_int = 'h12a00;
    'h13d1: romdata_int = 'h5814; // Line descriptor for 8_9
    'h13d2: romdata_int = 'h0;
    'h13d3: romdata_int = 'h322;
    'h13d4: romdata_int = 'h1ec4;
    'h13d5: romdata_int = 'h22e7;
    'h13d6: romdata_int = 'h2800;
    'h13d7: romdata_int = 'h3338;
    'h13d8: romdata_int = 'h4479;
    'h13d9: romdata_int = 'h5000;
    'h13da: romdata_int = 'h6425;
    'h13db: romdata_int = 'h72ee;
    'h13dc: romdata_int = 'h7800;
    'h13dd: romdata_int = 'h9a1e;
    'h13de: romdata_int = 'h9e3f;
    'h13df: romdata_int = 'ha000;
    'h13e0: romdata_int = 'ha616;
    'h13e1: romdata_int = 'hb750;
    'h13e2: romdata_int = 'hc800;
    'h13e3: romdata_int = 'hdace;
    'h13e4: romdata_int = 'hdad6;
    'h13e5: romdata_int = 'hf000;
    'h13e6: romdata_int = 'hf35c;
    'h13e7: romdata_int = 'h110d8;
    'h13e8: romdata_int = 'h11800;
    'h13e9: romdata_int = 'h13050;
    'h13ea: romdata_int = 'h13222;
    'h13eb: romdata_int = 'h5814; // Line descriptor for 8_9
    'h13ec: romdata_int = 'h200;
    'h13ed: romdata_int = 'h75c;
    'h13ee: romdata_int = 'h10bc;
    'h13ef: romdata_int = 'h2277;
    'h13f0: romdata_int = 'h2a00;
    'h13f1: romdata_int = 'h3d48;
    'h13f2: romdata_int = 'h4631;
    'h13f3: romdata_int = 'h5200;
    'h13f4: romdata_int = 'h5650;
    'h13f5: romdata_int = 'h7733;
    'h13f6: romdata_int = 'h7a00;
    'h13f7: romdata_int = 'h7e35;
    'h13f8: romdata_int = 'h8523;
    'h13f9: romdata_int = 'ha200;
    'h13fa: romdata_int = 'hac4a;
    'h13fb: romdata_int = 'hb8e2;
    'h13fc: romdata_int = 'hca00;
    'h13fd: romdata_int = 'hd870;
    'h13fe: romdata_int = 'he74a;
    'h13ff: romdata_int = 'hf200;
    'h1400: romdata_int = 'h11132;
    'h1401: romdata_int = 'h112c6;
    'h1402: romdata_int = 'h11a00;
    'h1403: romdata_int = 'h1345a;
    'h1404: romdata_int = 'h13854;
    'h1405: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1406: romdata_int = 'ha1;
    'h1407: romdata_int = 'h400;
    'h1408: romdata_int = 'hf3d;
    'h1409: romdata_int = 'h224a;
    'h140a: romdata_int = 'h2c00;
    'h140b: romdata_int = 'h3b05;
    'h140c: romdata_int = 'h4cbe;
    'h140d: romdata_int = 'h5400;
    'h140e: romdata_int = 'h5719;
    'h140f: romdata_int = 'h6eeb;
    'h1410: romdata_int = 'h7c00;
    'h1411: romdata_int = 'h915d;
    'h1412: romdata_int = 'h98f2;
    'h1413: romdata_int = 'ha400;
    'h1414: romdata_int = 'hb6b5;
    'h1415: romdata_int = 'hc458;
    'h1416: romdata_int = 'hca67;
    'h1417: romdata_int = 'hcc00;
    'h1418: romdata_int = 'hd276;
    'h1419: romdata_int = 'hf400;
    'h141a: romdata_int = 'hf561;
    'h141b: romdata_int = 'h1007b;
    'h141c: romdata_int = 'h11c00;
    'h141d: romdata_int = 'h12904;
    'h141e: romdata_int = 'h12aec;
    'h141f: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1420: romdata_int = 'h600;
    'h1421: romdata_int = 'hab8;
    'h1422: romdata_int = 'h1a43;
    'h1423: romdata_int = 'h1b28;
    'h1424: romdata_int = 'h2e00;
    'h1425: romdata_int = 'h3475;
    'h1426: romdata_int = 'h48d0;
    'h1427: romdata_int = 'h5600;
    'h1428: romdata_int = 'h5b21;
    'h1429: romdata_int = 'h6a70;
    'h142a: romdata_int = 'h7e00;
    'h142b: romdata_int = 'h7ead;
    'h142c: romdata_int = 'h9ef5;
    'h142d: romdata_int = 'ha41d;
    'h142e: romdata_int = 'ha600;
    'h142f: romdata_int = 'hb4c8;
    'h1430: romdata_int = 'hce00;
    'h1431: romdata_int = 'he446;
    'h1432: romdata_int = 'he703;
    'h1433: romdata_int = 'hf600;
    'h1434: romdata_int = 'h10738;
    'h1435: romdata_int = 'h10cad;
    'h1436: romdata_int = 'h11e00;
    'h1437: romdata_int = 'h122ca;
    'h1438: romdata_int = 'h1387b;
    'h1439: romdata_int = 'h5814; // Line descriptor for 8_9
    'h143a: romdata_int = 'h800;
    'h143b: romdata_int = 'h939;
    'h143c: romdata_int = 'h120d;
    'h143d: romdata_int = 'h2052;
    'h143e: romdata_int = 'h2a4b;
    'h143f: romdata_int = 'h2c5f;
    'h1440: romdata_int = 'h3000;
    'h1441: romdata_int = 'h5800;
    'h1442: romdata_int = 'h581a;
    'h1443: romdata_int = 'h6693;
    'h1444: romdata_int = 'h8000;
    'h1445: romdata_int = 'h8eb3;
    'h1446: romdata_int = 'h94f8;
    'h1447: romdata_int = 'ha2a1;
    'h1448: romdata_int = 'ha800;
    'h1449: romdata_int = 'hba3a;
    'h144a: romdata_int = 'hd000;
    'h144b: romdata_int = 'hed35;
    'h144c: romdata_int = 'hef52;
    'h144d: romdata_int = 'hf6b4;
    'h144e: romdata_int = 'hf800;
    'h144f: romdata_int = 'h10884;
    'h1450: romdata_int = 'h12000;
    'h1451: romdata_int = 'h12a97;
    'h1452: romdata_int = 'h13cd6;
    'h1453: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1454: romdata_int = 'ha00;
    'h1455: romdata_int = 'ha79;
    'h1456: romdata_int = 'h18f3;
    'h1457: romdata_int = 'h192c;
    'h1458: romdata_int = 'h3200;
    'h1459: romdata_int = 'h3711;
    'h145a: romdata_int = 'h3eee;
    'h145b: romdata_int = 'h592c;
    'h145c: romdata_int = 'h5a00;
    'h145d: romdata_int = 'h7072;
    'h145e: romdata_int = 'h7a07;
    'h145f: romdata_int = 'h8200;
    'h1460: romdata_int = 'h98f6;
    'h1461: romdata_int = 'haa00;
    'h1462: romdata_int = 'hb267;
    'h1463: romdata_int = 'hbc62;
    'h1464: romdata_int = 'hd200;
    'h1465: romdata_int = 'hdd23;
    'h1466: romdata_int = 'he410;
    'h1467: romdata_int = 'hfa00;
    'h1468: romdata_int = 'hfe7d;
    'h1469: romdata_int = 'h11238;
    'h146a: romdata_int = 'h120c2;
    'h146b: romdata_int = 'h12200;
    'h146c: romdata_int = 'h12d10;
    'h146d: romdata_int = 'h5814; // Line descriptor for 8_9
    'h146e: romdata_int = 'hc00;
    'h146f: romdata_int = 'h1291;
    'h1470: romdata_int = 'h18a4;
    'h1471: romdata_int = 'h26bd;
    'h1472: romdata_int = 'h2934;
    'h1473: romdata_int = 'h3400;
    'h1474: romdata_int = 'h412a;
    'h1475: romdata_int = 'h5132;
    'h1476: romdata_int = 'h5c00;
    'h1477: romdata_int = 'h6280;
    'h1478: romdata_int = 'h78fd;
    'h1479: romdata_int = 'h7a41;
    'h147a: romdata_int = 'h8400;
    'h147b: romdata_int = 'ha937;
    'h147c: romdata_int = 'hac00;
    'h147d: romdata_int = 'hbe03;
    'h147e: romdata_int = 'hd400;
    'h147f: romdata_int = 'hd43d;
    'h1480: romdata_int = 'heaf2;
    'h1481: romdata_int = 'hfc00;
    'h1482: romdata_int = 'h100f0;
    'h1483: romdata_int = 'h10f09;
    'h1484: romdata_int = 'h11f37;
    'h1485: romdata_int = 'h12048;
    'h1486: romdata_int = 'h12400;
    'h1487: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1488: romdata_int = 'h42e;
    'h1489: romdata_int = 'ha60;
    'h148a: romdata_int = 'he00;
    'h148b: romdata_int = 'h1328;
    'h148c: romdata_int = 'h2e9f;
    'h148d: romdata_int = 'h2f2d;
    'h148e: romdata_int = 'h3600;
    'h148f: romdata_int = 'h5e00;
    'h1490: romdata_int = 'h6c2b;
    'h1491: romdata_int = 'h76b0;
    'h1492: romdata_int = 'h814c;
    'h1493: romdata_int = 'h8600;
    'h1494: romdata_int = 'h8c32;
    'h1495: romdata_int = 'had56;
    'h1496: romdata_int = 'hae00;
    'h1497: romdata_int = 'hb069;
    'h1498: romdata_int = 'hd600;
    'h1499: romdata_int = 'he31d;
    'h149a: romdata_int = 'hef64;
    'h149b: romdata_int = 'hfe00;
    'h149c: romdata_int = 'hfeaa;
    'h149d: romdata_int = 'h1074b;
    'h149e: romdata_int = 'h11b49;
    'h149f: romdata_int = 'h122c3;
    'h14a0: romdata_int = 'h12600;
    'h14a1: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14a2: romdata_int = 'h8e;
    'h14a3: romdata_int = 'h30b;
    'h14a4: romdata_int = 'h1000;
    'h14a5: romdata_int = 'h1079;
    'h14a6: romdata_int = 'h3800;
    'h14a7: romdata_int = 'h3a4f;
    'h14a8: romdata_int = 'h4ec5;
    'h14a9: romdata_int = 'h6000;
    'h14aa: romdata_int = 'h6661;
    'h14ab: romdata_int = 'h6946;
    'h14ac: romdata_int = 'h786b;
    'h14ad: romdata_int = 'h8800;
    'h14ae: romdata_int = 'h8cf6;
    'h14af: romdata_int = 'ha497;
    'h14b0: romdata_int = 'hb000;
    'h14b1: romdata_int = 'hb53f;
    'h14b2: romdata_int = 'hce3d;
    'h14b3: romdata_int = 'hd6e3;
    'h14b4: romdata_int = 'hd800;
    'h14b5: romdata_int = 'h10000;
    'h14b6: romdata_int = 'h1050b;
    'h14b7: romdata_int = 'h10afe;
    'h14b8: romdata_int = 'h12800;
    'h14b9: romdata_int = 'h12e5b;
    'h14ba: romdata_int = 'h13d1e;
    'h14bb: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14bc: romdata_int = 'hd3b;
    'h14bd: romdata_int = 'h1200;
    'h14be: romdata_int = 'h1ab0;
    'h14bf: romdata_int = 'h1ce5;
    'h14c0: romdata_int = 'h3a00;
    'h14c1: romdata_int = 'h4262;
    'h14c2: romdata_int = 'h42c1;
    'h14c3: romdata_int = 'h525f;
    'h14c4: romdata_int = 'h6200;
    'h14c5: romdata_int = 'h643e;
    'h14c6: romdata_int = 'h8a00;
    'h14c7: romdata_int = 'h908f;
    'h14c8: romdata_int = 'h9d45;
    'h14c9: romdata_int = 'ha0a8;
    'h14ca: romdata_int = 'hb052;
    'h14cb: romdata_int = 'hb200;
    'h14cc: romdata_int = 'hda00;
    'h14cd: romdata_int = 'he8e4;
    'h14ce: romdata_int = 'he93e;
    'h14cf: romdata_int = 'hfca6;
    'h14d0: romdata_int = 'h10200;
    'h14d1: romdata_int = 'h10cc2;
    'h14d2: romdata_int = 'h128d5;
    'h14d3: romdata_int = 'h12a00;
    'h14d4: romdata_int = 'h13685;
    'h14d5: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14d6: romdata_int = 'h404;
    'h14d7: romdata_int = 'he99;
    'h14d8: romdata_int = 'h1400;
    'h14d9: romdata_int = 'h1461;
    'h14da: romdata_int = 'h2c06;
    'h14db: romdata_int = 'h328f;
    'h14dc: romdata_int = 'h3c00;
    'h14dd: romdata_int = 'h542a;
    'h14de: romdata_int = 'h62ab;
    'h14df: romdata_int = 'h6400;
    'h14e0: romdata_int = 'h88c4;
    'h14e1: romdata_int = 'h8c00;
    'h14e2: romdata_int = 'h96dc;
    'h14e3: romdata_int = 'hb400;
    'h14e4: romdata_int = 'hbb60;
    'h14e5: romdata_int = 'hc094;
    'h14e6: romdata_int = 'hc830;
    'h14e7: romdata_int = 'hccf3;
    'h14e8: romdata_int = 'hdc00;
    'h14e9: romdata_int = 'hf487;
    'h14ea: romdata_int = 'hfa05;
    'h14eb: romdata_int = 'h10400;
    'h14ec: romdata_int = 'h12c00;
    'h14ed: romdata_int = 'h12e12;
    'h14ee: romdata_int = 'h1354e;
    'h14ef: romdata_int = 'h5814; // Line descriptor for 8_9
    'h14f0: romdata_int = 'h1600;
    'h14f1: romdata_int = 'h16ae;
    'h14f2: romdata_int = 'h203b;
    'h14f3: romdata_int = 'h2553;
    'h14f4: romdata_int = 'h3441;
    'h14f5: romdata_int = 'h3e00;
    'h14f6: romdata_int = 'h44b2;
    'h14f7: romdata_int = 'h5b06;
    'h14f8: romdata_int = 'h6040;
    'h14f9: romdata_int = 'h6600;
    'h14fa: romdata_int = 'h7c2b;
    'h14fb: romdata_int = 'h8a0a;
    'h14fc: romdata_int = 'h8e00;
    'h14fd: romdata_int = 'ha097;
    'h14fe: romdata_int = 'hb600;
    'h14ff: romdata_int = 'hbed8;
    'h1500: romdata_int = 'hd759;
    'h1501: romdata_int = 'hde00;
    'h1502: romdata_int = 'he111;
    'h1503: romdata_int = 'hf061;
    'h1504: romdata_int = 'h10600;
    'h1505: romdata_int = 'h11745;
    'h1506: romdata_int = 'h11c37;
    'h1507: romdata_int = 'h12e00;
    'h1508: romdata_int = 'h13b02;
    'h1509: romdata_int = 'h5814; // Line descriptor for 8_9
    'h150a: romdata_int = 'h2ae;
    'h150b: romdata_int = 'h83a;
    'h150c: romdata_int = 'h1800;
    'h150d: romdata_int = 'h1c6a;
    'h150e: romdata_int = 'h4000;
    'h150f: romdata_int = 'h4158;
    'h1510: romdata_int = 'h46e7;
    'h1511: romdata_int = 'h5c08;
    'h1512: romdata_int = 'h5c65;
    'h1513: romdata_int = 'h6800;
    'h1514: romdata_int = 'h84f6;
    'h1515: romdata_int = 'h9000;
    'h1516: romdata_int = 'h9250;
    'h1517: romdata_int = 'hae60;
    'h1518: romdata_int = 'hb800;
    'h1519: romdata_int = 'hc2e8;
    'h151a: romdata_int = 'hc880;
    'h151b: romdata_int = 'he000;
    'h151c: romdata_int = 'hed62;
    'h151d: romdata_int = 'h10800;
    'h151e: romdata_int = 'h10ad2;
    'h151f: romdata_int = 'h11627;
    'h1520: romdata_int = 'h12d3e;
    'h1521: romdata_int = 'h13000;
    'h1522: romdata_int = 'h13b2a;
    'h1523: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1524: romdata_int = 'h101e;
    'h1525: romdata_int = 'h14d5;
    'h1526: romdata_int = 'h16e6;
    'h1527: romdata_int = 'h1a00;
    'h1528: romdata_int = 'h387d;
    'h1529: romdata_int = 'h4200;
    'h152a: romdata_int = 'h4a30;
    'h152b: romdata_int = 'h521c;
    'h152c: romdata_int = 'h6a00;
    'h152d: romdata_int = 'h6cba;
    'h152e: romdata_int = 'h9200;
    'h152f: romdata_int = 'h9232;
    'h1530: romdata_int = 'h942f;
    'h1531: romdata_int = 'haedd;
    'h1532: romdata_int = 'hba00;
    'h1533: romdata_int = 'hbcb4;
    'h1534: romdata_int = 'hcf59;
    'h1535: romdata_int = 'he0bd;
    'h1536: romdata_int = 'he200;
    'h1537: romdata_int = 'hf638;
    'h1538: romdata_int = 'h108fd;
    'h1539: romdata_int = 'h10a00;
    'h153a: romdata_int = 'h1248f;
    'h153b: romdata_int = 'h12656;
    'h153c: romdata_int = 'h13200;
    'h153d: romdata_int = 'h5814; // Line descriptor for 8_9
    'h153e: romdata_int = 'hcb9;
    'h153f: romdata_int = 'hf65;
    'h1540: romdata_int = 'h1c00;
    'h1541: romdata_int = 'h252c;
    'h1542: romdata_int = 'h3e66;
    'h1543: romdata_int = 'h4400;
    'h1544: romdata_int = 'h4ebd;
    'h1545: romdata_int = 'h54c9;
    'h1546: romdata_int = 'h6c00;
    'h1547: romdata_int = 'h6e44;
    'h1548: romdata_int = 'h8115;
    'h1549: romdata_int = 'h8a9a;
    'h154a: romdata_int = 'h9400;
    'h154b: romdata_int = 'haa36;
    'h154c: romdata_int = 'hb8b8;
    'h154d: romdata_int = 'hbc00;
    'h154e: romdata_int = 'hdc17;
    'h154f: romdata_int = 'hde6b;
    'h1550: romdata_int = 'he400;
    'h1551: romdata_int = 'hf8b8;
    'h1552: romdata_int = 'h1020a;
    'h1553: romdata_int = 'h10c00;
    'h1554: romdata_int = 'h118c4;
    'h1555: romdata_int = 'h13267;
    'h1556: romdata_int = 'h13400;
    'h1557: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1558: romdata_int = 'h137;
    'h1559: romdata_int = 'hc7c;
    'h155a: romdata_int = 'h1cc9;
    'h155b: romdata_int = 'h1e00;
    'h155c: romdata_int = 'h3c1a;
    'h155d: romdata_int = 'h4600;
    'h155e: romdata_int = 'h48a0;
    'h155f: romdata_int = 'h5e5d;
    'h1560: romdata_int = 'h5e7b;
    'h1561: romdata_int = 'h6e00;
    'h1562: romdata_int = 'h8e3d;
    'h1563: romdata_int = 'h9600;
    'h1564: romdata_int = 'h96e3;
    'h1565: romdata_int = 'ha94c;
    'h1566: romdata_int = 'haaf4;
    'h1567: romdata_int = 'hbe00;
    'h1568: romdata_int = 'hd413;
    'h1569: romdata_int = 'he24f;
    'h156a: romdata_int = 'he600;
    'h156b: romdata_int = 'hfa43;
    'h156c: romdata_int = 'h10e00;
    'h156d: romdata_int = 'h1143b;
    'h156e: romdata_int = 'h12718;
    'h156f: romdata_int = 'h130ea;
    'h1570: romdata_int = 'h13600;
    'h1571: romdata_int = 'h5814; // Line descriptor for 8_9
    'h1572: romdata_int = 'h6e1;
    'h1573: romdata_int = 'h1455;
    'h1574: romdata_int = 'h2000;
    'h1575: romdata_int = 'h2549;
    'h1576: romdata_int = 'h2901;
    'h1577: romdata_int = 'h2ad9;
    'h1578: romdata_int = 'h4800;
    'h1579: romdata_int = 'h509f;
    'h157a: romdata_int = 'h6ab4;
    'h157b: romdata_int = 'h7000;
    'h157c: romdata_int = 'h86ed;
    'h157d: romdata_int = 'h873d;
    'h157e: romdata_int = 'h9800;
    'h157f: romdata_int = 'hc000;
    'h1580: romdata_int = 'hc059;
    'h1581: romdata_int = 'hc71e;
    'h1582: romdata_int = 'hd291;
    'h1583: romdata_int = 'he800;
    'h1584: romdata_int = 'hea2c;
    'h1585: romdata_int = 'hfd50;
    'h1586: romdata_int = 'h102d2;
    'h1587: romdata_int = 'h11000;
    'h1588: romdata_int = 'h11d49;
    'h1589: romdata_int = 'h13800;
    'h158a: romdata_int = 'h13e54;
    'h158b: romdata_int = 'h5814; // Line descriptor for 8_9
    'h158c: romdata_int = 'h489;
    'h158d: romdata_int = 'h8a1;
    'h158e: romdata_int = 'h1f50;
    'h158f: romdata_int = 'h2200;
    'h1590: romdata_int = 'h394a;
    'h1591: romdata_int = 'h4a00;
    'h1592: romdata_int = 'h4a9b;
    'h1593: romdata_int = 'h6018;
    'h1594: romdata_int = 'h7200;
    'h1595: romdata_int = 'h72c3;
    'h1596: romdata_int = 'h8323;
    'h1597: romdata_int = 'h9a00;
    'h1598: romdata_int = 'h9c78;
    'h1599: romdata_int = 'ha2b1;
    'h159a: romdata_int = 'hc200;
    'h159b: romdata_int = 'hc4ee;
    'h159c: romdata_int = 'hcce5;
    'h159d: romdata_int = 'hd033;
    'h159e: romdata_int = 'hea00;
    'h159f: romdata_int = 'hf29b;
    'h15a0: romdata_int = 'hf820;
    'h15a1: romdata_int = 'h11200;
    'h15a2: romdata_int = 'h11e48;
    'h15a3: romdata_int = 'h13644;
    'h15a4: romdata_int = 'h13a00;
    'h15a5: romdata_int = 'h5814; // Line descriptor for 8_9
    'h15a6: romdata_int = 'h212b;
    'h15a7: romdata_int = 'h2400;
    'h15a8: romdata_int = 'h2688;
    'h15a9: romdata_int = 'h2727;
    'h15aa: romdata_int = 'h314f;
    'h15ab: romdata_int = 'h4c00;
    'h15ac: romdata_int = 'h4d35;
    'h15ad: romdata_int = 'h70ea;
    'h15ae: romdata_int = 'h7400;
    'h15af: romdata_int = 'h74ca;
    'h15b0: romdata_int = 'h8814;
    'h15b1: romdata_int = 'h9b20;
    'h15b2: romdata_int = 'h9c00;
    'h15b3: romdata_int = 'ha6a2;
    'h15b4: romdata_int = 'hc2a0;
    'h15b5: romdata_int = 'hc400;
    'h15b6: romdata_int = 'hd8e6;
    'h15b7: romdata_int = 'hdf15;
    'h15b8: romdata_int = 'hec00;
    'h15b9: romdata_int = 'hf13d;
    'h15ba: romdata_int = 'h10e17;
    'h15bb: romdata_int = 'h11400;
    'h15bc: romdata_int = 'h1188a;
    'h15bd: romdata_int = 'h11aa1;
    'h15be: romdata_int = 'h13c00;
    'h15bf: romdata_int = 'h7814; // Line descriptor for 8_9
    'h15c0: romdata_int = 'h6ec;
    'h15c1: romdata_int = 'h1734;
    'h15c2: romdata_int = 'h1e4e;
    'h15c3: romdata_int = 'h2600;
    'h15c4: romdata_int = 'h3025;
    'h15c5: romdata_int = 'h3633;
    'h15c6: romdata_int = 'h4e00;
    'h15c7: romdata_int = 'h6890;
    'h15c8: romdata_int = 'h745c;
    'h15c9: romdata_int = 'h7600;
    'h15ca: romdata_int = 'h7c73;
    'h15cb: romdata_int = 'h8210;
    'h15cc: romdata_int = 'h9e00;
    'h15cd: romdata_int = 'hb269;
    'h15ce: romdata_int = 'hc600;
    'h15cf: romdata_int = 'hc645;
    'h15d0: romdata_int = 'hcb49;
    'h15d1: romdata_int = 'hd0cf;
    'h15d2: romdata_int = 'hee00;
    'h15d3: romdata_int = 'h10518;
    'h15d4: romdata_int = 'h1151c;
    'h15d5: romdata_int = 'h11600;
    'h15d6: romdata_int = 'h12555;
    'h15d7: romdata_int = 'h13e00;
    'h15d8: romdata_int = 'h13e48;
    'h15d9: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h15da: romdata_int = 'h0;
    'h15db: romdata_int = 'h322;
    'h15dc: romdata_int = 'h172c;
    'h15dd: romdata_int = 'h1ac4;
    'h15de: romdata_int = 'h2400;
    'h15df: romdata_int = 'h3538;
    'h15e0: romdata_int = 'h4679;
    'h15e1: romdata_int = 'h4800;
    'h15e2: romdata_int = 'h4ad0;
    'h15e3: romdata_int = 'h6a7e;
    'h15e4: romdata_int = 'h6c00;
    'h15e5: romdata_int = 'h7272;
    'h15e6: romdata_int = 'h8123;
    'h15e7: romdata_int = 'h9000;
    'h15e8: romdata_int = 'ha84a;
    'h15e9: romdata_int = 'hac67;
    'h15ea: romdata_int = 'hb400;
    'h15eb: romdata_int = 'hb608;
    'h15ec: romdata_int = 'hc2ed;
    'h15ed: romdata_int = 'hd800;
    'h15ee: romdata_int = 'he15c;
    'h15ef: romdata_int = 'hf8d8;
    'h15f0: romdata_int = 'hfc00;
    'h15f1: romdata_int = 'hfc5e;
    'h15f2: romdata_int = 'h1063a;
    'h15f3: romdata_int = 'h12000;
    'h15f4: romdata_int = 'h13241;
    'h15f5: romdata_int = 'h13440;
    'h15f6: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h15f7: romdata_int = 'h200;
    'h15f8: romdata_int = 'h75c;
    'h15f9: romdata_int = 'hebc;
    'h15fa: romdata_int = 'h1928;
    'h15fb: romdata_int = 'h2600;
    'h15fc: romdata_int = 'h3d05;
    'h15fd: romdata_int = 'h3f48;
    'h15fe: romdata_int = 'h4a00;
    'h15ff: romdata_int = 'h5850;
    'h1600: romdata_int = 'h5919;
    'h1601: romdata_int = 'h6e00;
    'h1602: romdata_int = 'h70eb;
    'h1603: romdata_int = 'h7cad;
    'h1604: romdata_int = 'h9200;
    'h1605: romdata_int = 'h961e;
    'h1606: romdata_int = 'haec8;
    'h1607: romdata_int = 'hb600;
    'h1608: romdata_int = 'hbc67;
    'h1609: romdata_int = 'hc8d6;
    'h160a: romdata_int = 'hda00;
    'h160b: romdata_int = 'hed28;
    'h160c: romdata_int = 'hee24;
    'h160d: romdata_int = 'hfe00;
    'h160e: romdata_int = 'h11824;
    'h160f: romdata_int = 'h11eea;
    'h1610: romdata_int = 'h12141;
    'h1611: romdata_int = 'h12200;
    'h1612: romdata_int = 'h13d2c;
    'h1613: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1614: romdata_int = 'ha1;
    'h1615: romdata_int = 'h400;
    'h1616: romdata_int = 'h100d;
    'h1617: romdata_int = 'h204a;
    'h1618: romdata_int = 'h2800;
    'h1619: romdata_int = 'h3675;
    'h161a: romdata_int = 'h44c1;
    'h161b: romdata_int = 'h4831;
    'h161c: romdata_int = 'h4c00;
    'h161d: romdata_int = 'h50bd;
    'h161e: romdata_int = 'h7000;
    'h161f: romdata_int = 'h74ee;
    'h1620: romdata_int = 'h7c35;
    'h1621: romdata_int = 'h9400;
    'h1622: romdata_int = 'h9ee5;
    'h1623: romdata_int = 'ha4f3;
    'h1624: romdata_int = 'hb800;
    'h1625: romdata_int = 'hc470;
    'h1626: romdata_int = 'hc8ce;
    'h1627: romdata_int = 'hdb21;
    'h1628: romdata_int = 'hdc00;
    'h1629: romdata_int = 'hf932;
    'h162a: romdata_int = 'h10000;
    'h162b: romdata_int = 'h11304;
    'h162c: romdata_int = 'h11e50;
    'h162d: romdata_int = 'h12400;
    'h162e: romdata_int = 'h12454;
    'h162f: romdata_int = 'h13f1a;
    'h1630: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1631: romdata_int = 'h600;
    'h1632: romdata_int = 'hab8;
    'h1633: romdata_int = 'h1843;
    'h1634: romdata_int = 'h2077;
    'h1635: romdata_int = 'h28bd;
    'h1636: romdata_int = 'h2a00;
    'h1637: romdata_int = 'h2e5f;
    'h1638: romdata_int = 'h4e00;
    'h1639: romdata_int = 'h4ebe;
    'h163a: romdata_int = 'h6825;
    'h163b: romdata_int = 'h7200;
    'h163c: romdata_int = 'h8ab3;
    'h163d: romdata_int = 'h8e32;
    'h163e: romdata_int = 'h9600;
    'h163f: romdata_int = 'h9c1d;
    'h1640: romdata_int = 'h9e3c;
    'h1641: romdata_int = 'hba00;
    'h1642: romdata_int = 'hd246;
    'h1643: romdata_int = 'hd503;
    'h1644: romdata_int = 'hd8b0;
    'h1645: romdata_int = 'hdd35;
    'h1646: romdata_int = 'hde00;
    'h1647: romdata_int = 'h10200;
    'h1648: romdata_int = 'h10eca;
    'h1649: romdata_int = 'h114a9;
    'h164a: romdata_int = 'h1247b;
    'h164b: romdata_int = 'h12600;
    'h164c: romdata_int = 'h1304b;
    'h164d: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h164e: romdata_int = 'h800;
    'h164f: romdata_int = 'h939;
    'h1650: romdata_int = 'ha79;
    'h1651: romdata_int = 'h1c52;
    'h1652: romdata_int = 'h2c00;
    'h1653: romdata_int = 'h2c4b;
    'h1654: romdata_int = 'h309f;
    'h1655: romdata_int = 'h5000;
    'h1656: romdata_int = 'h5a21;
    'h1657: romdata_int = 'h6680;
    'h1658: romdata_int = 'h7400;
    'h1659: romdata_int = 'h7a41;
    'h165a: romdata_int = 'h88f6;
    'h165b: romdata_int = 'h9800;
    'h165c: romdata_int = 'h9aa1;
    'h165d: romdata_int = 'ha081;
    'h165e: romdata_int = 'hb462;
    'h165f: romdata_int = 'hb4b4;
    'h1660: romdata_int = 'hbc00;
    'h1661: romdata_int = 'he000;
    'h1662: romdata_int = 'he4b4;
    'h1663: romdata_int = 'he6df;
    'h1664: romdata_int = 'hfd44;
    'h1665: romdata_int = 'h10400;
    'h1666: romdata_int = 'h10cc2;
    'h1667: romdata_int = 'h12800;
    'h1668: romdata_int = 'h13115;
    'h1669: romdata_int = 'h1372a;
    'h166a: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h166b: romdata_int = 'ha00;
    'h166c: romdata_int = 'h1091;
    'h166d: romdata_int = 'h16a4;
    'h166e: romdata_int = 'h20e7;
    'h166f: romdata_int = 'h252c;
    'h1670: romdata_int = 'h2e00;
    'h1671: romdata_int = 'h40ee;
    'h1672: romdata_int = 'h5200;
    'h1673: romdata_int = 'h5c1a;
    'h1674: romdata_int = 'h5d2c;
    'h1675: romdata_int = 'h7600;
    'h1676: romdata_int = 'h7733;
    'h1677: romdata_int = 'h7a07;
    'h1678: romdata_int = 'h94f2;
    'h1679: romdata_int = 'h94f6;
    'h167a: romdata_int = 'h9a00;
    'h167b: romdata_int = 'hb858;
    'h167c: romdata_int = 'hbe00;
    'h167d: romdata_int = 'hd210;
    'h167e: romdata_int = 'he200;
    'h167f: romdata_int = 'hf2d3;
    'h1680: romdata_int = 'hf4ad;
    'h1681: romdata_int = 'h10600;
    'h1682: romdata_int = 'h1095f;
    'h1683: romdata_int = 'h10b37;
    'h1684: romdata_int = 'h12a00;
    'h1685: romdata_int = 'h12a54;
    'h1686: romdata_int = 'h13e95;
    'h1687: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1688: romdata_int = 'h42e;
    'h1689: romdata_int = 'ha60;
    'h168a: romdata_int = 'hc00;
    'h168b: romdata_int = 'h1128;
    'h168c: romdata_int = 'h26a6;
    'h168d: romdata_int = 'h2b34;
    'h168e: romdata_int = 'h3000;
    'h168f: romdata_int = 'h50c5;
    'h1690: romdata_int = 'h5400;
    'h1691: romdata_int = 'h683e;
    'h1692: romdata_int = 'h7800;
    'h1693: romdata_int = 'h78fd;
    'h1694: romdata_int = 'h8832;
    'h1695: romdata_int = 'h9c00;
    'h1696: romdata_int = 'h9c97;
    'h1697: romdata_int = 'haf3f;
    'h1698: romdata_int = 'hbb1e;
    'h1699: romdata_int = 'hbe96;
    'h169a: romdata_int = 'hc000;
    'h169b: romdata_int = 'he291;
    'h169c: romdata_int = 'he400;
    'h169d: romdata_int = 'hf317;
    'h169e: romdata_int = 'h10800;
    'h169f: romdata_int = 'h10ec3;
    'h16a0: romdata_int = 'h11691;
    'h16a1: romdata_int = 'h128d6;
    'h16a2: romdata_int = 'h12c00;
    'h16a3: romdata_int = 'h12f25;
    'h16a4: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16a5: romdata_int = 'h8e;
    'h16a6: romdata_int = 'h30b;
    'h16a7: romdata_int = 'he00;
    'h16a8: romdata_int = 'he79;
    'h16a9: romdata_int = 'h312d;
    'h16aa: romdata_int = 'h3200;
    'h16ab: romdata_int = 'h3911;
    'h16ac: romdata_int = 'h48e7;
    'h16ad: romdata_int = 'h5332;
    'h16ae: romdata_int = 'h5600;
    'h16af: romdata_int = 'h7044;
    'h16b0: romdata_int = 'h74c3;
    'h16b1: romdata_int = 'h7a00;
    'h16b2: romdata_int = 'h9e00;
    'h16b3: romdata_int = 'ha337;
    'h16b4: romdata_int = 'ha956;
    'h16b5: romdata_int = 'hb677;
    'h16b6: romdata_int = 'hb8ee;
    'h16b7: romdata_int = 'hc200;
    'h16b8: romdata_int = 'he600;
    'h16b9: romdata_int = 'he87d;
    'h16ba: romdata_int = 'he8aa;
    'h16bb: romdata_int = 'h10a00;
    'h16bc: romdata_int = 'h10c48;
    'h16bd: romdata_int = 'h1107f;
    'h16be: romdata_int = 'h1291e;
    'h16bf: romdata_int = 'h12e00;
    'h16c0: romdata_int = 'h1384e;
    'h16c1: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16c2: romdata_int = 'hd3b;
    'h16c3: romdata_int = 'h1000;
    'h16c4: romdata_int = 'h16f3;
    'h16c5: romdata_int = 'h220e;
    'h16c6: romdata_int = 'h3400;
    'h16c7: romdata_int = 'h348f;
    'h16c8: romdata_int = 'h3c4f;
    'h16c9: romdata_int = 'h5800;
    'h16ca: romdata_int = 'h5f06;
    'h16cb: romdata_int = 'h5f21;
    'h16cc: romdata_int = 'h6e2b;
    'h16cd: romdata_int = 'h7c00;
    'h16ce: romdata_int = 'h7e3c;
    'h16cf: romdata_int = 'ha000;
    'h16d0: romdata_int = 'hb0b5;
    'h16d1: romdata_int = 'hb150;
    'h16d2: romdata_int = 'hc400;
    'h16d3: romdata_int = 'hcd55;
    'h16d4: romdata_int = 'hd762;
    'h16d5: romdata_int = 'hda75;
    'h16d6: romdata_int = 'he800;
    'h16d7: romdata_int = 'hec42;
    'h16d8: romdata_int = 'h10652;
    'h16d9: romdata_int = 'h10c00;
    'h16da: romdata_int = 'h11b5a;
    'h16db: romdata_int = 'h12caf;
    'h16dc: romdata_int = 'h13000;
    'h16dd: romdata_int = 'h142bc;
    'h16de: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16df: romdata_int = 'h404;
    'h16e0: romdata_int = 'h1200;
    'h16e1: romdata_int = 'h1261;
    'h16e2: romdata_int = 'h1ed5;
    'h16e3: romdata_int = 'h2e06;
    'h16e4: romdata_int = 'h3600;
    'h16e5: romdata_int = 'h3641;
    'h16e6: romdata_int = 'h545f;
    'h16e7: romdata_int = 'h562a;
    'h16e8: romdata_int = 'h5a00;
    'h16e9: romdata_int = 'h786b;
    'h16ea: romdata_int = 'h7e00;
    'h16eb: romdata_int = 'h8c8f;
    'h16ec: romdata_int = 'h902f;
    'h16ed: romdata_int = 'ha14d;
    'h16ee: romdata_int = 'ha200;
    'h16ef: romdata_int = 'hc226;
    'h16f0: romdata_int = 'hc600;
    'h16f1: romdata_int = 'hd54a;
    'h16f2: romdata_int = 'hea00;
    'h16f3: romdata_int = 'hf0fe;
    'h16f4: romdata_int = 'hf709;
    'h16f5: romdata_int = 'h10156;
    'h16f6: romdata_int = 'h10e00;
    'h16f7: romdata_int = 'h118b5;
    'h16f8: romdata_int = 'h12285;
    'h16f9: romdata_int = 'h13200;
    'h16fa: romdata_int = 'h14061;
    'h16fb: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h16fc: romdata_int = 'h1400;
    'h16fd: romdata_int = 'h14ae;
    'h16fe: romdata_int = 'h1c3b;
    'h16ff: romdata_int = 'h2283;
    'h1700: romdata_int = 'h3800;
    'h1701: romdata_int = 'h4066;
    'h1702: romdata_int = 'h432a;
    'h1703: romdata_int = 'h4c30;
    'h1704: romdata_int = 'h5c00;
    'h1705: romdata_int = 'h66ab;
    'h1706: romdata_int = 'h6d46;
    'h1707: romdata_int = 'h8000;
    'h1708: romdata_int = 'h869a;
    'h1709: romdata_int = 'h92dc;
    'h170a: romdata_int = 'ha400;
    'h170b: romdata_int = 'hb2b8;
    'h170c: romdata_int = 'hba45;
    'h170d: romdata_int = 'hc800;
    'h170e: romdata_int = 'hd11d;
    'h170f: romdata_int = 'hd904;
    'h1710: romdata_int = 'he438;
    'h1711: romdata_int = 'hec00;
    'h1712: romdata_int = 'h108e0;
    'h1713: romdata_int = 'h11000;
    'h1714: romdata_int = 'h1169c;
    'h1715: romdata_int = 'h13400;
    'h1716: romdata_int = 'h134f2;
    'h1717: romdata_int = 'h14011;
    'h1718: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1719: romdata_int = 'h2ae;
    'h171a: romdata_int = 'h83a;
    'h171b: romdata_int = 'h1600;
    'h171c: romdata_int = 'h18b0;
    'h171d: romdata_int = 'h3a00;
    'h171e: romdata_int = 'h3a7d;
    'h171f: romdata_int = 'h4462;
    'h1720: romdata_int = 'h4c9b;
    'h1721: romdata_int = 'h5e00;
    'h1722: romdata_int = 'h6008;
    'h1723: romdata_int = 'h6eba;
    'h1724: romdata_int = 'h8200;
    'h1725: romdata_int = 'h860a;
    'h1726: romdata_int = 'h90f8;
    'h1727: romdata_int = 'h92e3;
    'h1728: romdata_int = 'ha600;
    'h1729: romdata_int = 'hca00;
    'h172a: romdata_int = 'hcb1c;
    'h172b: romdata_int = 'hccb8;
    'h172c: romdata_int = 'hde61;
    'h172d: romdata_int = 'hee00;
    'h172e: romdata_int = 'hf0d2;
    'h172f: romdata_int = 'h1047b;
    'h1730: romdata_int = 'h11200;
    'h1731: romdata_int = 'h112d5;
    'h1732: romdata_int = 'h12737;
    'h1733: romdata_int = 'h13600;
    'h1734: romdata_int = 'h1426e;
    'h1735: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1736: romdata_int = 'hcb9;
    'h1737: romdata_int = 'he1e;
    'h1738: romdata_int = 'h12d5;
    'h1739: romdata_int = 'h1800;
    'h173a: romdata_int = 'h3c00;
    'h173b: romdata_int = 'h3e1a;
    'h173c: romdata_int = 'h46b2;
    'h173d: romdata_int = 'h541c;
    'h173e: romdata_int = 'h6000;
    'h173f: romdata_int = 'h6440;
    'h1740: romdata_int = 'h80f6;
    'h1741: romdata_int = 'h8400;
    'h1742: romdata_int = 'h84c4;
    'h1743: romdata_int = 'h983f;
    'h1744: romdata_int = 'ha636;
    'h1745: romdata_int = 'ha800;
    'h1746: romdata_int = 'hc0ba;
    'h1747: romdata_int = 'hcc00;
    'h1748: romdata_int = 'hd6fc;
    'h1749: romdata_int = 'hdd62;
    'h174a: romdata_int = 'heed9;
    'h174b: romdata_int = 'hf000;
    'h174c: romdata_int = 'h102c4;
    'h174d: romdata_int = 'h10560;
    'h174e: romdata_int = 'h11400;
    'h174f: romdata_int = 'h12058;
    'h1750: romdata_int = 'h13800;
    'h1751: romdata_int = 'h13c55;
    'h1752: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1753: romdata_int = 'h137;
    'h1754: romdata_int = 'h1a00;
    'h1755: romdata_int = 'h1e62;
    'h1756: romdata_int = 'h1ef2;
    'h1757: romdata_int = 'h285c;
    'h1758: romdata_int = 'h3b4a;
    'h1759: romdata_int = 'h3e00;
    'h175a: romdata_int = 'h56c9;
    'h175b: romdata_int = 'h5b38;
    'h175c: romdata_int = 'h6200;
    'h175d: romdata_int = 'h72ea;
    'h175e: romdata_int = 'h8600;
    'h175f: romdata_int = 'h8a3d;
    'h1760: romdata_int = 'ha457;
    'h1761: romdata_int = 'haa00;
    'h1762: romdata_int = 'hab29;
    'h1763: romdata_int = 'hca33;
    'h1764: romdata_int = 'hce00;
    'h1765: romdata_int = 'hce6b;
    'h1766: romdata_int = 'heaaa;
    'h1767: romdata_int = 'hf200;
    'h1768: romdata_int = 'hfaf3;
    'h1769: romdata_int = 'h1111e;
    'h176a: romdata_int = 'h11423;
    'h176b: romdata_int = 'h11600;
    'h176c: romdata_int = 'h12244;
    'h176d: romdata_int = 'h13a00;
    'h176e: romdata_int = 'h13b39;
    'h176f: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h1770: romdata_int = 'h6e1;
    'h1771: romdata_int = 'hc7c;
    'h1772: romdata_int = 'h14e6;
    'h1773: romdata_int = 'h1c00;
    'h1774: romdata_int = 'h26f2;
    'h1775: romdata_int = 'h2b01;
    'h1776: romdata_int = 'h4000;
    'h1777: romdata_int = 'h529f;
    'h1778: romdata_int = 'h6065;
    'h1779: romdata_int = 'h6400;
    'h177a: romdata_int = 'h82ed;
    'h177b: romdata_int = 'h8800;
    'h177c: romdata_int = 'h8d5d;
    'h177d: romdata_int = 'h9720;
    'h177e: romdata_int = 'ha34c;
    'h177f: romdata_int = 'hac00;
    'h1780: romdata_int = 'hbf0b;
    'h1781: romdata_int = 'hc629;
    'h1782: romdata_int = 'hd000;
    'h1783: romdata_int = 'he242;
    'h1784: romdata_int = 'hf400;
    'h1785: romdata_int = 'hf4c2;
    'h1786: romdata_int = 'hff1c;
    'h1787: romdata_int = 'h11800;
    'h1788: romdata_int = 'h11ca3;
    'h1789: romdata_int = 'h12627;
    'h178a: romdata_int = 'h13339;
    'h178b: romdata_int = 'h13c00;
    'h178c: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h178d: romdata_int = 'h489;
    'h178e: romdata_int = 'h1b50;
    'h178f: romdata_int = 'h1e00;
    'h1790: romdata_int = 'h2318;
    'h1791: romdata_int = 'h2cd9;
    'h1792: romdata_int = 'h3833;
    'h1793: romdata_int = 'h4200;
    'h1794: romdata_int = 'h625d;
    'h1795: romdata_int = 'h627b;
    'h1796: romdata_int = 'h6600;
    'h1797: romdata_int = 'h7ead;
    'h1798: romdata_int = 'h8414;
    'h1799: romdata_int = 'h8a00;
    'h179a: romdata_int = 'ha6f4;
    'h179b: romdata_int = 'haadc;
    'h179c: romdata_int = 'hae00;
    'h179d: romdata_int = 'hc674;
    'h179e: romdata_int = 'hd04f;
    'h179f: romdata_int = 'hd200;
    'h17a0: romdata_int = 'he09b;
    'h17a1: romdata_int = 'he725;
    'h17a2: romdata_int = 'hf600;
    'h17a3: romdata_int = 'h1013d;
    'h17a4: romdata_int = 'h1028a;
    'h17a5: romdata_int = 'h11a00;
    'h17a6: romdata_int = 'h12e92;
    'h17a7: romdata_int = 'h136c5;
    'h17a8: romdata_int = 'h13e00;
    'h17a9: romdata_int = 'h5b12; // Line descriptor for 9_10
    'h17aa: romdata_int = 'h8a1;
    'h17ab: romdata_int = 'h1255;
    'h17ac: romdata_int = 'h1d2b;
    'h17ad: romdata_int = 'h2000;
    'h17ae: romdata_int = 'h2553;
    'h17af: romdata_int = 'h4358;
    'h17b0: romdata_int = 'h4400;
    'h17b1: romdata_int = 'h4aa0;
    'h17b2: romdata_int = 'h6800;
    'h17b3: romdata_int = 'h6b3f;
    'h17b4: romdata_int = 'h76b0;
    'h17b5: romdata_int = 'h833d;
    'h17b6: romdata_int = 'h8c00;
    'h17b7: romdata_int = 'h98f5;
    'h17b8: romdata_int = 'h9ab1;
    'h17b9: romdata_int = 'hb000;
    'h17ba: romdata_int = 'hc4e6;
    'h17bb: romdata_int = 'hcf15;
    'h17bc: romdata_int = 'hd400;
    'h17bd: romdata_int = 'hdf3d;
    'h17be: romdata_int = 'hf800;
    'h17bf: romdata_int = 'hfae2;
    'h17c0: romdata_int = 'hfe3b;
    'h17c1: romdata_int = 'h11c00;
    'h17c2: romdata_int = 'h11c23;
    'h17c3: romdata_int = 'h12a48;
    'h17c4: romdata_int = 'h12c8d;
    'h17c5: romdata_int = 'h14000;
    'h17c6: romdata_int = 'h7b12; // Line descriptor for 9_10
    'h17c7: romdata_int = 'h6ec;
    'h17c8: romdata_int = 'h1534;
    'h17c9: romdata_int = 'h1a4e;
    'h17ca: romdata_int = 'h2200;
    'h17cb: romdata_int = 'h3225;
    'h17cc: romdata_int = 'h334f;
    'h17cd: romdata_int = 'h4600;
    'h17ce: romdata_int = 'h4f35;
    'h17cf: romdata_int = 'h6418;
    'h17d0: romdata_int = 'h6a00;
    'h17d1: romdata_int = 'h6c90;
    'h17d2: romdata_int = 'h8e00;
    'h17d3: romdata_int = 'h8e50;
    'h17d4: romdata_int = 'hac69;
    'h17d5: romdata_int = 'hb200;
    'h17d6: romdata_int = 'hb2e2;
    'h17d7: romdata_int = 'hbd49;
    'h17d8: romdata_int = 'hc051;
    'h17d9: romdata_int = 'hd600;
    'h17da: romdata_int = 'hea89;
    'h17db: romdata_int = 'hf617;
    'h17dc: romdata_int = 'hfa00;
    'h17dd: romdata_int = 'h10a48;
    'h17de: romdata_int = 'h11a20;
    'h17df: romdata_int = 'h11e00;
    'h17e0: romdata_int = 'h138c6;
    'h17e1: romdata_int = 'h13b02;
    'h17e2: romdata_int = 'h14200;
    'h17e3: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h17e4: romdata_int = 'h667;
    'h17e5: romdata_int = 'h4;
    'h17e6: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17e7: romdata_int = 'h6bd;
    'h17e8: romdata_int = 'ha5e;
    'h17e9: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17ea: romdata_int = 'h261;
    'h17eb: romdata_int = 'h334;
    'h17ec: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17ed: romdata_int = 'h4c9;
    'h17ee: romdata_int = 'he41;
    'h17ef: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17f0: romdata_int = 'h2e;
    'h17f1: romdata_int = 'h89;
    'h17f2: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17f3: romdata_int = 'h6a6;
    'h17f4: romdata_int = 'h2e0;
    'h17f5: romdata_int = 'h24; // Line descriptor for 1_5s
    'h17f6: romdata_int = 'h6f2;
    'h17f7: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h17f8: romdata_int = 'h137;
    'h17f9: romdata_int = 'h26b;
    'h17fa: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17fb: romdata_int = 'h4d5;
    'h17fc: romdata_int = 'h477;
    'h17fd: romdata_int = 'h124; // Line descriptor for 1_5s
    'h17fe: romdata_int = 'h92b;
    'h17ff: romdata_int = 'h108a;
    'h1800: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1801: romdata_int = 'h44a;
    'h1802: romdata_int = 'h52b;
    'h1803: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1804: romdata_int = 'hb0;
    'h1805: romdata_int = 'h255;
    'h1806: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1807: romdata_int = 'h688;
    'h1808: romdata_int = 'h1111;
    'h1809: romdata_int = 'h24; // Line descriptor for 1_5s
    'h180a: romdata_int = 'h464;
    'h180b: romdata_int = 'h24; // Line descriptor for 1_5s
    'h180c: romdata_int = 'h10b;
    'h180d: romdata_int = 'h4024; // Line descriptor for 1_5s
    'h180e: romdata_int = 'h86;
    'h180f: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1810: romdata_int = 'h8;
    'h1811: romdata_int = 'h2e6;
    'h1812: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1813: romdata_int = 'h536;
    'h1814: romdata_int = 'h31e;
    'h1815: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1816: romdata_int = 'hb2d;
    'h1817: romdata_int = 'h1161;
    'h1818: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1819: romdata_int = 'h855;
    'h181a: romdata_int = 'h2d5;
    'h181b: romdata_int = 'h24; // Line descriptor for 1_5s
    'h181c: romdata_int = 'h28a;
    'h181d: romdata_int = 'h124; // Line descriptor for 1_5s
    'h181e: romdata_int = 'h722;
    'h181f: romdata_int = 'h462;
    'h1820: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1821: romdata_int = 'hd4d;
    'h1822: romdata_int = 'h65c;
    'h1823: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h1824: romdata_int = 'h9a;
    'h1825: romdata_int = 'ha9f;
    'h1826: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1827: romdata_int = 'h490;
    'h1828: romdata_int = 'h2a5;
    'h1829: romdata_int = 'h124; // Line descriptor for 1_5s
    'h182a: romdata_int = 'h554;
    'h182b: romdata_int = 'h749;
    'h182c: romdata_int = 'h24; // Line descriptor for 1_5s
    'h182d: romdata_int = 'h267;
    'h182e: romdata_int = 'h24; // Line descriptor for 1_5s
    'h182f: romdata_int = 'hd5;
    'h1830: romdata_int = 'h24; // Line descriptor for 1_5s
    'h1831: romdata_int = 'hc25;
    'h1832: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1833: romdata_int = 'h15c;
    'h1834: romdata_int = 'he75;
    'h1835: romdata_int = 'h24; // Line descriptor for 1_5s
    'h1836: romdata_int = 'h727;
    'h1837: romdata_int = 'h4124; // Line descriptor for 1_5s
    'h1838: romdata_int = 'h4b6;
    'h1839: romdata_int = 'hae;
    'h183a: romdata_int = 'h124; // Line descriptor for 1_5s
    'h183b: romdata_int = 'h8d9;
    'h183c: romdata_int = 'h734;
    'h183d: romdata_int = 'h124; // Line descriptor for 1_5s
    'h183e: romdata_int = 'heab;
    'h183f: romdata_int = 'h701;
    'h1840: romdata_int = 'h124; // Line descriptor for 1_5s
    'h1841: romdata_int = 'h4f2;
    'h1842: romdata_int = 'hd52;
    'h1843: romdata_int = 'h2124; // Line descriptor for 1_5s
    'h1844: romdata_int = 'h328;
    'h1845: romdata_int = 'h648;
    'h1846: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1847: romdata_int = 'h48f;
    'h1848: romdata_int = 'h680;
    'h1849: romdata_int = 'h154b;
    'h184a: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h184b: romdata_int = 'h91d;
    'h184c: romdata_int = 'h2c9;
    'h184d: romdata_int = 'h83d;
    'h184e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h184f: romdata_int = 'h95d;
    'h1850: romdata_int = 'hcef;
    'h1851: romdata_int = 'h61;
    'h1852: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1853: romdata_int = 'h67b;
    'h1854: romdata_int = 'h12fc;
    'h1855: romdata_int = 'he0;
    'h1856: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1857: romdata_int = 'h425;
    'h1858: romdata_int = 'h1839;
    'h1859: romdata_int = 'h1c6f;
    'h185a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h185b: romdata_int = 'ha32;
    'h185c: romdata_int = 'h277;
    'h185d: romdata_int = 'h6cf;
    'h185e: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h185f: romdata_int = 'h2d5;
    'h1860: romdata_int = 'h6b;
    'h1861: romdata_int = 'h24a;
    'h1862: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1863: romdata_int = 'h552;
    'h1864: romdata_int = 'h65d;
    'h1865: romdata_int = 'h165a;
    'h1866: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1867: romdata_int = 'h32b;
    'h1868: romdata_int = 'hb03;
    'h1869: romdata_int = 'h1a81;
    'h186a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h186b: romdata_int = 'h4ab;
    'h186c: romdata_int = 'h54f;
    'h186d: romdata_int = 'h1740;
    'h186e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h186f: romdata_int = 'h55;
    'h1870: romdata_int = 'h6ab;
    'h1871: romdata_int = 'h1156;
    'h1872: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h1873: romdata_int = 'he83;
    'h1874: romdata_int = 'h264;
    'h1875: romdata_int = 'h44c;
    'h1876: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1877: romdata_int = 'he6;
    'h1878: romdata_int = 'h336;
    'h1879: romdata_int = 'habd;
    'h187a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h187b: romdata_int = 'h18e5;
    'h187c: romdata_int = 'h8b3;
    'h187d: romdata_int = 'h11e;
    'h187e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h187f: romdata_int = 'h40e;
    'h1880: romdata_int = 'h16a1;
    'h1881: romdata_int = 'h101e;
    'h1882: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1883: romdata_int = 'h832;
    'h1884: romdata_int = 'h441;
    'h1885: romdata_int = 'hd5;
    'h1886: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h1887: romdata_int = 'h722;
    'h1888: romdata_int = 'h8a;
    'h1889: romdata_int = 'h88f;
    'h188a: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h188b: romdata_int = 'h262;
    'h188c: romdata_int = 'h1d13;
    'h188d: romdata_int = 'h1d51;
    'h188e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h188f: romdata_int = 'h354;
    'h1890: romdata_int = 'h54d;
    'h1891: romdata_int = 'h14a8;
    'h1892: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1893: romdata_int = 'ha5;
    'h1894: romdata_int = 'h8a2;
    'h1895: romdata_int = 'h290;
    'h1896: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h1897: romdata_int = 'h8cb;
    'h1898: romdata_int = 'h6b4;
    'h1899: romdata_int = 'hce3;
    'h189a: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h189b: romdata_int = 'h640;
    'h189c: romdata_int = 'hef2;
    'h189d: romdata_int = 'h872;
    'h189e: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h189f: romdata_int = 'h1278;
    'h18a0: romdata_int = 'h698;
    'h18a1: romdata_int = 'h67;
    'h18a2: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18a3: romdata_int = 'h470;
    'h18a4: romdata_int = 'hcdc;
    'h18a5: romdata_int = 'h618;
    'h18a6: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18a7: romdata_int = 'h1497;
    'h18a8: romdata_int = 'h8f6;
    'h18a9: romdata_int = 'h538;
    'h18aa: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18ab: romdata_int = 'h2b6;
    'h18ac: romdata_int = 'h6fd;
    'h18ad: romdata_int = 'he74;
    'h18ae: romdata_int = 'h421e; // Line descriptor for 1_3s
    'h18af: romdata_int = 'hd;
    'h18b0: romdata_int = 'h475;
    'h18b1: romdata_int = 'h8a4;
    'h18b2: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18b3: romdata_int = 'h1b4d;
    'h18b4: romdata_int = 'h6eb;
    'h18b5: romdata_int = 'h186b;
    'h18b6: romdata_int = 'h21e; // Line descriptor for 1_3s
    'h18b7: romdata_int = 'h2f2;
    'h18b8: romdata_int = 'h1338;
    'h18b9: romdata_int = 'h1a9e;
    'h18ba: romdata_int = 'h221e; // Line descriptor for 1_3s
    'h18bb: romdata_int = 'h128;
    'h18bc: romdata_int = 'h93e;
    'h18bd: romdata_int = 'h1120;
    'h18be: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18bf: romdata_int = 'h6a4;
    'h18c0: romdata_int = 'h80c;
    'h18c1: romdata_int = 'hb67;
    'h18c2: romdata_int = 'h234a;
    'h18c3: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18c4: romdata_int = 'h2ba;
    'h18c5: romdata_int = 'h68c;
    'h18c6: romdata_int = 'h10ac;
    'h18c7: romdata_int = 'h1cf9;
    'h18c8: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18c9: romdata_int = 'h144;
    'h18ca: romdata_int = 'ha43;
    'h18cb: romdata_int = 'ha74;
    'h18cc: romdata_int = 'h1ac6;
    'h18cd: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18ce: romdata_int = 'h300;
    'h18cf: romdata_int = 'h445;
    'h18d0: romdata_int = 'h451;
    'h18d1: romdata_int = 'h1cd1;
    'h18d2: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18d3: romdata_int = 'h698;
    'h18d4: romdata_int = 'hc35;
    'h18d5: romdata_int = 'h113b;
    'h18d6: romdata_int = 'h20bd;
    'h18d7: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18d8: romdata_int = 'h8d9;
    'h18d9: romdata_int = 'h924;
    'h18da: romdata_int = 'hc3d;
    'h18db: romdata_int = 'h18b7;
    'h18dc: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18dd: romdata_int = 'h6fc;
    'h18de: romdata_int = 'h54c;
    'h18df: romdata_int = 'h8ed;
    'h18e0: romdata_int = 'h1b54;
    'h18e1: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18e2: romdata_int = 'ha95;
    'h18e3: romdata_int = 'h759;
    'h18e4: romdata_int = 'hd1;
    'h18e5: romdata_int = 'h1911;
    'h18e6: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18e7: romdata_int = 'h4e3;
    'h18e8: romdata_int = 'h89d;
    'h18e9: romdata_int = 'h6d9;
    'h18ea: romdata_int = 'h134c;
    'h18eb: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h18ec: romdata_int = 'h14f4;
    'h18ed: romdata_int = 'ha5d;
    'h18ee: romdata_int = 'h1b;
    'h18ef: romdata_int = 'hef2;
    'h18f0: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18f1: romdata_int = 'h20f;
    'h18f2: romdata_int = 'h2233;
    'h18f3: romdata_int = 'habe;
    'h18f4: romdata_int = 'h100;
    'h18f5: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18f6: romdata_int = 'h1ea4;
    'h18f7: romdata_int = 'h23e;
    'h18f8: romdata_int = 'h808;
    'h18f9: romdata_int = 'ha47;
    'h18fa: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h18fb: romdata_int = 'h41;
    'h18fc: romdata_int = 'h99;
    'h18fd: romdata_int = 'h547;
    'h18fe: romdata_int = 'h12d6;
    'h18ff: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1900: romdata_int = 'ha52;
    'h1901: romdata_int = 'h260;
    'h1902: romdata_int = 'h653;
    'h1903: romdata_int = 'h168e;
    'h1904: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1905: romdata_int = 'h447;
    'h1906: romdata_int = 'ha12;
    'h1907: romdata_int = 'h17;
    'h1908: romdata_int = 'h2262;
    'h1909: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h190a: romdata_int = 'h241;
    'h190b: romdata_int = 'h1757;
    'h190c: romdata_int = 'h41c;
    'h190d: romdata_int = 'hb59;
    'h190e: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h190f: romdata_int = 'h15;
    'h1910: romdata_int = 'hf6;
    'h1911: romdata_int = 'h1941;
    'h1912: romdata_int = 'h520;
    'h1913: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1914: romdata_int = 'h718;
    'h1915: romdata_int = 'h71f;
    'h1916: romdata_int = 'hd2e;
    'h1917: romdata_int = 'h1442;
    'h1918: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1919: romdata_int = 'hab2;
    'h191a: romdata_int = 'h1695;
    'h191b: romdata_int = 'he7c;
    'h191c: romdata_int = 'h730;
    'h191d: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h191e: romdata_int = 'h215d;
    'h191f: romdata_int = 'h2cf;
    'h1920: romdata_int = 'h946;
    'h1921: romdata_int = 'he8a;
    'h1922: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1923: romdata_int = 'h8a1;
    'h1924: romdata_int = 'h21f;
    'h1925: romdata_int = 'h1ea6;
    'h1926: romdata_int = 'h442;
    'h1927: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h1928: romdata_int = 'h31;
    'h1929: romdata_int = 'h14a3;
    'h192a: romdata_int = 'h965;
    'h192b: romdata_int = 'h276;
    'h192c: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h192d: romdata_int = 'h420;
    'h192e: romdata_int = 'h50c;
    'h192f: romdata_int = 'h1a49;
    'h1930: romdata_int = 'h8b0;
    'h1931: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1932: romdata_int = 'h1f39;
    'h1933: romdata_int = 'h6c7;
    'h1934: romdata_int = 'h493;
    'h1935: romdata_int = 'ha1d;
    'h1936: romdata_int = 'h31b; // Line descriptor for 2_5s
    'h1937: romdata_int = 'hf8;
    'h1938: romdata_int = 'h328;
    'h1939: romdata_int = 'h820;
    'h193a: romdata_int = 'h1d4d;
    'h193b: romdata_int = 'h431b; // Line descriptor for 2_5s
    'h193c: romdata_int = 'h746;
    'h193d: romdata_int = 'h12a;
    'h193e: romdata_int = 'h1157;
    'h193f: romdata_int = 'h210f;
    'h1940: romdata_int = 'h231b; // Line descriptor for 2_5s
    'h1941: romdata_int = 'h2d2;
    'h1942: romdata_int = 'h303;
    'h1943: romdata_int = 'h94b;
    'h1944: romdata_int = 'h1311;
    'h1945: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1946: romdata_int = 'ha00;
    'h1947: romdata_int = 'h129a;
    'h1948: romdata_int = 'h268a;
    'h1949: romdata_int = 'h319; // Line descriptor for 4_9s
    'h194a: romdata_int = 'h2eb;
    'h194b: romdata_int = 'h425;
    'h194c: romdata_int = 'h4e4;
    'h194d: romdata_int = 'hc00;
    'h194e: romdata_int = 'h4419; // Line descriptor for 4_9s
    'h194f: romdata_int = 'h8f8;
    'h1950: romdata_int = 'h670;
    'h1951: romdata_int = 'h68f;
    'h1952: romdata_int = 'h1d3b;
    'h1953: romdata_int = 'he00;
    'h1954: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1955: romdata_int = 'h2fd;
    'h1956: romdata_int = 'h850;
    'h1957: romdata_int = 'h1000;
    'h1958: romdata_int = 'h2279;
    'h1959: romdata_int = 'h119; // Line descriptor for 4_9s
    'h195a: romdata_int = 'hfe;
    'h195b: romdata_int = 'h1200;
    'h195c: romdata_int = 'h219; // Line descriptor for 4_9s
    'h195d: romdata_int = 'h1a7b;
    'h195e: romdata_int = 'h1400;
    'h195f: romdata_int = 'hc72;
    'h1960: romdata_int = 'h119; // Line descriptor for 4_9s
    'h1961: romdata_int = 'h1600;
    'h1962: romdata_int = 'h1ab8;
    'h1963: romdata_int = 'h4219; // Line descriptor for 4_9s
    'h1964: romdata_int = 'h48c;
    'h1965: romdata_int = 'h1800;
    'h1966: romdata_int = 'h242a;
    'h1967: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1968: romdata_int = 'h1cb9;
    'h1969: romdata_int = 'hce;
    'h196a: romdata_int = 'h102e;
    'h196b: romdata_int = 'h1a00;
    'h196c: romdata_int = 'h219; // Line descriptor for 4_9s
    'h196d: romdata_int = 'h1e9b;
    'h196e: romdata_int = 'h1c00;
    'h196f: romdata_int = 'hb15;
    'h1970: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1971: romdata_int = 'h82f;
    'h1972: romdata_int = 'h2165;
    'h1973: romdata_int = 'h1e00;
    'h1974: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1975: romdata_int = 'h5f;
    'h1976: romdata_int = 'ha2;
    'h1977: romdata_int = 'h2728;
    'h1978: romdata_int = 'h2000;
    'h1979: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h197a: romdata_int = 'he08;
    'h197b: romdata_int = 'h2200;
    'h197c: romdata_int = 'h2a;
    'h197d: romdata_int = 'h1c;
    'h197e: romdata_int = 'h319; // Line descriptor for 4_9s
    'h197f: romdata_int = 'h461;
    'h1980: romdata_int = 'h832;
    'h1981: romdata_int = 'h2400;
    'h1982: romdata_int = 'h24ef;
    'h1983: romdata_int = 'h319; // Line descriptor for 4_9s
    'h1984: romdata_int = 'h27b;
    'h1985: romdata_int = 'h1089;
    'h1986: romdata_int = 'h221e;
    'h1987: romdata_int = 'h2600;
    'h1988: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1989: romdata_int = 'h47f;
    'h198a: romdata_int = 'h8cd;
    'h198b: romdata_int = 'h140b;
    'h198c: romdata_int = 'h119; // Line descriptor for 4_9s
    'h198d: romdata_int = 'h62b;
    'h198e: romdata_int = 'hc02;
    'h198f: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h1990: romdata_int = 'h8bd;
    'h1991: romdata_int = 'h163a;
    'h1992: romdata_int = 'h1859;
    'h1993: romdata_int = 'h6ba;
    'h1994: romdata_int = 'h219; // Line descriptor for 4_9s
    'h1995: romdata_int = 'h265;
    'h1996: romdata_int = 'h493;
    'h1997: romdata_int = 'h1f12;
    'h1998: romdata_int = 'h119; // Line descriptor for 4_9s
    'h1999: romdata_int = 'hf0b;
    'h199a: romdata_int = 'h40a;
    'h199b: romdata_int = 'h319; // Line descriptor for 4_9s
    'h199c: romdata_int = 'h0;
    'h199d: romdata_int = 'hc9;
    'h199e: romdata_int = 'h6b4;
    'h199f: romdata_int = 'h1938;
    'h19a0: romdata_int = 'h219; // Line descriptor for 4_9s
    'h19a1: romdata_int = 'h200;
    'h19a2: romdata_int = 'haa1;
    'h19a3: romdata_int = 'h20c7;
    'h19a4: romdata_int = 'h4319; // Line descriptor for 4_9s
    'h19a5: romdata_int = 'h903;
    'h19a6: romdata_int = 'h400;
    'h19a7: romdata_int = 'h2c0;
    'h19a8: romdata_int = 'h12b0;
    'h19a9: romdata_int = 'h219; // Line descriptor for 4_9s
    'h19aa: romdata_int = 'h2e5;
    'h19ab: romdata_int = 'h600;
    'h19ac: romdata_int = 'h25d;
    'h19ad: romdata_int = 'h2419; // Line descriptor for 4_9s
    'h19ae: romdata_int = 'h16a1;
    'h19af: romdata_int = 'h14ec;
    'h19b0: romdata_int = 'h800;
    'h19b1: romdata_int = 'h6b1;
    'h19b2: romdata_int = 'h6d4;
    'h19b3: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19b4: romdata_int = 'h165;
    'h19b5: romdata_int = 'h4ac;
    'h19b6: romdata_int = 'h6ee;
    'h19b7: romdata_int = 'hcd4;
    'h19b8: romdata_int = 'h1016;
    'h19b9: romdata_int = 'h1077;
    'h19ba: romdata_int = 'h1200;
    'h19bb: romdata_int = 'h168b;
    'h19bc: romdata_int = 'h250f;
    'h19bd: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19be: romdata_int = 'h313;
    'h19bf: romdata_int = 'h567;
    'h19c0: romdata_int = 'h854;
    'h19c1: romdata_int = 'ha6f;
    'h19c2: romdata_int = 'hd42;
    'h19c3: romdata_int = 'h10e2;
    'h19c4: romdata_int = 'h1278;
    'h19c5: romdata_int = 'h1400;
    'h19c6: romdata_int = 'h34e8;
    'h19c7: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19c8: romdata_int = 'h216;
    'h19c9: romdata_int = 'h4df;
    'h19ca: romdata_int = 'h55f;
    'h19cb: romdata_int = 'hc5a;
    'h19cc: romdata_int = 'h1031;
    'h19cd: romdata_int = 'h113a;
    'h19ce: romdata_int = 'h1600;
    'h19cf: romdata_int = 'h2035;
    'h19d0: romdata_int = 'h32fd;
    'h19d1: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19d2: romdata_int = 'h228;
    'h19d3: romdata_int = 'h337;
    'h19d4: romdata_int = 'h43e;
    'h19d5: romdata_int = 'h958;
    'h19d6: romdata_int = 'haab;
    'h19d7: romdata_int = 'hb47;
    'h19d8: romdata_int = 'h1451;
    'h19d9: romdata_int = 'h1800;
    'h19da: romdata_int = 'h2cea;
    'h19db: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19dc: romdata_int = 'h1e;
    'h19dd: romdata_int = 'h79;
    'h19de: romdata_int = 'h245;
    'h19df: romdata_int = 'h109d;
    'h19e0: romdata_int = 'h1063;
    'h19e1: romdata_int = 'h1107;
    'h19e2: romdata_int = 'h1a00;
    'h19e3: romdata_int = 'h233c;
    'h19e4: romdata_int = 'h30bc;
    'h19e5: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19e6: romdata_int = 'h10b;
    'h19e7: romdata_int = 'h291;
    'h19e8: romdata_int = 'h61f;
    'h19e9: romdata_int = 'h708;
    'h19ea: romdata_int = 'h803;
    'h19eb: romdata_int = 'he3e;
    'h19ec: romdata_int = 'h1c00;
    'h19ed: romdata_int = 'h1c60;
    'h19ee: romdata_int = 'h2aa1;
    'h19ef: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h19f0: romdata_int = 'h4c;
    'h19f1: romdata_int = 'h526;
    'h19f2: romdata_int = 'ha94;
    'h19f3: romdata_int = 'haf2;
    'h19f4: romdata_int = 'he79;
    'h19f5: romdata_int = 'h104b;
    'h19f6: romdata_int = 'h1e00;
    'h19f7: romdata_int = 'h1ed2;
    'h19f8: romdata_int = 'h2f21;
    'h19f9: romdata_int = 'h812; // Line descriptor for 3_5s
    'h19fa: romdata_int = 'h13d;
    'h19fb: romdata_int = 'h512;
    'h19fc: romdata_int = 'h6af;
    'h19fd: romdata_int = 'h8e9;
    'h19fe: romdata_int = 'hc2d;
    'h19ff: romdata_int = 'hc80;
    'h1a00: romdata_int = 'h1293;
    'h1a01: romdata_int = 'h2000;
    'h1a02: romdata_int = 'h26b4;
    'h1a03: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a04: romdata_int = 'hef;
    'h1a05: romdata_int = 'had3;
    'h1a06: romdata_int = 'hca1;
    'h1a07: romdata_int = 'hd32;
    'h1a08: romdata_int = 'hf0f;
    'h1a09: romdata_int = 'hf39;
    'h1a0a: romdata_int = 'h20ee;
    'h1a0b: romdata_int = 'h2200;
    'h1a0c: romdata_int = 'h2ac7;
    'h1a0d: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a0e: romdata_int = 'h6e7;
    'h1a0f: romdata_int = 'h8a6;
    'h1a10: romdata_int = 'h8d3;
    'h1a11: romdata_int = 'hb1d;
    'h1a12: romdata_int = 'hb2c;
    'h1a13: romdata_int = 'hcb6;
    'h1a14: romdata_int = 'h1b4c;
    'h1a15: romdata_int = 'h2400;
    'h1a16: romdata_int = 'h2f05;
    'h1a17: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a18: romdata_int = 'hbc;
    'h1a19: romdata_int = 'h55a;
    'h1a1a: romdata_int = 'h6bd;
    'h1a1b: romdata_int = 'h8f8;
    'h1a1c: romdata_int = 'hacf;
    'h1a1d: romdata_int = 'hf4e;
    'h1a1e: romdata_int = 'h1e6b;
    'h1a1f: romdata_int = 'h2600;
    'h1a20: romdata_int = 'h2c8e;
    'h1a21: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a22: romdata_int = 'h99;
    'h1a23: romdata_int = 'h672;
    'h1a24: romdata_int = 'h687;
    'h1a25: romdata_int = 'h85f;
    'h1a26: romdata_int = 'hc30;
    'h1a27: romdata_int = 'he81;
    'h1a28: romdata_int = 'h18dc;
    'h1a29: romdata_int = 'h2800;
    'h1a2a: romdata_int = 'h2908;
    'h1a2b: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a2c: romdata_int = 'h27a;
    'h1a2d: romdata_int = 'h2a2;
    'h1a2e: romdata_int = 'h40b;
    'h1a2f: romdata_int = 'h73a;
    'h1a30: romdata_int = 'hb62;
    'h1a31: romdata_int = 'he66;
    'h1a32: romdata_int = 'h144c;
    'h1a33: romdata_int = 'h2a00;
    'h1a34: romdata_int = 'h3510;
    'h1a35: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a36: romdata_int = 'h20b;
    'h1a37: romdata_int = 'h20e;
    'h1a38: romdata_int = 'hb42;
    'h1a39: romdata_int = 'he5e;
    'h1a3a: romdata_int = 'hec7;
    'h1a3b: romdata_int = 'h10d9;
    'h1a3c: romdata_int = 'h183a;
    'h1a3d: romdata_int = 'h28da;
    'h1a3e: romdata_int = 'h2c00;
    'h1a3f: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a40: romdata_int = 'h9d;
    'h1a41: romdata_int = 'hc7;
    'h1a42: romdata_int = 'h506;
    'h1a43: romdata_int = 'h6db;
    'h1a44: romdata_int = 'h817;
    'h1a45: romdata_int = 'heeb;
    'h1a46: romdata_int = 'h1b50;
    'h1a47: romdata_int = 'h240e;
    'h1a48: romdata_int = 'h2e00;
    'h1a49: romdata_int = 'h812; // Line descriptor for 3_5s
    'h1a4a: romdata_int = 'h2a;
    'h1a4b: romdata_int = 'h33e;
    'h1a4c: romdata_int = 'h74f;
    'h1a4d: romdata_int = 'hc45;
    'h1a4e: romdata_int = 'hcc4;
    'h1a4f: romdata_int = 'hf2c;
    'h1a50: romdata_int = 'h22bd;
    'h1a51: romdata_int = 'h3000;
    'h1a52: romdata_int = 'h331b;
    'h1a53: romdata_int = 'h4812; // Line descriptor for 3_5s
    'h1a54: romdata_int = 'h4ed;
    'h1a55: romdata_int = 'h75f;
    'h1a56: romdata_int = 'h886;
    'h1a57: romdata_int = 'h828;
    'h1a58: romdata_int = 'h906;
    'h1a59: romdata_int = 'hafb;
    'h1a5a: romdata_int = 'h1d4e;
    'h1a5b: romdata_int = 'h30da;
    'h1a5c: romdata_int = 'h3200;
    'h1a5d: romdata_int = 'h2812; // Line descriptor for 3_5s
    'h1a5e: romdata_int = 'h34c;
    'h1a5f: romdata_int = 'h540;
    'h1a60: romdata_int = 'hc42;
    'h1a61: romdata_int = 'he0f;
    'h1a62: romdata_int = 'h1047;
    'h1a63: romdata_int = 'h10a3;
    'h1a64: romdata_int = 'h16cd;
    'h1a65: romdata_int = 'h2710;
    'h1a66: romdata_int = 'h3400;
    'h1a67: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a68: romdata_int = 'h0;
    'h1a69: romdata_int = 'h134;
    'h1a6a: romdata_int = 'h2c0;
    'h1a6b: romdata_int = 'h162f;
    'h1a6c: romdata_int = 'h16bd;
    'h1a6d: romdata_int = 'h1e00;
    'h1a6e: romdata_int = 'h2443;
    'h1a6f: romdata_int = 'h2e68;
    'h1a70: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a71: romdata_int = 'hd5;
    'h1a72: romdata_int = 'he6;
    'h1a73: romdata_int = 'h200;
    'h1a74: romdata_int = 'h265;
    'h1a75: romdata_int = 'h1533;
    'h1a76: romdata_int = 'h1ea9;
    'h1a77: romdata_int = 'h2000;
    'h1a78: romdata_int = 'h2c0f;
    'h1a79: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a7a: romdata_int = 'h208;
    'h1a7b: romdata_int = 'h27b;
    'h1a7c: romdata_int = 'h400;
    'h1a7d: romdata_int = 'h407;
    'h1a7e: romdata_int = 'h88f;
    'h1a7f: romdata_int = 'h2200;
    'h1a80: romdata_int = 'h2755;
    'h1a81: romdata_int = 'h2a17;
    'h1a82: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a83: romdata_int = 'h67;
    'h1a84: romdata_int = 'h2cf;
    'h1a85: romdata_int = 'h600;
    'h1a86: romdata_int = 'he10;
    'h1a87: romdata_int = 'h1c74;
    'h1a88: romdata_int = 'h20ac;
    'h1a89: romdata_int = 'h2400;
    'h1a8a: romdata_int = 'h32c3;
    'h1a8b: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a8c: romdata_int = 'h2eb;
    'h1a8d: romdata_int = 'h2fd;
    'h1a8e: romdata_int = 'h411;
    'h1a8f: romdata_int = 'h6eb;
    'h1a90: romdata_int = 'h800;
    'h1a91: romdata_int = 'h2600;
    'h1a92: romdata_int = 'h3870;
    'h1a93: romdata_int = 'h3a4b;
    'h1a94: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1a95: romdata_int = 'h61;
    'h1a96: romdata_int = 'h4d0;
    'h1a97: romdata_int = 'ha00;
    'h1a98: romdata_int = 'ha7d;
    'h1a99: romdata_int = 'hd47;
    'h1a9a: romdata_int = 'h2800;
    'h1a9b: romdata_int = 'h306d;
    'h1a9c: romdata_int = 'h362a;
    'h1a9d: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1a9e: romdata_int = 'ha5;
    'h1a9f: romdata_int = 'h50a;
    'h1aa0: romdata_int = 'hb42;
    'h1aa1: romdata_int = 'hc00;
    'h1aa2: romdata_int = 'h18e4;
    'h1aa3: romdata_int = 'h2a00;
    'h1aa4: romdata_int = 'h2d1e;
    'h1aa5: romdata_int = 'h380f;
    'h1aa6: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1aa7: romdata_int = 'h11e;
    'h1aa8: romdata_int = 'h560;
    'h1aa9: romdata_int = 'he00;
    'h1aaa: romdata_int = 'h1290;
    'h1aab: romdata_int = 'h12a7;
    'h1aac: romdata_int = 'h275b;
    'h1aad: romdata_int = 'h2c00;
    'h1aae: romdata_int = 'h2e20;
    'h1aaf: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ab0: romdata_int = 'h6b;
    'h1ab1: romdata_int = 'h322;
    'h1ab2: romdata_int = 'h4ff;
    'h1ab3: romdata_int = 'h1000;
    'h1ab4: romdata_int = 'h1b00;
    'h1ab5: romdata_int = 'h2526;
    'h1ab6: romdata_int = 'h2e00;
    'h1ab7: romdata_int = 'h3425;
    'h1ab8: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1ab9: romdata_int = 'he0;
    'h1aba: romdata_int = 'h439;
    'h1abb: romdata_int = 'h4e2;
    'h1abc: romdata_int = 'hd01;
    'h1abd: romdata_int = 'h1200;
    'h1abe: romdata_int = 'h3000;
    'h1abf: romdata_int = 'h349d;
    'h1ac0: romdata_int = 'h3b03;
    'h1ac1: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ac2: romdata_int = 'h49c;
    'h1ac3: romdata_int = 'h4b0;
    'h1ac4: romdata_int = 'h1400;
    'h1ac5: romdata_int = 'h189d;
    'h1ac6: romdata_int = 'h1c5a;
    'h1ac7: romdata_int = 'h204e;
    'h1ac8: romdata_int = 'h288f;
    'h1ac9: romdata_int = 'h3200;
    'h1aca: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1acb: romdata_int = 'h55;
    'h1acc: romdata_int = 'h240;
    'h1acd: romdata_int = 'h105f;
    'h1ace: romdata_int = 'h10c8;
    'h1acf: romdata_int = 'h1600;
    'h1ad0: romdata_int = 'h2ab3;
    'h1ad1: romdata_int = 'h3105;
    'h1ad2: romdata_int = 'h3400;
    'h1ad3: romdata_int = 'h470f; // Line descriptor for 2_3s
    'h1ad4: romdata_int = 'hae;
    'h1ad5: romdata_int = 'h25d;
    'h1ad6: romdata_int = 'h616;
    'h1ad7: romdata_int = 'he66;
    'h1ad8: romdata_int = 'h1800;
    'h1ad9: romdata_int = 'h2266;
    'h1ada: romdata_int = 'h28c2;
    'h1adb: romdata_int = 'h3600;
    'h1adc: romdata_int = 'h70f; // Line descriptor for 2_3s
    'h1add: romdata_int = 'h218;
    'h1ade: romdata_int = 'h2e5;
    'h1adf: romdata_int = 'h917;
    'h1ae0: romdata_int = 'h1442;
    'h1ae1: romdata_int = 'h1a00;
    'h1ae2: romdata_int = 'h1e0a;
    'h1ae3: romdata_int = 'h362d;
    'h1ae4: romdata_int = 'h3800;
    'h1ae5: romdata_int = 'h670f; // Line descriptor for 2_3s
    'h1ae6: romdata_int = 'h8a;
    'h1ae7: romdata_int = 'h40a;
    'h1ae8: romdata_int = 'h43d;
    'h1ae9: romdata_int = 'h1aa4;
    'h1aea: romdata_int = 'h1c00;
    'h1aeb: romdata_int = 'h2221;
    'h1aec: romdata_int = 'h3209;
    'h1aed: romdata_int = 'h3a00;
    'h1aee: romdata_int = 'h70c; // Line descriptor for 11_15s
    'h1aef: romdata_int = 'hda;
    'h1af0: romdata_int = 'h1052;
    'h1af1: romdata_int = 'h1200;
    'h1af2: romdata_int = 'h168f;
    'h1af3: romdata_int = 'h180b;
    'h1af4: romdata_int = 'h2a00;
    'h1af5: romdata_int = 'h36d3;
    'h1af6: romdata_int = 'h40ea;
    'h1af7: romdata_int = 'h490c; // Line descriptor for 11_15s
    'h1af8: romdata_int = 'h54;
    'h1af9: romdata_int = 'h96;
    'h1afa: romdata_int = 'h719;
    'h1afb: romdata_int = 'hb58;
    'h1afc: romdata_int = 'h1400;
    'h1afd: romdata_int = 'h22a2;
    'h1afe: romdata_int = 'h2959;
    'h1aff: romdata_int = 'h2c00;
    'h1b00: romdata_int = 'h3053;
    'h1b01: romdata_int = 'h3318;
    'h1b02: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b03: romdata_int = 'h2e;
    'h1b04: romdata_int = 'h93f;
    'h1b05: romdata_int = 'he59;
    'h1b06: romdata_int = 'h1600;
    'h1b07: romdata_int = 'h1a35;
    'h1b08: romdata_int = 'h202d;
    'h1b09: romdata_int = 'h2e00;
    'h1b0a: romdata_int = 'h3452;
    'h1b0b: romdata_int = 'h3a6c;
    'h1b0c: romdata_int = 'h460c; // Line descriptor for 11_15s
    'h1b0d: romdata_int = 'h0;
    'h1b0e: romdata_int = 'h14fa;
    'h1b0f: romdata_int = 'h1800;
    'h1b10: romdata_int = 'h1d1f;
    'h1b11: romdata_int = 'h3000;
    'h1b12: romdata_int = 'h3145;
    'h1b13: romdata_int = 'h3c33;
    'h1b14: romdata_int = 'h70c; // Line descriptor for 11_15s
    'h1b15: romdata_int = 'ha0;
    'h1b16: romdata_int = 'h200;
    'h1b17: romdata_int = 'h1a00;
    'h1b18: romdata_int = 'h2422;
    'h1b19: romdata_int = 'h24a2;
    'h1b1a: romdata_int = 'h3200;
    'h1b1b: romdata_int = 'h3e89;
    'h1b1c: romdata_int = 'h3f03;
    'h1b1d: romdata_int = 'h4a0c; // Line descriptor for 11_15s
    'h1b1e: romdata_int = 'h7b;
    'h1b1f: romdata_int = 'h11e;
    'h1b20: romdata_int = 'h2df;
    'h1b21: romdata_int = 'h400;
    'h1b22: romdata_int = 'h91f;
    'h1b23: romdata_int = 'h1936;
    'h1b24: romdata_int = 'h1a97;
    'h1b25: romdata_int = 'h1c00;
    'h1b26: romdata_int = 'h2e3b;
    'h1b27: romdata_int = 'h3400;
    'h1b28: romdata_int = 'h38c8;
    'h1b29: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b2a: romdata_int = 'h10a;
    'h1b2b: romdata_int = 'h600;
    'h1b2c: romdata_int = 'hce4;
    'h1b2d: romdata_int = 'h1279;
    'h1b2e: romdata_int = 'h1e00;
    'h1b2f: romdata_int = 'h26ba;
    'h1b30: romdata_int = 'h345c;
    'h1b31: romdata_int = 'h3600;
    'h1b32: romdata_int = 'h3c0e;
    'h1b33: romdata_int = 'h490c; // Line descriptor for 11_15s
    'h1b34: romdata_int = 'h15e;
    'h1b35: romdata_int = 'h54f;
    'h1b36: romdata_int = 'h800;
    'h1b37: romdata_int = 'h10ba;
    'h1b38: romdata_int = 'h12fc;
    'h1b39: romdata_int = 'h2000;
    'h1b3a: romdata_int = 'h2254;
    'h1b3b: romdata_int = 'h2b00;
    'h1b3c: romdata_int = 'h32c1;
    'h1b3d: romdata_int = 'h3800;
    'h1b3e: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b3f: romdata_int = 'ha00;
    'h1b40: romdata_int = 'haab;
    'h1b41: romdata_int = 'hd5c;
    'h1b42: romdata_int = 'h146e;
    'h1b43: romdata_int = 'h1f2e;
    'h1b44: romdata_int = 'h2200;
    'h1b45: romdata_int = 'h2ace;
    'h1b46: romdata_int = 'h2c5a;
    'h1b47: romdata_int = 'h3a00;
    'h1b48: romdata_int = 'h470c; // Line descriptor for 11_15s
    'h1b49: romdata_int = 'h6db;
    'h1b4a: romdata_int = 'hc00;
    'h1b4b: romdata_int = 'h165e;
    'h1b4c: romdata_int = 'h1e68;
    'h1b4d: romdata_int = 'h2400;
    'h1b4e: romdata_int = 'h2cfb;
    'h1b4f: romdata_int = 'h3a9c;
    'h1b50: romdata_int = 'h3c00;
    'h1b51: romdata_int = 'h80c; // Line descriptor for 11_15s
    'h1b52: romdata_int = 'h27;
    'h1b53: romdata_int = 'he00;
    'h1b54: romdata_int = 'hf48;
    'h1b55: romdata_int = 'h1c93;
    'h1b56: romdata_int = 'h2133;
    'h1b57: romdata_int = 'h2600;
    'h1b58: romdata_int = 'h360b;
    'h1b59: romdata_int = 'h388c;
    'h1b5a: romdata_int = 'h3e00;
    'h1b5b: romdata_int = 'h690c; // Line descriptor for 11_15s
    'h1b5c: romdata_int = 'h38;
    'h1b5d: romdata_int = 'h2b1;
    'h1b5e: romdata_int = 'h502;
    'h1b5f: romdata_int = 'h1000;
    'h1b60: romdata_int = 'h2652;
    'h1b61: romdata_int = 'h2800;
    'h1b62: romdata_int = 'h289e;
    'h1b63: romdata_int = 'h2e72;
    'h1b64: romdata_int = 'h4000;
    'h1b65: romdata_int = 'h4075;
    'h1b66: romdata_int = 'h90a; // Line descriptor for 7_9s
    'h1b67: romdata_int = 'h541;
    'h1b68: romdata_int = 'ha00;
    'h1b69: romdata_int = 'hc17;
    'h1b6a: romdata_int = 'h14d3;
    'h1b6b: romdata_int = 'h1e00;
    'h1b6c: romdata_int = 'h20b4;
    'h1b6d: romdata_int = 'h2148;
    'h1b6e: romdata_int = 'h3200;
    'h1b6f: romdata_int = 'h36a1;
    'h1b70: romdata_int = 'h3f5a;
    'h1b71: romdata_int = 'h480a; // Line descriptor for 7_9s
    'h1b72: romdata_int = 'hc00;
    'h1b73: romdata_int = 'h185f;
    'h1b74: romdata_int = 'h1c8e;
    'h1b75: romdata_int = 'h2000;
    'h1b76: romdata_int = 'h2221;
    'h1b77: romdata_int = 'h2c0c;
    'h1b78: romdata_int = 'h3400;
    'h1b79: romdata_int = 'h34bc;
    'h1b7a: romdata_int = 'h370e;
    'h1b7b: romdata_int = 'ha0a; // Line descriptor for 7_9s
    'h1b7c: romdata_int = 'h415;
    'h1b7d: romdata_int = 'h83d;
    'h1b7e: romdata_int = 'he00;
    'h1b7f: romdata_int = 'h1256;
    'h1b80: romdata_int = 'h1b62;
    'h1b81: romdata_int = 'h1ee3;
    'h1b82: romdata_int = 'h2200;
    'h1b83: romdata_int = 'h24ff;
    'h1b84: romdata_int = 'h3248;
    'h1b85: romdata_int = 'h3600;
    'h1b86: romdata_int = 'h38ad;
    'h1b87: romdata_int = 'h490a; // Line descriptor for 7_9s
    'h1b88: romdata_int = 'h2f9;
    'h1b89: romdata_int = 'hb0a;
    'h1b8a: romdata_int = 'h1000;
    'h1b8b: romdata_int = 'h101c;
    'h1b8c: romdata_int = 'h2400;
    'h1b8d: romdata_int = 'h2822;
    'h1b8e: romdata_int = 'h288a;
    'h1b8f: romdata_int = 'h3800;
    'h1b90: romdata_int = 'h3948;
    'h1b91: romdata_int = 'h3c18;
    'h1b92: romdata_int = 'h90a; // Line descriptor for 7_9s
    'h1b93: romdata_int = 'h212;
    'h1b94: romdata_int = 'hf17;
    'h1b95: romdata_int = 'h1200;
    'h1b96: romdata_int = 'h16cb;
    'h1b97: romdata_int = 'h2600;
    'h1b98: romdata_int = 'h2a09;
    'h1b99: romdata_int = 'h2f15;
    'h1b9a: romdata_int = 'h329e;
    'h1b9b: romdata_int = 'h3a00;
    'h1b9c: romdata_int = 'h3d33;
    'h1b9d: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1b9e: romdata_int = 'h0;
    'h1b9f: romdata_int = 'h9c;
    'h1ba0: romdata_int = 'hd0d;
    'h1ba1: romdata_int = 'heca;
    'h1ba2: romdata_int = 'h1400;
    'h1ba3: romdata_int = 'h242e;
    'h1ba4: romdata_int = 'h2800;
    'h1ba5: romdata_int = 'h30b9;
    'h1ba6: romdata_int = 'h3c00;
    'h1ba7: romdata_int = 'h3e5e;
    'h1ba8: romdata_int = 'h4562;
    'h1ba9: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1baa: romdata_int = 'h59;
    'h1bab: romdata_int = 'h200;
    'h1bac: romdata_int = 'h1425;
    'h1bad: romdata_int = 'h1600;
    'h1bae: romdata_int = 'h16e4;
    'h1baf: romdata_int = 'h2a00;
    'h1bb0: romdata_int = 'h2a17;
    'h1bb1: romdata_int = 'h30d3;
    'h1bb2: romdata_int = 'h3e00;
    'h1bb3: romdata_int = 'h40ae;
    'h1bb4: romdata_int = 'h4238;
    'h1bb5: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1bb6: romdata_int = 'h400;
    'h1bb7: romdata_int = 'h648;
    'h1bb8: romdata_int = 'hac2;
    'h1bb9: romdata_int = 'h1800;
    'h1bba: romdata_int = 'h1c1e;
    'h1bbb: romdata_int = 'h1e77;
    'h1bbc: romdata_int = 'h2c00;
    'h1bbd: romdata_int = 'h2e95;
    'h1bbe: romdata_int = 'h3514;
    'h1bbf: romdata_int = 'h4000;
    'h1bc0: romdata_int = 'h428e;
    'h1bc1: romdata_int = 'h4a0a; // Line descriptor for 7_9s
    'h1bc2: romdata_int = 'h600;
    'h1bc3: romdata_int = 'h956;
    'h1bc4: romdata_int = 'h18ce;
    'h1bc5: romdata_int = 'h1a00;
    'h1bc6: romdata_int = 'h1b36;
    'h1bc7: romdata_int = 'h22e6;
    'h1bc8: romdata_int = 'h2667;
    'h1bc9: romdata_int = 'h2e00;
    'h1bca: romdata_int = 'h3a10;
    'h1bcb: romdata_int = 'h4200;
    'h1bcc: romdata_int = 'h4474;
    'h1bcd: romdata_int = 'h6a0a; // Line descriptor for 7_9s
    'h1bce: romdata_int = 'h685;
    'h1bcf: romdata_int = 'h800;
    'h1bd0: romdata_int = 'h112f;
    'h1bd1: romdata_int = 'h1320;
    'h1bd2: romdata_int = 'h1c00;
    'h1bd3: romdata_int = 'h26f7;
    'h1bd4: romdata_int = 'h2d05;
    'h1bd5: romdata_int = 'h3000;
    'h1bd6: romdata_int = 'h3a6d;
    'h1bd7: romdata_int = 'h40cc;
    'h1bd8: romdata_int = 'h4400;
    'h1bd9: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1bda: romdata_int = 'h11b;
    'h1bdb: romdata_int = 'h499;
    'h1bdc: romdata_int = 'ha00;
    'h1bdd: romdata_int = 'hb08;
    'h1bde: romdata_int = 'h109e;
    'h1bdf: romdata_int = 'h1a00;
    'h1be0: romdata_int = 'h1e8a;
    'h1be1: romdata_int = 'h1ed4;
    'h1be2: romdata_int = 'h2a00;
    'h1be3: romdata_int = 'h2a20;
    'h1be4: romdata_int = 'h3522;
    'h1be5: romdata_int = 'h3a00;
    'h1be6: romdata_int = 'h452b;
    'h1be7: romdata_int = 'h48d5;
    'h1be8: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1be9: romdata_int = 'hb9;
    'h1bea: romdata_int = 'h12d;
    'h1beb: romdata_int = 'hc00;
    'h1bec: romdata_int = 'he44;
    'h1bed: romdata_int = 'h180a;
    'h1bee: romdata_int = 'h1c00;
    'h1bef: romdata_int = 'h1c15;
    'h1bf0: romdata_int = 'h263e;
    'h1bf1: romdata_int = 'h2c00;
    'h1bf2: romdata_int = 'h2e9d;
    'h1bf3: romdata_int = 'h3099;
    'h1bf4: romdata_int = 'h3b28;
    'h1bf5: romdata_int = 'h3c00;
    'h1bf6: romdata_int = 'h3c07;
    'h1bf7: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1bf8: romdata_int = 'h669;
    'h1bf9: romdata_int = 'h708;
    'h1bfa: romdata_int = 'he00;
    'h1bfb: romdata_int = 'h131a;
    'h1bfc: romdata_int = 'h160e;
    'h1bfd: romdata_int = 'h1e00;
    'h1bfe: romdata_int = 'h20ef;
    'h1bff: romdata_int = 'h22b5;
    'h1c00: romdata_int = 'h2b36;
    'h1c01: romdata_int = 'h2e00;
    'h1c02: romdata_int = 'h2ecf;
    'h1c03: romdata_int = 'h3e00;
    'h1c04: romdata_int = 'h3e83;
    'h1c05: romdata_int = 'h42d9;
    'h1c06: romdata_int = 'h4d08; // Line descriptor for 37_45s
    'h1c07: romdata_int = 'h0;
    'h1c08: romdata_int = 'h3e;
    'h1c09: romdata_int = 'he66;
    'h1c0a: romdata_int = 'h1000;
    'h1c0b: romdata_int = 'h1918;
    'h1c0c: romdata_int = 'h2000;
    'h1c0d: romdata_int = 'h240b;
    'h1c0e: romdata_int = 'h28c5;
    'h1c0f: romdata_int = 'h3000;
    'h1c10: romdata_int = 'h354e;
    'h1c11: romdata_int = 'h3636;
    'h1c12: romdata_int = 'h3c3c;
    'h1c13: romdata_int = 'h4000;
    'h1c14: romdata_int = 'h4614;
    'h1c15: romdata_int = 'h5008; // Line descriptor for 37_45s
    'h1c16: romdata_int = 'h71;
    'h1c17: romdata_int = 'h59;
    'h1c18: romdata_int = 'h139;
    'h1c19: romdata_int = 'h200;
    'h1c1a: romdata_int = 'h81a;
    'h1c1b: romdata_int = 'hd25;
    'h1c1c: romdata_int = 'h1200;
    'h1c1d: romdata_int = 'h1478;
    'h1c1e: romdata_int = 'h2200;
    'h1c1f: romdata_int = 'h2242;
    'h1c20: romdata_int = 'h2716;
    'h1c21: romdata_int = 'h3200;
    'h1c22: romdata_int = 'h327a;
    'h1c23: romdata_int = 'h381c;
    'h1c24: romdata_int = 'h4200;
    'h1c25: romdata_int = 'h4208;
    'h1c26: romdata_int = 'h494a;
    'h1c27: romdata_int = 'h4f08; // Line descriptor for 37_45s
    'h1c28: romdata_int = 'h29;
    'h1c29: romdata_int = 'h15e;
    'h1c2a: romdata_int = 'h400;
    'h1c2b: romdata_int = 'h847;
    'h1c2c: romdata_int = 'h12d4;
    'h1c2d: romdata_int = 'h1400;
    'h1c2e: romdata_int = 'h172d;
    'h1c2f: romdata_int = 'h1a9b;
    'h1c30: romdata_int = 'h1ac5;
    'h1c31: romdata_int = 'h2400;
    'h1c32: romdata_int = 'h2c8b;
    'h1c33: romdata_int = 'h2c9d;
    'h1c34: romdata_int = 'h3400;
    'h1c35: romdata_int = 'h3aeb;
    'h1c36: romdata_int = 'h4400;
    'h1c37: romdata_int = 'h4650;
    'h1c38: romdata_int = 'h5008; // Line descriptor for 37_45s
    'h1c39: romdata_int = 'h9e;
    'h1c3a: romdata_int = 'hd4;
    'h1c3b: romdata_int = 'h2f0;
    'h1c3c: romdata_int = 'h433;
    'h1c3d: romdata_int = 'h600;
    'h1c3e: romdata_int = 'hd1d;
    'h1c3f: romdata_int = 'h1414;
    'h1c40: romdata_int = 'h1600;
    'h1c41: romdata_int = 'h2479;
    'h1c42: romdata_int = 'h2600;
    'h1c43: romdata_int = 'h2922;
    'h1c44: romdata_int = 'h30b8;
    'h1c45: romdata_int = 'h3600;
    'h1c46: romdata_int = 'h369f;
    'h1c47: romdata_int = 'h3e68;
    'h1c48: romdata_int = 'h40f8;
    'h1c49: romdata_int = 'h4600;
    'h1c4a: romdata_int = 'h6e08; // Line descriptor for 37_45s
    'h1c4b: romdata_int = 'h45;
    'h1c4c: romdata_int = 'h331;
    'h1c4d: romdata_int = 'h800;
    'h1c4e: romdata_int = 'hb29;
    'h1c4f: romdata_int = 'h1011;
    'h1c50: romdata_int = 'h1800;
    'h1c51: romdata_int = 'h1c60;
    'h1c52: romdata_int = 'h2161;
    'h1c53: romdata_int = 'h2800;
    'h1c54: romdata_int = 'h3339;
    'h1c55: romdata_int = 'h3800;
    'h1c56: romdata_int = 'h383e;
    'h1c57: romdata_int = 'h4099;
    'h1c58: romdata_int = 'h4476;
    'h1c59: romdata_int = 'h4800;
    'h1c5a: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c5b: romdata_int = 'h0;
    'h1c5c: romdata_int = 'ha1;
    'h1c5d: romdata_int = 'h322;
    'h1c5e: romdata_int = 'h879;
    'h1c5f: romdata_int = 'ha00;
    'h1c60: romdata_int = 'h102a;
    'h1c61: romdata_int = 'h10ef;
    'h1c62: romdata_int = 'h1400;
    'h1c63: romdata_int = 'h1aa7;
    'h1c64: romdata_int = 'h1b2c;
    'h1c65: romdata_int = 'h1e00;
    'h1c66: romdata_int = 'h20e7;
    'h1c67: romdata_int = 'h272b;
    'h1c68: romdata_int = 'h2800;
    'h1c69: romdata_int = 'h284d;
    'h1c6a: romdata_int = 'h2ec0;
    'h1c6b: romdata_int = 'h3200;
    'h1c6c: romdata_int = 'h34cb;
    'h1c6d: romdata_int = 'h38ee;
    'h1c6e: romdata_int = 'h3c00;
    'h1c6f: romdata_int = 'h3c7e;
    'h1c70: romdata_int = 'h44e7;
    'h1c71: romdata_int = 'h4600;
    'h1c72: romdata_int = 'h46c8;
    'h1c73: romdata_int = 'h4d2f;
    'h1c74: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c75: romdata_int = 'h200;
    'h1c76: romdata_int = 'h55c;
    'h1c77: romdata_int = 'h6a1;
    'h1c78: romdata_int = 'h739;
    'h1c79: romdata_int = 'hab9;
    'h1c7a: romdata_int = 'hc00;
    'h1c7b: romdata_int = 'he1e;
    'h1c7c: romdata_int = 'h1600;
    'h1c7d: romdata_int = 'h1911;
    'h1c7e: romdata_int = 'h1d2b;
    'h1c7f: romdata_int = 'h1ec9;
    'h1c80: romdata_int = 'h1f54;
    'h1c81: romdata_int = 'h2000;
    'h1c82: romdata_int = 'h2a00;
    'h1c83: romdata_int = 'h2a1e;
    'h1c84: romdata_int = 'h3122;
    'h1c85: romdata_int = 'h3400;
    'h1c86: romdata_int = 'h36fc;
    'h1c87: romdata_int = 'h3af9;
    'h1c88: romdata_int = 'h3e00;
    'h1c89: romdata_int = 'h3e54;
    'h1c8a: romdata_int = 'h446f;
    'h1c8b: romdata_int = 'h467e;
    'h1c8c: romdata_int = 'h4800;
    'h1c8d: romdata_int = 'h4c65;
    'h1c8e: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1c8f: romdata_int = 'h8e;
    'h1c90: romdata_int = 'h30b;
    'h1c91: romdata_int = 'h400;
    'h1c92: romdata_int = 'h860;
    'h1c93: romdata_int = 'hc9b;
    'h1c94: romdata_int = 'he00;
    'h1c95: romdata_int = 'h128a;
    'h1c96: romdata_int = 'h1455;
    'h1c97: romdata_int = 'h1800;
    'h1c98: romdata_int = 'h1c64;
    'h1c99: romdata_int = 'h2013;
    'h1c9a: romdata_int = 'h2200;
    'h1c9b: romdata_int = 'h2283;
    'h1c9c: romdata_int = 'h2a49;
    'h1c9d: romdata_int = 'h2c00;
    'h1c9e: romdata_int = 'h2c28;
    'h1c9f: romdata_int = 'h3358;
    'h1ca0: romdata_int = 'h3600;
    'h1ca1: romdata_int = 'h3b26;
    'h1ca2: romdata_int = 'h4000;
    'h1ca3: romdata_int = 'h424e;
    'h1ca4: romdata_int = 'h4273;
    'h1ca5: romdata_int = 'h4892;
    'h1ca6: romdata_int = 'h4a00;
    'h1ca7: romdata_int = 'h4eea;
    'h1ca8: romdata_int = 'h5805; // Line descriptor for 8_9s
    'h1ca9: romdata_int = 'h137;
    'h1caa: romdata_int = 'h2ae;
    'h1cab: romdata_int = 'h600;
    'h1cac: romdata_int = 'h8b8;
    'h1cad: romdata_int = 'hb3b;
    'h1cae: romdata_int = 'he79;
    'h1caf: romdata_int = 'h1000;
    'h1cb0: romdata_int = 'h1461;
    'h1cb1: romdata_int = 'h16a5;
    'h1cb2: romdata_int = 'h1a00;
    'h1cb3: romdata_int = 'h2318;
    'h1cb4: romdata_int = 'h2400;
    'h1cb5: romdata_int = 'h2522;
    'h1cb6: romdata_int = 'h2d08;
    'h1cb7: romdata_int = 'h2e00;
    'h1cb8: romdata_int = 'h2e3f;
    'h1cb9: romdata_int = 'h32db;
    'h1cba: romdata_int = 'h351d;
    'h1cbb: romdata_int = 'h3800;
    'h1cbc: romdata_int = 'h3c65;
    'h1cbd: romdata_int = 'h40b3;
    'h1cbe: romdata_int = 'h4200;
    'h1cbf: romdata_int = 'h4911;
    'h1cc0: romdata_int = 'h4b09;
    'h1cc1: romdata_int = 'h4c00;
    'h1cc2: romdata_int = 'h7805; // Line descriptor for 8_9s
    'h1cc3: romdata_int = 'h4e1;
    'h1cc4: romdata_int = 'h4ec;
    'h1cc5: romdata_int = 'h63a;
    'h1cc6: romdata_int = 'h800;
    'h1cc7: romdata_int = 'hd12;
    'h1cc8: romdata_int = 'h1200;
    'h1cc9: romdata_int = 'h1328;
    'h1cca: romdata_int = 'h16e0;
    'h1ccb: romdata_int = 'h18ae;
    'h1ccc: romdata_int = 'h1c00;
    'h1ccd: romdata_int = 'h247c;
    'h1cce: romdata_int = 'h2600;
    'h1ccf: romdata_int = 'h2655;
    'h1cd0: romdata_int = 'h28a1;
    'h1cd1: romdata_int = 'h3000;
    'h1cd2: romdata_int = 'h30cf;
    'h1cd3: romdata_int = 'h3738;
    'h1cd4: romdata_int = 'h386c;
    'h1cd5: romdata_int = 'h3a00;
    'h1cd6: romdata_int = 'h3f54;
    'h1cd7: romdata_int = 'h4038;
    'h1cd8: romdata_int = 'h4400;
    'h1cd9: romdata_int = 'h4a41;
    'h1cda: romdata_int = 'h4e00;
    default: romdata_int = 'h4edc;
  endcase
endmodule

