library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
Library UNISIM;
use UNISIM.vcomponents.all;

entity ucecho is
   port(
      pd        : in unsigned(7 downto 0);
      pb        : out unsigned(7 downto 0);
      fxclk_in  : in std_logic
   );
end ucecho;


architecture RTL of ucecho is

--signal declaration
signal pb_buf : unsigned(7 downto 0);
signal clk : std_logic;
signal fxclk_fb : std_logic;

begin
    -- PLL used as clock filter
    fxclk_pll : PLLE2_BASE
    generic map (
       BANDWIDTH => "OPTIMIZED",  -- OPTIMIZED, HIGH, LOW
       CLKFBOUT_MULT => 20,       -- Multiply value for all CLKOUT, (2-64)
       CLKFBOUT_PHASE => 0.0,     -- Phase offset in degrees of CLKFB, (-360.000-360.000).
       CLKIN1_PERIOD => 0.0,      -- Input clock period in ns to ps resolution (i.e. 33.333 is 30 MHz).
       -- CLKOUT0_DIVIDE - CLKOUT5_DIVIDE: Divide amount for each CLKOUT (1-128)
       CLKOUT0_DIVIDE => 10,
       CLKOUT1_DIVIDE => 1,
       CLKOUT2_DIVIDE => 1,
       CLKOUT3_DIVIDE => 1,
       CLKOUT4_DIVIDE => 1,
       CLKOUT5_DIVIDE => 1,
       -- CLKOUT0_DUTY_CYCLE - CLKOUT5_DUTY_CYCLE: Duty cycle for each CLKOUT (0.001-0.999).
       CLKOUT0_DUTY_CYCLE => 0.5,
       CLKOUT1_DUTY_CYCLE => 0.5,
       CLKOUT2_DUTY_CYCLE => 0.5,
       CLKOUT3_DUTY_CYCLE => 0.5,
       CLKOUT4_DUTY_CYCLE => 0.5,
       CLKOUT5_DUTY_CYCLE => 0.5,
       -- CLKOUT0_PHASE - CLKOUT5_PHASE: Phase offset for each CLKOUT (-360.000-360.000).
       CLKOUT0_PHASE => 0.0,
       CLKOUT1_PHASE => 0.0,
       CLKOUT2_PHASE => 0.0,
       CLKOUT3_PHASE => 0.0,
       CLKOUT4_PHASE => 0.0,
       CLKOUT5_PHASE => 0.0,
       DIVCLK_DIVIDE => 1,        -- Master division value, (1-56)
       REF_JITTER1 => 0.0,        -- Reference input jitter in UI, (0.000-0.999).
       STARTUP_WAIT => "FALSE"    -- Delay DONE until PLL Locks, ("TRUE"/"FALSE")
    )
    port map (
       CLKOUT0 => clk,
       CLKFBOUT => fxclk_fb,   -- 1-bit output: Feedback clock
       CLKIN1 => fxclk_in,     -- 1-bit input: Input clock
       PWRDWN => '0',          -- 1-bit input: Power-down
       RST => '0',             -- 1-bit input: Reset
       CLKFBIN => fxclk_fb     -- 1-bit input: Feedback clock
    );

    dpUCECHO: process(CLK)
    begin
         if CLK' event and CLK = '1' then
	    if ( pd >= 97 ) and ( pd <= 122)
	    then
		pb_buf <= pd - 32;
	    else
		pb_buf <= pd;
	    end if;
	    pb <= pb_buf;
	end if;
    end process dpUCECHO;
    
end RTL;
