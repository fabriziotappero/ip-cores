-------------------------------------------------------------------------------
--
-- Generic testbench elements
--
-- $Id: tb_elems-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration tb_elems_behav_c0 of tb_elems is

  for behav
  end for;

end tb_elems_behav_c0;
