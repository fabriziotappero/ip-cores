/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

module rom (clk, addr, out);
   input clk;
   input [8:0] addr;
   output reg [27:0] out;
   
   always @(posedge clk)
      case (addr)
         0: out <= 28'hc30042;
         1: out <= 28'h1450045;
         2: out <= 28'h1868041;
         3: out <= 28'h1c78041;
         4: out <= 28'h30046;
         5: out <= 28'h580ea00;
         6: out <= 28'h5c08041;
         7: out <= 28'h5c5ea17;
         8: out <= 28'h605ea07;
         9: out <= 28'h658ea07;
         10: out <= 28'h3d74059;
         11: out <= 28'h3c5404f;
         12: out <= 28'h5d8ea05;
         13: out <= 28'h617ea00;
         14: out <= 28'h587ea16;
         15: out <= 28'h4580056;
         16: out <= 28'h4850041;
         17: out <= 28'h4c7ea00;
         18: out <= 28'h4d34057;
         19: out <= 28'h5014041;
         20: out <= 28'h5474041;
         21: out <= 28'hf8041;
         22: out <= 28'h5918041;
         23: out <= 28'h5d28041;
         24: out <= 28'h6138041;
         25: out <= 28'h6548041;
         26: out <= 28'h6958041;
         27: out <= 28'h3c00057;
         28: out <= 28'h3cf0059;
         29: out <= 28'h4560058;
         30: out <= 28'h451005a;
         31: out <= 28'h4510051;
         32: out <= 28'h4974059;
         33: out <= 28'h4da4058;
         34: out <= 28'h5190041;
         35: out <= 28'h55a005a;
         36: out <= 28'h1868081;
         37: out <= 28'h1864042;
         38: out <= 28'h1c78081;
         39: out <= 28'h1c70047;
         40: out <= 28'h30046;
         41: out <= 28'h5800040;
         42: out <= 28'h5c5ea07;
         43: out <= 28'h16ea00;
         44: out <= 28'h6000056;
         45: out <= 28'h6404056;
         46: out <= 28'h68f0054;
         47: out <= 28'h6da0052;
         48: out <= 28'h71a4052;
         49: out <= 28'h74f4054;
         50: out <= 28'h79d4053;
         51: out <= 28'h75d0053;
         52: out <= 28'h7d10055;
         53: out <= 28'h81f0053;
         54: out <= 28'h85f4053;
         55: out <= 28'h8970056;
         56: out <= 28'h5974056;
         57: out <= 28'h8d14055;
         58: out <= 28'h9230052;
         59: out <= 28'h8e34052;
         60: out <= 28'h9580057;
         61: out <= 28'h99b0060;
         62: out <= 28'h9c00062;
         63: out <= 28'ha1e0064;
         64: out <= 28'ha590057;
         65: out <= 28'ha9c0061;
         66: out <= 28'hac00056;
         67: out <= 28'hb1d0063;
         68: out <= 28'h618ea1b;
         69: out <= 28'h6e5ea26;
         70: out <= 28'h817ea20;
         71: out <= 28'h780ea1e;
         72: out <= 28'h967ea28;
         73: out <= 28'h8a2ea24;
         74: out <= 28'h659ea1c;
         75: out <= 28'h729ea2a;
         76: out <= 28'h5d7ea21;
         77: out <= 28'hea1d;
         78: out <= 28'h76bea2c;
         79: out <= 28'h596ea23;
         80: out <= 28'h8580065;
         81: out <= 28'h8e0005d;
         82: out <= 28'h9204057;
         83: out <= 28'h9994058;
         84: out <= 28'h5d70060;
         85: out <= 28'h5e24057;
         86: out <= 28'h5d70056;
         87: out <= 28'h6190058;
         88: out <= 28'h618405e;
         89: out <= 28'h6184040;
         90: out <= 28'h6634061;
         91: out <= 28'h659405e;
         92: out <= 28'h5990056;
         93: out <= 28'h6610063;
         94: out <= 28'h659405b;
         95: out <= 28'h6590062;
         96: out <= 28'h190040;
         97: out <= 28'h6640066;
         98: out <= 28'h7a44066;
         99: out <= 28'h79e005c;
         100: out <= 28'h79e405b;
         101: out <= 28'h8170058;
         102: out <= 28'h5d74058;
         103: out <= 28'h5d7005c;
         104: out <= 28'h5d7005b;
         105: out <= 28'h5d74065;
         106: out <= 28'h5d7405d;
         107: out <= 28'h3d64052;
         108: out <= 28'h4404053;
         109: out <= 28'h194052;
         110: out <= 28'h4054;
         111: out <= 28'h59e4053;
         112: out <= 28'h5964055;
         113: out <= 28'h520405a;
         114: out <= 28'h557405f;
         115: out <= 28'h4804041;
         116: out <= 28'h4d64041;
         117: out <= 28'h24f8041;
         118: out <= 28'hf0052;
         119: out <= 28'h54;
         120: out <= 28'h58fea0f;
         121: out <= 28'h5cfea12;
         122: out <= 28'h612ea14;
         123: out <= 28'h654ea14;
         124: out <= 28'hea00;
         125: out <= 28'h5d70058;
         126: out <= 28'h6164058;
         127: out <= 28'h6594057;
         128: out <= 28'h57;
         129: out <= 28'h4056;
         130: out <= 28'h5910053;
         131: out <= 28'h5960055;
         132: out <= 28'h5d1ea11;
         133: out <= 28'h691ea13;
         134: out <= 28'h6d3ea15;
         135: out <= 28'h715ea15;
         136: out <= 28'h596ea16;
         137: out <= 28'h69a005b;
         138: out <= 28'h6d7405b;
         139: out <= 28'h71c405a;
         140: out <= 28'h596005a;
         141: out <= 28'h5964057;
         142: out <= 28'h5cf0052;
         143: out <= 28'h68f0054;
         144: out <= 28'h7520054;
         145: out <= 28'h7910053;
         146: out <= 28'h7d10055;
         147: out <= 28'h8130055;
         148: out <= 28'h84fea11;
         149: out <= 28'h892ea13;
         150: out <= 28'h8d4ea15;
         151: out <= 28'h5d7ea1e;
         152: out <= 28'h69aea1f;
         153: out <= 28'h75dea20;
         154: out <= 28'h7a14062;
         155: out <= 28'h7de4063;
         156: out <= 28'h7df005d;
         157: out <= 28'h5d7405e;
         158: out <= 28'h5d7005d;
         159: out <= 28'h69a405e;
         160: out <= 28'h758405b;
         161: out <= 28'h799405c;
         162: out <= 28'h8004056;
         163: out <= 28'h618005b;
         164: out <= 28'h659005c;
         165: out <= 28'h56;
         166: out <= 28'h5980059;
         167: out <= 28'h6d84040;
         168: out <= 28'h7194058;
         169: out <= 28'h840405c;
         170: out <= 28'h898ea18;
         171: out <= 28'h8d9ea19;
         172: out <= 28'h900ea00;
         173: out <= 28'h658ea19;
         174: out <= 28'h618ea00;
         175: out <= 28'hea16;
         176: out <= 28'h5a2ea1b;
         177: out <= 28'h6e3ea1c;
         178: out <= 28'h724ea21;
         179: out <= 28'h596005b;
         180: out <= 28'h596005c;
         181: out <= 28'h6d60041;
         182: out <= 28'h71b8041;
         183: out <= 28'h71bea1c;
         184: out <= 28'h71c8041;
         185: out <= 28'h71bea1c;
         186: out <= 28'h85c8041;
         187: out <= 28'h6dbea21;
         188: out <= 28'h85b80c1;
         189: out <= 28'h71cea21;
         190: out <= 28'h71c8101;
         191: out <= 28'h71bea1c;
         192: out <= 28'h85c8101;
         193: out <= 28'h6dbea21;
         194: out <= 28'h85b83c1;
         195: out <= 28'h6dbea21;
         196: out <= 28'h85b8781;
         197: out <= 28'h6dbea21;
         198: out <= 28'h85b8f01;
         199: out <= 28'h6dbea21;
         200: out <= 28'h85b82c1;
         201: out <= 28'h71cea21;
         202: out <= 28'h71c9e01;
         203: out <= 28'h6dbea1c;
         204: out <= 28'h71bbec1;
         205: out <= 28'h6dbea1c;
         206: out <= 28'h6db8041;
         207: out <= 28'h59bea16;
         208: out <= 28'h59bea16;
         209: out <= 28'h6e34064;
         210: out <= 28'h722405b;
         211: out <= 28'h1c4040;
         212: out <= 28'h6644059;
         213: out <= 28'h61b4058;
         214: out <= 28'h16ea00;
         215: out <= 28'h656ea19;
         216: out <= 28'h596ea18;
         217: out <= 28'h61d005e;
         218: out <= 28'h6dd0060;
         219: out <= 28'h71e0060;
         220: out <= 28'h8400059;
         221: out <= 28'h8800056;
         222: out <= 28'h8d90056;
         223: out <= 28'h75dea00;
         224: out <= 28'h79eea19;
         225: out <= 28'h820ea16;
         226: out <= 28'h618ea21;
         227: out <= 28'h6dbea22;
         228: out <= 28'h71cea23;
         229: out <= 28'h75d405e;
         230: out <= 28'h79d4060;
         231: out <= 28'h79e005c;
         232: out <= 28'h618405d;
         233: out <= 28'h618005c;
         234: out <= 28'h6db405d;
         235: out <= 28'h71f0057;
         236: out <= 28'h75f005a;
         237: out <= 28'h817005a;
         238: out <= 28'h8400059;
         239: out <= 28'h8800056;
         240: out <= 28'h8d90056;
         241: out <= 28'h1fea00;
         242: out <= 28'h5d7ea19;
         243: out <= 28'h59aea16;
         244: out <= 28'h65cea21;
         245: out <= 28'h69dea22;
         246: out <= 28'h720ea23;
         247: out <= 28'h4057;
         248: out <= 28'h5804056;
         249: out <= 28'h596005c;
         250: out <= 28'h5d94040;
         251: out <= 28'h5d7005c;
         252: out <= 28'h1a4040;
         253: out <= 28'h65e0056;
         254: out <= 28'h6980057;
         255: out <= 28'h71b4040;
         256: out <= 28'h75eea1b;
         257: out <= 28'h7d6ea00;
         258: out <= 28'h6d8ea1b;
         259: out <= 28'h17ea00;
         260: out <= 28'h819ea1c;
         261: out <= 28'h596ea18;
         262: out <= 28'h5deea17;
         263: out <= 28'h619ea1a;
         264: out <= 28'h65aea1c;
         265: out <= 28'h6960057;
         266: out <= 28'h61a4058;
         267: out <= 28'h69b0040;
         268: out <= 28'h69a005a;
         269: out <= 28'h405b;
         270: out <= 28'h6df405d;
         271: out <= 28'h6db0060;
         272: out <= 28'h702005d;
         273: out <= 28'h71c005f;
         274: out <= 28'h71c405a;
         275: out <= 28'h5974056;
         276: out <= 28'h59b0056;
         277: out <= 28'h5d80041;
         278: out <= 28'h7590040;
         279: out <= 28'h6dd005b;
         280: out <= 28'h618005a;
         281: out <= 28'h6180058;
         282: out <= 28'h190040;
         283: out <= 28'h40;
         284: out <= 28'h65c8041;
         285: out <= 28'h6968041;
         286: out <= 28'h7578041;
         287: out <= 28'h79b8041;
         288: out <= 28'h7d88041;
         289: out <= 28'h8008041;
         290: out <= 28'h659005d;
         291: out <= 28'h659005f;
         292: out <= 28'h69a005a;
         293: out <= 28'h69a405e;
         294: out <= 28'h69a4060;
         295: out <= 28'h75d405f;
         296: out <= 28'h7a0405e;
         297: out <= 28'h8200060;
         298: out <= 28'h6598041;
         299: out <= 28'h69a8041;
         300: out <= 28'h75d8041;
         301: out <= 28'h79e8041;
         302: out <= 28'h7df8041;
         303: out <= 28'h8208041;
         304: out <= 28'h659005d;
         305: out <= 28'h659005f;
         306: out <= 28'h69a005a;
         307: out <= 28'h69a405e;
         308: out <= 28'h69a4060;
         309: out <= 28'h75d405f;
         310: out <= 28'h7a0405e;
         311: out <= 28'h8200060;
         312: out <= 28'h85c0056;
         313: out <= 28'h897005b;
         314: out <= 28'h8d84040;
         315: out <= 28'h91cea18;
         316: out <= 28'h956ea00;
         317: out <= 28'h617ea18;
         318: out <= 28'h1bea00;
         319: out <= 28'h9a1ea23;
         320: out <= 28'h596ea17;
         321: out <= 28'h5dcea1b;
         322: out <= 28'h6e1ea22;
         323: out <= 28'h722ea23;
         324: out <= 28'h8560057;
         325: out <= 28'h6e1405b;
         326: out <= 28'h8580040;
         327: out <= 28'h8610061;
         328: out <= 28'h4058;
         329: out <= 28'h6254064;
         330: out <= 28'h6180066;
         331: out <= 28'h8820064;
         332: out <= 28'h8a20065;
         333: out <= 28'h8a24061;
         334: out <= 28'h5974056;
         335: out <= 28'h5980056;
         336: out <= 28'h5db0041;
         337: out <= 28'h8dc0040;
         338: out <= 28'h6230058;
         339: out <= 28'h6db0061;
         340: out <= 28'h6db005b;
         341: out <= 28'h1c0040;
         342: out <= 28'h40;
         343: out <= 28'h69a005a;
         344: out <= 28'h71e005e;
         345: out <= 28'h7a00060;
         346: out <= 28'h819005f;
         347: out <= 28'h860005d;
         348: out <= 28'h820405d;
         349: out <= 28'h8e2005b;
         350: out <= 28'h9230057;
         351: out <= 28'h8e34057;
         352: out <= 28'h659405f;
         353: out <= 28'h959405c;
         354: out <= 28'h659005c;
         355: out <= 28'h8a2405b;
         356: out <= 28'h9a24058;
         357: out <= 28'h8a20058;
         358: out <= 28'h9da005e;
         359: out <= 28'ha27005c;
         360: out <= 28'h727405c;
         361: out <= 28'h9d60040;
         362: out <= 28'ha670058;
         363: out <= 28'h6274058;
         364: out <= 28'h69a405e;
         365: out <= 28'h9da005d;
         366: out <= 28'h69a405d;
         367: out <= 28'h5964040;
         368: out <= 28'h7560057;
         369: out <= 28'h5964057;
         370: out <= 28'h5e10068;
         371: out <= 28'haa40069;
         372: out <= 28'hae50067;
         373: out <= 28'hb26005d;
         374: out <= 28'hb60005c;
         375: out <= 28'hba30058;
         376: out <= 28'hbd9005a;
         377: out <= 28'hc220056;
         378: out <= 28'hc5f005e;
         379: out <= 28'hc9b0040;
         380: out <= 28'h861ea24;
         381: out <= 28'h5d7ea2a;
         382: out <= 28'h928ea29;
         383: out <= 28'h965ea26;
         384: out <= 28'h9abea2c;
         385: out <= 28'h767ea1d;
         386: out <= 28'h820ea23;
         387: out <= 28'h8edea2e;
         388: out <= 28'h61cea18;
         389: out <= 28'h659ea22;
         390: out <= 28'h72fea30;
         391: out <= 28'h59aea16;
         392: out <= 28'h69fea1b;
         393: out <= 28'h6f1ea32;
         394: out <= 28'h1eea00;
         395: out <= 28'h7a10066;
         396: out <= 28'h79e005a;
         397: out <= 28'h7e4005c;
         398: out <= 28'h7df0040;
         399: out <= 28'h6a0005a;
         400: out <= 28'h180040;
         401: out <= 28'h40;
         402: out <= 28'h623005b;
         403: out <= 28'h8000064;
         404: out <= 28'h89a4061;
         405: out <= 28'h4064;
         406: out <= 28'h5d;
         407: out <= 28'h56;
         408: out <= 28'h69a0061;
         409: out <= 28'h69a4065;
         410: out <= 28'h69a4059;
         411: out <= 28'h25f405e;
         412: out <= 28'h2494065;
         413: out <= 28'h2490056;
         414: out <= 28'h29e005f;
         415: out <= 28'h28a4057;
         416: out <= 28'h28a005d;
         417: out <= 28'h28a0059;
         418: out <= 28'h28a405b;
         419: out <= 28'h2e00062;
         420: out <= 28'h3204062;
         421: out <= 28'h30c0058;
         422: out <= 28'h30c4057;
         423: out <= 28'h340005a;
         424: out <= 28'h380405a;
         425: out <= 28'h38e0058;
         426: out <= 28'h38e0057;
         427: out <= 28'h38e4066;
         428: out <= 28'h38e405c;
         default: out <= 0;
      endcase
endmodule
