library verilog;
use verilog.vl_types.all;
entity ac97_prc is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        valid           : in     vl_logic;
        in_valid        : in     vl_logic_vector(2 downto 0);
        out_slt0        : out    vl_logic_vector(15 downto 0);
        in_slt0         : in     vl_logic_vector(15 downto 0);
        in_slt1         : in     vl_logic_vector(19 downto 0);
        crac_valid      : in     vl_logic;
        crac_wr         : in     vl_logic;
        oc0_cfg         : in     vl_logic_vector(7 downto 0);
        oc1_cfg         : in     vl_logic_vector(7 downto 0);
        oc2_cfg         : in     vl_logic_vector(7 downto 0);
        oc3_cfg         : in     vl_logic_vector(7 downto 0);
        oc4_cfg         : in     vl_logic_vector(7 downto 0);
        oc5_cfg         : in     vl_logic_vector(7 downto 0);
        ic0_cfg         : in     vl_logic_vector(7 downto 0);
        ic1_cfg         : in     vl_logic_vector(7 downto 0);
        ic2_cfg         : in     vl_logic_vector(7 downto 0);
        o3_empty        : in     vl_logic;
        o4_empty        : in     vl_logic;
        o6_empty        : in     vl_logic;
        o7_empty        : in     vl_logic;
        o8_empty        : in     vl_logic;
        o9_empty        : in     vl_logic;
        i3_full         : in     vl_logic;
        i4_full         : in     vl_logic;
        i6_full         : in     vl_logic;
        o3_re           : out    vl_logic;
        o4_re           : out    vl_logic;
        o6_re           : out    vl_logic;
        o7_re           : out    vl_logic;
        o8_re           : out    vl_logic;
        o9_re           : out    vl_logic;
        i3_we           : out    vl_logic;
        i4_we           : out    vl_logic;
        i6_we           : out    vl_logic
    );
end ac97_prc;
