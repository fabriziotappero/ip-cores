module notech_and4 (A,B,C,D,Z);
input A,B,C,D;
output Z;
assign Z=A&B&C&D;
endmodule
