--------------------------------------------------------------------------------
--
-- Title       : ramb_teylor_init_pkg
-- Design      : fp24fftk
-- Author      : Kapitanov
-- Company     :
--
-- Description : FP TWIDDLE GENERATOR
--
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
--		(c) Copyright 2015 													 
--		Kapitanov.                                          				 
--		All rights reserved.                                                 
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use work.fp24_type_pkg.all;

package ramb_teylor_init_pkg is

constant mem_init0:	bit_array_1024x48:=(
(0)=>    "000000000000000000000000000000011001001000011110",
(1)=>    "111111111111111011000011000000011001001000011110",
(2)=>    "111111111111110110000111000000011001001000011100",
(3)=>    "111111111111110001001100000000011001001000011011",
(4)=>    "111111111111101100010000000000011001001000011000",
(5)=>    "111111111111100111010100000000011001001000010011",
(6)=>    "111111111111100010011001000000011001001000001101",
(7)=>    "111111111111011101011101000000011001001000000110",
(8)=>    "111111111111011000100001000000011001001000000000",
(9)=>    "111111111111010011100101000000011001000111111000",
(10)=>    "111111111111001110101010000000011001000111101111",
(11)=>    "111111111111001001101110000000011001000111100100",
(12)=>    "111111111111000100110010000000011001000111011001",
(13)=>    "111111111110111111110110000000011001000111001100",
(14)=>    "111111111110111010111011000000011001000111000000",
(15)=>    "111111111110110110000001000000011001000110110010",
(16)=>    "111111111110110001000101000000011001000110100011",
(17)=>    "111111111110101100001001000000011001000110010010",
(18)=>    "111111111110100111001101000000011001000110000010",
(19)=>    "111111111110100010010010000000011001000101110000",
(20)=>    "111111111110011101010111000000011001000101011101",
(21)=>    "111111111110011000011100000000011001000101001010",
(22)=>    "111111111110010011100000000000011001000100110100",
(23)=>    "111111111110001110100110000000011001000100011110",
(24)=>    "111111111110001001101010000000011001000100001000",
(25)=>    "111111111110000100110000000000011001000011110000",
(26)=>    "111111111101111111110100000000011001000011010111",
(27)=>    "111111111101111010111010000000011001000010111110",
(28)=>    "111111111101110110000000000000011001000010100011",
(29)=>    "111111111101110001000100000000011001000010000111",
(30)=>    "111111111101101100001010000000011001000001101011",
(31)=>    "111111111101100111010000000000011001000001001101",
(32)=>    "111111111101100010010110000000011001000000101111",
(33)=>    "111111111101011101011100000000011001000000010000",
(34)=>    "111111111101011000100001000000011000111111101111",
(35)=>    "111111111101010011100111000000011000111111001110",
(36)=>    "111111111101001110101101000000011000111110101011",
(37)=>    "111111111101001001110011000000011000111110001001",
(38)=>    "111111111101000100111001000000011000111101100100",
(39)=>    "111111111101000000000000000000011000111100111111",
(40)=>    "111111111100111011000110000000011000111100011001",
(41)=>    "111111111100110110001101000000011000111011110010",
(42)=>    "111111111100110001010011000000011000111011001001",
(43)=>    "111111111100101100011011000000011000111010100000",
(44)=>    "111111111100100111100010000000011000111001110110",
(45)=>    "111111111100100010101000000000011000111001001011",
(46)=>    "111111111100011101101111000000011000111000011111",
(47)=>    "111111111100011000110111000000011000110111110010",
(48)=>    "111111111100010011111110000000011000110111000100",
(49)=>    "111111111100001111000111000000011000110110010101",
(50)=>    "111111111100001010001111000000011000110101100110",
(51)=>    "111111111100000101010110000000011000110100110101",
(52)=>    "111111111100000000011111000000011000110100000011",
(53)=>    "111111111011111011100110000000011000110011010001",
(54)=>    "111111111011110110101111000000011000110010011101",
(55)=>    "111111111011110001110111000000011000110001101001",
(56)=>    "111111111011101101000000000000011000110000110100",
(57)=>    "111111111011101000001001000000011000101111111101",
(58)=>    "111111111011100011010010000000011000101111000110",
(59)=>    "111111111011011110011100000000011000101110001101",
(60)=>    "111111111011011001100101000000011000101101010011",
(61)=>    "111111111011010100101110000000011000101100011001",
(62)=>    "111111111011001111111001000000011000101011011101",
(63)=>    "111111111011001011000010000000011000101010100010",
(64)=>    "111111111011000110001100000000011000101001100100",
(65)=>    "111111111011000001010111000000011000101000100111",
(66)=>    "111111111010111100100001000000011000100111101000",
(67)=>    "111111111010110111101100000000011000100110101000",
(68)=>    "111111111010110010110110000000011000100101100111",
(69)=>    "111111111010101110000011000000011000100100100101",
(70)=>    "111111111010101001001101000000011000100011100010",
(71)=>    "111111111010100100011001000000011000100010011110",
(72)=>    "111111111010011111100100000000011000100001011001",
(73)=>    "111111111010011010110000000000011000100000010100",
(74)=>    "111111111010010101111100000000011000011111001101",
(75)=>    "111111111010010001001010000000011000011110000101",
(76)=>    "111111111010001100010110000000011000011100111101",
(77)=>    "111111111010000111100010000000011000011011110011",
(78)=>    "111111111010000010110000000000011000011010101001",
(79)=>    "111111111001111101111101000000011000011001011110",
(80)=>    "111111111001111001001011000000011000011000010001",
(81)=>    "111111111001110100011001000000011000010111000100",
(82)=>    "111111111001101111100110000000011000010101110111",
(83)=>    "111111111001101010110100000000011000010100100111",
(84)=>    "111111111001100110000011000000011000010011010111",
(85)=>    "111111111001100001010001000000011000010010000111",
(86)=>    "111111111001011100100000000000011000010000110101",
(87)=>    "111111111001010111110000000000011000001111100010",
(88)=>    "111111111001010010111111000000011000001110001110",
(89)=>    "111111111001001110010000000000011000001100111010",
(90)=>    "111111111001001001011111000000011000001011100011",
(91)=>    "111111111001000100110000000000011000001010001101",
(92)=>    "111111111000111111111111000000011000001000110101",
(93)=>    "111111111000111011010000000000011000000111011101",
(94)=>    "111111111000110110100010000000011000000110000011",
(95)=>    "111111111000110001110011000000011000000100101010",
(96)=>    "111111111000101101000100000000011000000011001111",
(97)=>    "111111111000101000010110000000011000000001110010",
(98)=>    "111111111000100011101001000000011000000000010101",
(99)=>    "111111111000011110111011000000010111111110110111",
(100)=>    "111111111000011010001110000000010111111101010111",
(101)=>    "111111111000010101100010000000010111111011110111",
(102)=>    "111111111000010000110100000000010111111010011000",
(103)=>    "111111111000001100001000000000010111111000110110",
(104)=>    "111111111000000111011100000000010111110111010011",
(105)=>    "111111111000000010110000000000010111110101101111",
(106)=>    "111111110111111110000110000000010111110100001010",
(107)=>    "111111110111111001011001000000010111110010100110",
(108)=>    "111111110111110100101111000000010111110001000000",
(109)=>    "111111110111110000000101000000010111101111011000",
(110)=>    "111111110111101011011010000000010111101101110000",
(111)=>    "111111110111100110110000000000010111101100000111",
(112)=>    "111111110111100010000111000000010111101010011110",
(113)=>    "111111110111011101011110000000010111101000110011",
(114)=>    "111111110111011000110101000000010111100111000111",
(115)=>    "111111110111010100001100000000010111100101011010",
(116)=>    "111111110111001111100101000000010111100011101100",
(117)=>    "111111110111001010111100000000010111100001111110",
(118)=>    "111111110111000110010101000000010111100000001111",
(119)=>    "111111110111000001101101000000010111011110011110",
(120)=>    "111111110110111101000110000000010111011100101101",
(121)=>    "111111110110111000100000000000010111011010111010",
(122)=>    "111111110110110011111011000000010111011001000111",
(123)=>    "111111110110101111010101000000010111010111010011",
(124)=>    "111111110110101010101111000000010111010101011111",
(125)=>    "111111110110100110001001000000010111010011101001",
(126)=>    "111111110110100001100101000000010111010001110011",
(127)=>    "111111110110011101000001000000010111001111111100",
(128)=>    "111111110110011000011101000000010111001110000011",
(129)=>    "111111110110010011111001000000010111001100001010",
(130)=>    "111111110110001111010110000000010111001010001111",
(131)=>    "111111110110001010110011000000010111001000010011",
(132)=>    "111111110110000110010001000000010111000110011001",
(133)=>    "111111110110000001101110000000010111000100011011",
(134)=>    "111111110101111101001101000000010111000010011101",
(135)=>    "111111110101111000101100000000010111000000011110",
(136)=>    "111111110101110100001011000000010110111110011111",
(137)=>    "111111110101101111101010000000010110111100011110",
(138)=>    "111111110101101011001001000000010110111010011101",
(139)=>    "111111110101100110101010000000010110111000011011",
(140)=>    "111111110101100010001010000000010110110110011001",
(141)=>    "111111110101011101101100000000010110110100010101",
(142)=>    "111111110101011001001101000000010110110010001111",
(143)=>    "111111110101010100101111000000010110110000001010",
(144)=>    "111111110101010000010001000000010110101110000010",
(145)=>    "111111110101001011110101000000010110101011111011",
(146)=>    "111111110101000111010111000000010110101001110011",
(147)=>    "111111110101000010111011000000010110100111101010",
(148)=>    "111111110100111110011110000000010110100101100000",
(149)=>    "111111110100111010000100000000010110100011010110",
(150)=>    "111111110100110101101001000000010110100001001010",
(151)=>    "111111110100110001001110000000010110011110111100",
(152)=>    "111111110100101100110011000000010110011100101111",
(153)=>    "111111110100101000011001000000010110011010100000",
(154)=>    "111111110100100011111111000000010110011000010001",
(155)=>    "111111110100011111100110000000010110010110000001",
(156)=>    "111111110100011011001111000000010110010011110000",
(157)=>    "111111110100010110110101000000010110010001011110",
(158)=>    "111111110100010010011110000000010110001111001100",
(159)=>    "111111110100001110001000000000010110001100111000",
(160)=>    "111111110100001001110000000000010110001010100011",
(161)=>    "111111110100000101011010000000010110001000001110",
(162)=>    "111111110100000001000100000000010110000101110111",
(163)=>    "111111110011111100101110000000010110000011100000",
(164)=>    "111111110011111000011010000000010110000001001001",
(165)=>    "111111110011110100000101000000010101111110110000",
(166)=>    "111111110011101111110001000000010101111100010111",
(167)=>    "111111110011101011011110000000010101111001111100",
(168)=>    "111111110011100111001011000000010101110111100010",
(169)=>    "111111110011100010111000000000010101110101000101",
(170)=>    "111111110011011110100111000000010101110010101000",
(171)=>    "111111110011011010010100000000010101110000001010",
(172)=>    "111111110011010110000100000000010101101101101100",
(173)=>    "111111110011010001110011000000010101101011001100",
(174)=>    "111111110011001101100011000000010101101000101011",
(175)=>    "111111110011001001010011000000010101100110001011",
(176)=>    "111111110011000101000100000000010101100011101001",
(177)=>    "111111110011000000110101000000010101100001000110",
(178)=>    "111111110010111100100111000000010101011110100011",
(179)=>    "111111110010111000011001000000010101011011111110",
(180)=>    "111111110010110100001100000000010101011001011001",
(181)=>    "111111110010110000000000000000010101010110110010",
(182)=>    "111111110010101011110011000000010101010100001100",
(183)=>    "111111110010100111101000000000010101010001100100",
(184)=>    "111111110010100011011101000000010101001110111100",
(185)=>    "111111110010011111010010000000010101001100010010",
(186)=>    "111111110010011011001001000000010101001001101000",
(187)=>    "111111110010010110111111000000010101000110111101",
(188)=>    "111111110010010010110110000000010101000100010000",
(189)=>    "111111110010001110101110000000010101000001100100",
(190)=>    "111111110010001010100110000000010100111110110111",
(191)=>    "111111110010000110011110000000010100111100001000",
(192)=>    "111111110010000010011000000000010100111001011010",
(193)=>    "111111110001111110010001000000010100110110101010",
(194)=>    "111111110001111010001011000000010100110011111001",
(195)=>    "111111110001110110000110000000010100110001000111",
(196)=>    "111111110001110010000001000000010100101110010110",
(197)=>    "111111110001101101111101000000010100101011100011",
(198)=>    "111111110001101001111010000000010100101000101110",
(199)=>    "111111110001100101110110000000010100100101111001",
(200)=>    "111111110001100001110011000000010100100011000101",
(201)=>    "111111110001011101110010000000010100100000001110",
(202)=>    "111111110001011001110000000000010100011101010111",
(203)=>    "111111110001010101110000000000010100011010011111",
(204)=>    "111111110001010001110000000000010100010111100111",
(205)=>    "111111110001001101110000000000010100010100101110",
(206)=>    "111111110001001001110000000000010100010001110011",
(207)=>    "111111110001000101110001000000010100001110111000",
(208)=>    "111111110001000001110100000000010100001011111101",
(209)=>    "111111110000111101110110000000010100001000111111",
(210)=>    "111111110000111001111001000000010100000110000010",
(211)=>    "111111110000110101111110000000010100000011000100",
(212)=>    "111111110000110010000010000000010100000000000101",
(213)=>    "111111110000101110000111000000010011111101000101",
(214)=>    "111111110000101010001100000000010011111010000101",
(215)=>    "111111110000100110010010000000010011110111000100",
(216)=>    "111111110000100010011010000000010011110100000011",
(217)=>    "111111110000011110100000000000010011110001000000",
(218)=>    "111111110000011010101000000000010011101101111100",
(219)=>    "111111110000010110110001000000010011101010110111",
(220)=>    "111111110000010010111011000000010011100111110011",
(221)=>    "111111110000001111000100000000010011100100101101",
(222)=>    "111111110000001011001111000000010011100001100111",
(223)=>    "111111110000000111011010000000010011011110100000",
(224)=>    "111111110000000011100101000000010011011011011000",
(225)=>    "111111101111111111110001000000010011011000001111",
(226)=>    "111111101111111011111110000000010011010101000101",
(227)=>    "111111101111111000001010000000010011010001111100",
(228)=>    "111111101111110100011001000000010011001110110001",
(229)=>    "111111101111110000101000000000010011001011100101",
(230)=>    "111111101111101100110110000000010011001000011000",
(231)=>    "111111101111101001001000000000010011000101001011",
(232)=>    "111111101111100101010111000000010011000001111101",
(233)=>    "111111101111100001101000000000010010111110101110",
(234)=>    "111111101111011101111010000000010010111011011110",
(235)=>    "111111101111011010001101000000010010111000001111",
(236)=>    "111111101111010110011111000000010010110100111110",
(237)=>    "111111101111010010110100000000010010110001101011",
(238)=>    "111111101111001111001000000000010010101110011011",
(239)=>    "111111101111001011011100000000010010101011000111",
(240)=>    "111111101111000111110010000000010010100111110010",
(241)=>    "111111101111000100001000000000010010100100011110",
(242)=>    "111111101111000000100000000000010010100001001010",
(243)=>    "111111101110111100110111000000010010011101110011",
(244)=>    "111111101110111001010001000000010010011010011101",
(245)=>    "111111101110110101101010000000010010010111000110",
(246)=>    "111111101110110010000011000000010010010011101110",
(247)=>    "111111101110101110011101000000010010010000010101",
(248)=>    "111111101110101010111000000000010010001100111100",
(249)=>    "111111101110100111010011000000010010001001100010",
(250)=>    "111111101110100011101111000000010010000110000111",
(251)=>    "111111101110100000001101000000010010000010101011",
(252)=>    "111111101110011100101011000000010001111111001111",
(253)=>    "111111101110011001001000000000010001111011110010",
(254)=>    "111111101110010101101000000000010001111000010101",
(255)=>    "111111101110010010000111000000010001110100110101",
(256)=>    "111111101110001110101000000000010001110001010110",
(257)=>    "111111101110001011001001000000010001101101110111",
(258)=>    "111111101110000111101010000000010001101010010111",
(259)=>    "111111101110000100001100000000010001100110110110",
(260)=>    "111111101110000000101111000000010001100011010100",
(261)=>    "111111101101111101010011000000010001011111110010",
(262)=>    "111111101101111001110111000000010001011100010000",
(263)=>    "111111101101110110011101000000010001011000101100",
(264)=>    "111111101101110011000010000000010001010101000110",
(265)=>    "111111101101101111101010000000010001010001100001",
(266)=>    "111111101101101100010001000000010001001101111100",
(267)=>    "111111101101101000111000000000010001001010010101",
(268)=>    "111111101101100101100001000000010001000110101110",
(269)=>    "111111101101100010001011000000010001000011000111",
(270)=>    "111111101101011110110100000000010000111111011111",
(271)=>    "111111101101011011100000000000010000111011110110",
(272)=>    "111111101101011000001100000000010000111000001100",
(273)=>    "111111101101010100111000000000010000110100100010",
(274)=>    "111111101101010001100100000000010000110000110110",
(275)=>    "111111101101001110010011000000010000101101001011",
(276)=>    "111111101101001011000000000000010000101001011111",
(277)=>    "111111101101000111110000000000010000100101110010",
(278)=>    "111111101101000100100000000000010000100010000101",
(279)=>    "111111101101000001010001000000010000011110010110",
(280)=>    "111111101100111110000010000000010000011010100111",
(281)=>    "111111101100111010110100000000010000010110110111",
(282)=>    "111111101100110111100110000000010000010011001000",
(283)=>    "111111101100110100011010000000010000001111010110",
(284)=>    "111111101100110001001110000000010000001011100110",
(285)=>    "111111101100101110000011000000010000000111110100",
(286)=>    "111111101100101010111010000000010000000100000000",
(287)=>    "111111101100100111101111000000010000000000001101",
(288)=>    "111111101100100100100110000000001111111100011010",
(289)=>    "111111101100100001011111000000001111111000100100",
(290)=>    "111111101100011110010111000000001111110100101111",
(291)=>    "111111101100011011010001000000001111110000111010",
(292)=>    "111111101100011000001011000000001111101101000100",
(293)=>    "111111101100010101000111000000001111101001001101",
(294)=>    "111111101100010010000011000000001111100101010111",
(295)=>    "111111101100001110111110000000001111100001011110",
(296)=>    "111111101100001011111100000000001111011101100101",
(297)=>    "111111101100001000111010000000001111011001101100",
(298)=>    "111111101100000101111001000000001111010101110011",
(299)=>    "111111101100000010111001000000001111010001110111",
(300)=>    "111111101011111111111010000000001111001101111100",
(301)=>    "111111101011111100111010000000001111001010000001",
(302)=>    "111111101011111001111100000000001111000110000101",
(303)=>    "111111101011110111000000000000001111000010001000",
(304)=>    "111111101011110100000010000000001110111110001010",
(305)=>    "111111101011110001000111000000001110111010001101",
(306)=>    "111111101011101110001100000000001110110110001111",
(307)=>    "111111101011101011010001000000001110110010001111",
(308)=>    "111111101011101000010111000000001110101110001111",
(309)=>    "111111101011100101100000000000001110101010001111",
(310)=>    "111111101011100010101000000000001110100110001110",
(311)=>    "111111101011011111110000000000001110100010001101",
(312)=>    "111111101011011100111010000000001110011110001011",
(313)=>    "111111101011011010000101000000001110011010001000",
(314)=>    "111111101011010111010001000000001110010110000101",
(315)=>    "111111101011010100011100000000001110010010000010",
(316)=>    "111111101011010001101001000000001110001101111101",
(317)=>    "111111101011001110110111000000001110001001111000",
(318)=>    "111111101011001100000110000000001110000101110011",
(319)=>    "111111101011001001010100000000001110000001101101",
(320)=>    "111111101011000110100100000000001101111101100111",
(321)=>    "111111101011000011110110000000001101111001100000",
(322)=>    "111111101011000001001000000000001101110101011001",
(323)=>    "111111101010111110011011000000001101110001010001",
(324)=>    "111111101010111011101110000000001101101101001001",
(325)=>    "111111101010111001000001000000001101101000111111",
(326)=>    "111111101010110110010110000000001101100100110110",
(327)=>    "111111101010110011101100000000001101100000101100",
(328)=>    "111111101010110001000011000000001101011100100001",
(329)=>    "111111101010101110011011000000001101011000010110",
(330)=>    "111111101010101011110011000000001101010100001011",
(331)=>    "111111101010101001001100000000001101001111111111",
(332)=>    "111111101010100110100110000000001101001011110010",
(333)=>    "111111101010100100000001000000001101000111100101",
(334)=>    "111111101010100001011100000000001101000011010111",
(335)=>    "111111101010011110111000000000001100111111001001",
(336)=>    "111111101010011100010101000000001100111010111011",
(337)=>    "111111101010011001110011000000001100110110101011",
(338)=>    "111111101010010111010011000000001100110010011011",
(339)=>    "111111101010010100110011000000001100101110001100",
(340)=>    "111111101010010010010011000000001100101001111010",
(341)=>    "111111101010001111110100000000001100100101101011",
(342)=>    "111111101010001101010111000000001100100001011000",
(343)=>    "111111101010001010111010000000001100011101000110",
(344)=>    "111111101010001000011101000000001100011000110100",
(345)=>    "111111101010000110000011000000001100010100100001",
(346)=>    "111111101010000011100111000000001100010000001110",
(347)=>    "111111101010000001001111000000001100001011111001",
(348)=>    "111111101001111110110101000000001100000111100101",
(349)=>    "111111101001111100011110000000001100000011010000",
(350)=>    "111111101001111010000111000000001011111110111010",
(351)=>    "111111101001110111110001000000001011111010100100",
(352)=>    "111111101001110101011011000000001011110110001110",
(353)=>    "111111101001110011000110000000001011110001110111",
(354)=>    "111111101001110000110010000000001011101101100001",
(355)=>    "111111101001101110100000000000001011101001001001",
(356)=>    "111111101001101100001110000000001011100100110000",
(357)=>    "111111101001101001111110000000001011100000011000",
(358)=>    "111111101001100111101101000000001011011011111111",
(359)=>    "111111101001100101011110000000001011010111100110",
(360)=>    "111111101001100011001111000000001011010011001011",
(361)=>    "111111101001100001000010000000001011001110110000",
(362)=>    "111111101001011110110101000000001011001010010110",
(363)=>    "111111101001011100101001000000001011000101111011",
(364)=>    "111111101001011010011111000000001011000001100000",
(365)=>    "111111101001011000010100000000001010111101000100",
(366)=>    "111111101001010110001100000000001010111000101000",
(367)=>    "111111101001010100000011000000001010110100001010",
(368)=>    "111111101001010001111100000000001010101111101101",
(369)=>    "111111101001001111110101000000001010101011001111",
(370)=>    "111111101001001101101111000000001010100110110010",
(371)=>    "111111101001001011101010000000001010100010010010",
(372)=>    "111111101001001001100110000000001010011101110100",
(373)=>    "111111101001000111100100000000001010011001010101",
(374)=>    "111111101001000101100001000000001010010100110101",
(375)=>    "111111101001000011100000000000001010010000010100",
(376)=>    "111111101001000001100000000000001010001011110011",
(377)=>    "111111101000111111100000000000001010000111010010",
(378)=>    "111111101000111101100001000000001010000010110001",
(379)=>    "111111101000111011100011000000001001111110010000",
(380)=>    "111111101000111001100110000000001001111001101110",
(381)=>    "111111101000110111101011000000001001110101001011",
(382)=>    "111111101000110101101111000000001001110000101000",
(383)=>    "111111101000110011110101000000001001101100000110",
(384)=>    "111111101000110001111100000000001001100111100010",
(385)=>    "111111101000110000000011000000001001100010111101",
(386)=>    "111111101000101110001011000000001001011110011001",
(387)=>    "111111101000101100010110000000001001011001110101",
(388)=>    "111111101000101010100000000000001001010101001111",
(389)=>    "111111101000101000101011000000001001010000101010",
(390)=>    "111111101000100110110111000000001001001100000100",
(391)=>    "111111101000100101000101000000001001000111011110",
(392)=>    "111111101000100011010010000000001001000010111000",
(393)=>    "111111101000100001100001000000001000111110010001",
(394)=>    "111111101000011111110000000000001000111001101010",
(395)=>    "111111101000011110000000000000001000110101000010",
(396)=>    "111111101000011100010010000000001000110000011010",
(397)=>    "111111101000011010100100000000001000101011110010",
(398)=>    "111111101000011000111000000000001000100111001001",
(399)=>    "111111101000010111001011000000001000100010100001",
(400)=>    "111111101000010101100001000000001000011101111000",
(401)=>    "111111101000010011110111000000001000011001001111",
(402)=>    "111111101000010010001110000000001000010100100100",
(403)=>    "111111101000010000100111000000001000001111111010",
(404)=>    "111111101000001110111111000000001000001011001111",
(405)=>    "111111101000001101011001000000001000000110100101",
(406)=>    "111111101000001011110100000000001000000001111001",
(407)=>    "111111101000001010010000000000000111111101001110",
(408)=>    "111111101000001000101011000000000111111000100010",
(409)=>    "111111101000000111001000000000000111110011110110",
(410)=>    "111111101000000101100111000000000111101111001010",
(411)=>    "111111101000000100000111000000000111101010011101",
(412)=>    "111111101000000010100111000000000111100101110001",
(413)=>    "111111101000000001000111000000000111100001000011",
(414)=>    "111111100111111111101001000000000111011100010110",
(415)=>    "111111100111111110001100000000000111010111101000",
(416)=>    "111111100111111100110000000000000111010010111010",
(417)=>    "111111100111111011010101000000000111001110001011",
(418)=>    "111111100111111001111011000000000111001001011100",
(419)=>    "111111100111111000100010000000000111000100101110",
(420)=>    "111111100111110111001010000000000110111111111111",
(421)=>    "111111100111110101110010000000000110111011001111",
(422)=>    "111111100111110100011011000000000110110110011111",
(423)=>    "111111100111110011000101000000000110110001101111",
(424)=>    "111111100111110001110000000000000110101101000000",
(425)=>    "111111100111110000011101000000000110101000001111",
(426)=>    "111111100111101111001010000000000110100011011110",
(427)=>    "111111100111101101111000000000000110011110101101",
(428)=>    "111111100111101100101000000000000110011001111011",
(429)=>    "111111100111101011011000000000000110010101001010",
(430)=>    "111111100111101010000111000000000110010000011000",
(431)=>    "111111100111101000111011000000000110001011100110",
(432)=>    "111111100111100111101110000000000110000110110011",
(433)=>    "111111100111100110100001000000000110000010000001",
(434)=>    "111111100111100101010101000000000101111101001111",
(435)=>    "111111100111100100001011000000000101111000011100",
(436)=>    "111111100111100011000010000000000101110011101001",
(437)=>    "111111100111100001111001000000000101101110110101",
(438)=>    "111111100111100000110001000000000101101010000010",
(439)=>    "111111100111011111101010000000000101100101001111",
(440)=>    "111111100111011110100101000000000101100000011011",
(441)=>    "111111100111011101100000000000000101011011100101",
(442)=>    "111111100111011100011101000000000101010110110001",
(443)=>    "111111100111011011011001000000000101010001111100",
(444)=>    "111111100111011010010111000000000101001101001000",
(445)=>    "111111100111011001010111000000000101001000010011",
(446)=>    "111111100111011000010110000000000101000011011101",
(447)=>    "111111100111010111010111000000000100111110101000",
(448)=>    "111111100111010110011010000000000100111001110010",
(449)=>    "111111100111010101011101000000000100110100111101",
(450)=>    "111111100111010100100001000000000100110000000110",
(451)=>    "111111100111010011100101000000000100101011010000",
(452)=>    "111111100111010010101011000000000100100110011001",
(453)=>    "111111100111010001110001000000000100100001100010",
(454)=>    "111111100111010000111001000000000100011100101101",
(455)=>    "111111100111010000000010000000000100010111110110",
(456)=>    "111111100111001111001011000000000100010010111111",
(457)=>    "111111100111001110010101000000000100001110001000",
(458)=>    "111111100111001101100010000000000100001001001111",
(459)=>    "111111100111001100101110000000000100000100011000",
(460)=>    "111111100111001011111011000000000011111111100000",
(461)=>    "111111100111001011001001000000000011111010101001",
(462)=>    "111111100111001010011000000000000011110101110000",
(463)=>    "111111100111001001101001000000000011110000110111",
(464)=>    "111111100111001000111010000000000011101100000000",
(465)=>    "111111100111001000001101000000000011100111001000",
(466)=>    "111111100111000111011111000000000011100010001111",
(467)=>    "111111100111000110110011000000000011011101010111",
(468)=>    "111111100111000110001001000000000011011000011100",
(469)=>    "111111100111000101011110000000000011010011100100",
(470)=>    "111111100111000100110101000000000011001110101011",
(471)=>    "111111100111000100001101000000000011001001110001",
(472)=>    "111111100111000011100101000000000011000100111000",
(473)=>    "111111100111000011000000000000000010111111111110",
(474)=>    "111111100111000010011010000000000010111011000110",
(475)=>    "111111100111000001110110000000000010110110001100",
(476)=>    "111111100111000001010011000000000010110001010001",
(477)=>    "111111100111000000110001000000000010101100010111",
(478)=>    "111111100111000000010000000000000010100111011101",
(479)=>    "111111100110111111101111000000000010100010100011",
(480)=>    "111111100110111111001111000000000010011101101001",
(481)=>    "111111100110111110110001000000000010011000101111",
(482)=>    "111111100110111110010100000000000010010011110100",
(483)=>    "111111100110111101110111000000000010001110111010",
(484)=>    "111111100110111101011011000000000010001001111111",
(485)=>    "111111100110111101000000000000000010000101000100",
(486)=>    "111111100110111100100111000000000010000000001010",
(487)=>    "111111100110111100001110000000000001111011001110",
(488)=>    "111111100110111011110111000000000001110110010100",
(489)=>    "111111100110111011100001000000000001110001011001",
(490)=>    "111111100110111011001011000000000001101100011110",
(491)=>    "111111100110111010110101000000000001100111100011",
(492)=>    "111111100110111010100010000000000001100010100111",
(493)=>    "111111100110111010001111000000000001011101101101",
(494)=>    "111111100110111001111100000000000001011000110001",
(495)=>    "111111100110111001101100000000000001010011110101",
(496)=>    "111111100110111001011011000000000001001110111010",
(497)=>    "111111100110111001001101000000000001001001111110",
(498)=>    "111111100110111000111111000000000001000101000100",
(499)=>    "111111100110111000110010000000000001000000001000",
(500)=>    "111111100110111000100110000000000000111011001100",
(501)=>    "111111100110111000011011000000000000110110010001",
(502)=>    "111111100110111000010000000000000000110001010101",
(503)=>    "111111100110111000000110000000000000101100011001",
(504)=>    "111111100110110111111110000000000000100111011101",
(505)=>    "111111100110110111111000000000000000100010100010",
(506)=>    "111111100110110111110010000000000000011101100110",
(507)=>    "111111100110110111101011000000000000011000101010",
(508)=>    "111111100110110111100111000000000000010011101110",
(509)=>    "111111100110110111100100000000000000001110110011",
(510)=>    "111111100110110111100010000000000000001001110111",
(511)=>    "111111100110110111100010000000000000000100111011",
(512)=>    "111111100110110111100010000000000000000000000000",
(513)=>    "111111100110110111100010111111111111111011000011",
(514)=>    "111111100110110111100010111111111111110110000111",
(515)=>    "111111100110110111100100111111111111110001001100",
(516)=>    "111111100110110111100111111111111111101100010000",
(517)=>    "111111100110110111101011111111111111100111010100",
(518)=>    "111111100110110111110010111111111111100010011001",
(519)=>    "111111100110110111111000111111111111011101011101",
(520)=>    "111111100110110111111110111111111111011000100001",
(521)=>    "111111100110111000000110111111111111010011100101",
(522)=>    "111111100110111000010000111111111111001110101010",
(523)=>    "111111100110111000011011111111111111001001101110",
(524)=>    "111111100110111000100110111111111111000100110010",
(525)=>    "111111100110111000110010111111111110111111110110",
(526)=>    "111111100110111000111111111111111110111010111011",
(527)=>    "111111100110111001001101111111111110110110000001",
(528)=>    "111111100110111001011011111111111110110001000101",
(529)=>    "111111100110111001101100111111111110101100001001",
(530)=>    "111111100110111001111100111111111110100111001101",
(531)=>    "111111100110111010001111111111111110100010010010",
(532)=>    "111111100110111010100010111111111110011101010111",
(533)=>    "111111100110111010110101111111111110011000011100",
(534)=>    "111111100110111011001011111111111110010011100000",
(535)=>    "111111100110111011100001111111111110001110100110",
(536)=>    "111111100110111011110111111111111110001001101010",
(537)=>    "111111100110111100001110111111111110000100110000",
(538)=>    "111111100110111100100111111111111101111111110100",
(539)=>    "111111100110111101000000111111111101111010111010",
(540)=>    "111111100110111101011011111111111101110110000000",
(541)=>    "111111100110111101110111111111111101110001000100",
(542)=>    "111111100110111110010100111111111101101100001010",
(543)=>    "111111100110111110110001111111111101100111010000",
(544)=>    "111111100110111111001111111111111101100010010110",
(545)=>    "111111100110111111101111111111111101011101011100",
(546)=>    "111111100111000000010000111111111101011000100001",
(547)=>    "111111100111000000110001111111111101010011100111",
(548)=>    "111111100111000001010011111111111101001110101101",
(549)=>    "111111100111000001110110111111111101001001110011",
(550)=>    "111111100111000010011010111111111101000100111001",
(551)=>    "111111100111000011000000111111111101000000000000",
(552)=>    "111111100111000011100101111111111100111011000110",
(553)=>    "111111100111000100001101111111111100110110001101",
(554)=>    "111111100111000100110101111111111100110001010011",
(555)=>    "111111100111000101011110111111111100101100011011",
(556)=>    "111111100111000110001001111111111100100111100010",
(557)=>    "111111100111000110110011111111111100100010101000",
(558)=>    "111111100111000111011111111111111100011101101111",
(559)=>    "111111100111001000001101111111111100011000110111",
(560)=>    "111111100111001000111010111111111100010011111110",
(561)=>    "111111100111001001101001111111111100001111000111",
(562)=>    "111111100111001010011000111111111100001010001111",
(563)=>    "111111100111001011001001111111111100000101010110",
(564)=>    "111111100111001011111011111111111100000000011111",
(565)=>    "111111100111001100101110111111111011111011100110",
(566)=>    "111111100111001101100010111111111011110110101111",
(567)=>    "111111100111001110010101111111111011110001110111",
(568)=>    "111111100111001111001011111111111011101101000000",
(569)=>    "111111100111010000000010111111111011101000001001",
(570)=>    "111111100111010000111001111111111011100011010010",
(571)=>    "111111100111010001110001111111111011011110011100",
(572)=>    "111111100111010010101011111111111011011001100101",
(573)=>    "111111100111010011100101111111111011010100101110",
(574)=>    "111111100111010100100001111111111011001111111001",
(575)=>    "111111100111010101011101111111111011001011000010",
(576)=>    "111111100111010110011010111111111011000110001100",
(577)=>    "111111100111010111010111111111111011000001010111",
(578)=>    "111111100111011000010110111111111010111100100001",
(579)=>    "111111100111011001010111111111111010110111101100",
(580)=>    "111111100111011010010111111111111010110010110110",
(581)=>    "111111100111011011011001111111111010101110000011",
(582)=>    "111111100111011100011101111111111010101001001101",
(583)=>    "111111100111011101100000111111111010100100011001",
(584)=>    "111111100111011110100101111111111010011111100100",
(585)=>    "111111100111011111101010111111111010011010110000",
(586)=>    "111111100111100000110001111111111010010101111100",
(587)=>    "111111100111100001111001111111111010010001001010",
(588)=>    "111111100111100011000010111111111010001100010110",
(589)=>    "111111100111100100001011111111111010000111100010",
(590)=>    "111111100111100101010101111111111010000010110000",
(591)=>    "111111100111100110100001111111111001111101111101",
(592)=>    "111111100111100111101110111111111001111001001011",
(593)=>    "111111100111101000111011111111111001110100011001",
(594)=>    "111111100111101010000111111111111001101111100110",
(595)=>    "111111100111101011011000111111111001101010110100",
(596)=>    "111111100111101100101000111111111001100110000011",
(597)=>    "111111100111101101111000111111111001100001010001",
(598)=>    "111111100111101111001010111111111001011100100000",
(599)=>    "111111100111110000011101111111111001010111110000",
(600)=>    "111111100111110001110000111111111001010010111111",
(601)=>    "111111100111110011000101111111111001001110010000",
(602)=>    "111111100111110100011011111111111001001001011111",
(603)=>    "111111100111110101110010111111111001000100110000",
(604)=>    "111111100111110111001010111111111000111111111111",
(605)=>    "111111100111111000100010111111111000111011010000",
(606)=>    "111111100111111001111011111111111000110110100010",
(607)=>    "111111100111111011010101111111111000110001110011",
(608)=>    "111111100111111100110000111111111000101101000100",
(609)=>    "111111100111111110001100111111111000101000010110",
(610)=>    "111111100111111111101001111111111000100011101001",
(611)=>    "111111101000000001000111111111111000011110111011",
(612)=>    "111111101000000010100111111111111000011010001110",
(613)=>    "111111101000000100000111111111111000010101100010",
(614)=>    "111111101000000101100111111111111000010000110100",
(615)=>    "111111101000000111001000111111111000001100001000",
(616)=>    "111111101000001000101011111111111000000111011100",
(617)=>    "111111101000001010010000111111111000000010110000",
(618)=>    "111111101000001011110100111111110111111110000110",
(619)=>    "111111101000001101011001111111110111111001011001",
(620)=>    "111111101000001110111111111111110111110100101111",
(621)=>    "111111101000010000100111111111110111110000000101",
(622)=>    "111111101000010010001110111111110111101011011010",
(623)=>    "111111101000010011110111111111110111100110110000",
(624)=>    "111111101000010101100001111111110111100010000111",
(625)=>    "111111101000010111001011111111110111011101011110",
(626)=>    "111111101000011000111000111111110111011000110101",
(627)=>    "111111101000011010100100111111110111010100001100",
(628)=>    "111111101000011100010010111111110111001111100101",
(629)=>    "111111101000011110000000111111110111001010111100",
(630)=>    "111111101000011111110000111111110111000110010101",
(631)=>    "111111101000100001100001111111110111000001101101",
(632)=>    "111111101000100011010010111111110110111101000110",
(633)=>    "111111101000100101000101111111110110111000100000",
(634)=>    "111111101000100110110111111111110110110011111011",
(635)=>    "111111101000101000101011111111110110101111010101",
(636)=>    "111111101000101010100000111111110110101010101111",
(637)=>    "111111101000101100010110111111110110100110001001",
(638)=>    "111111101000101110001011111111110110100001100101",
(639)=>    "111111101000110000000011111111110110011101000001",
(640)=>    "111111101000110001111100111111110110011000011101",
(641)=>    "111111101000110011110101111111110110010011111001",
(642)=>    "111111101000110101101111111111110110001111010110",
(643)=>    "111111101000110111101011111111110110001010110011",
(644)=>    "111111101000111001100110111111110110000110010001",
(645)=>    "111111101000111011100011111111110110000001101110",
(646)=>    "111111101000111101100001111111110101111101001101",
(647)=>    "111111101000111111100000111111110101111000101100",
(648)=>    "111111101001000001100000111111110101110100001011",
(649)=>    "111111101001000011100000111111110101101111101010",
(650)=>    "111111101001000101100001111111110101101011001001",
(651)=>    "111111101001000111100100111111110101100110101010",
(652)=>    "111111101001001001100110111111110101100010001010",
(653)=>    "111111101001001011101010111111110101011101101100",
(654)=>    "111111101001001101101111111111110101011001001101",
(655)=>    "111111101001001111110101111111110101010100101111",
(656)=>    "111111101001010001111100111111110101010000010001",
(657)=>    "111111101001010100000011111111110101001011110101",
(658)=>    "111111101001010110001100111111110101000111010111",
(659)=>    "111111101001011000010100111111110101000010111011",
(660)=>    "111111101001011010011111111111110100111110011110",
(661)=>    "111111101001011100101001111111110100111010000100",
(662)=>    "111111101001011110110101111111110100110101101001",
(663)=>    "111111101001100001000010111111110100110001001110",
(664)=>    "111111101001100011001111111111110100101100110011",
(665)=>    "111111101001100101011110111111110100101000011001",
(666)=>    "111111101001100111101101111111110100100011111111",
(667)=>    "111111101001101001111110111111110100011111100110",
(668)=>    "111111101001101100001110111111110100011011001111",
(669)=>    "111111101001101110100000111111110100010110110101",
(670)=>    "111111101001110000110010111111110100010010011110",
(671)=>    "111111101001110011000110111111110100001110001000",
(672)=>    "111111101001110101011011111111110100001001110000",
(673)=>    "111111101001110111110001111111110100000101011010",
(674)=>    "111111101001111010000111111111110100000001000100",
(675)=>    "111111101001111100011110111111110011111100101110",
(676)=>    "111111101001111110110101111111110011111000011010",
(677)=>    "111111101010000001001111111111110011110100000101",
(678)=>    "111111101010000011100111111111110011101111110001",
(679)=>    "111111101010000110000011111111110011101011011110",
(680)=>    "111111101010001000011101111111110011100111001011",
(681)=>    "111111101010001010111010111111110011100010111000",
(682)=>    "111111101010001101010111111111110011011110100111",
(683)=>    "111111101010001111110100111111110011011010010100",
(684)=>    "111111101010010010010011111111110011010110000100",
(685)=>    "111111101010010100110011111111110011010001110011",
(686)=>    "111111101010010111010011111111110011001101100011",
(687)=>    "111111101010011001110011111111110011001001010011",
(688)=>    "111111101010011100010101111111110011000101000100",
(689)=>    "111111101010011110111000111111110011000000110101",
(690)=>    "111111101010100001011100111111110010111100100111",
(691)=>    "111111101010100100000001111111110010111000011001",
(692)=>    "111111101010100110100110111111110010110100001100",
(693)=>    "111111101010101001001100111111110010110000000000",
(694)=>    "111111101010101011110011111111110010101011110011",
(695)=>    "111111101010101110011011111111110010100111101000",
(696)=>    "111111101010110001000011111111110010100011011101",
(697)=>    "111111101010110011101100111111110010011111010010",
(698)=>    "111111101010110110010110111111110010011011001001",
(699)=>    "111111101010111001000001111111110010010110111111",
(700)=>    "111111101010111011101110111111110010010010110110",
(701)=>    "111111101010111110011011111111110010001110101110",
(702)=>    "111111101011000001001000111111110010001010100110",
(703)=>    "111111101011000011110110111111110010000110011110",
(704)=>    "111111101011000110100100111111110010000010011000",
(705)=>    "111111101011001001010100111111110001111110010001",
(706)=>    "111111101011001100000110111111110001111010001011",
(707)=>    "111111101011001110110111111111110001110110000110",
(708)=>    "111111101011010001101001111111110001110010000001",
(709)=>    "111111101011010100011100111111110001101101111101",
(710)=>    "111111101011010111010001111111110001101001111010",
(711)=>    "111111101011011010000101111111110001100101110110",
(712)=>    "111111101011011100111010111111110001100001110011",
(713)=>    "111111101011011111110000111111110001011101110010",
(714)=>    "111111101011100010101000111111110001011001110000",
(715)=>    "111111101011100101100000111111110001010101110000",
(716)=>    "111111101011101000010111111111110001010001110000",
(717)=>    "111111101011101011010001111111110001001101110000",
(718)=>    "111111101011101110001100111111110001001001110000",
(719)=>    "111111101011110001000111111111110001000101110001",
(720)=>    "111111101011110100000010111111110001000001110100",
(721)=>    "111111101011110111000000111111110000111101110110",
(722)=>    "111111101011111001111100111111110000111001111001",
(723)=>    "111111101011111100111010111111110000110101111110",
(724)=>    "111111101011111111111010111111110000110010000010",
(725)=>    "111111101100000010111001111111110000101110000111",
(726)=>    "111111101100000101111001111111110000101010001100",
(727)=>    "111111101100001000111010111111110000100110010010",
(728)=>    "111111101100001011111100111111110000100010011010",
(729)=>    "111111101100001110111110111111110000011110100000",
(730)=>    "111111101100010010000011111111110000011010101000",
(731)=>    "111111101100010101000111111111110000010110110001",
(732)=>    "111111101100011000001011111111110000010010111011",
(733)=>    "111111101100011011010001111111110000001111000100",
(734)=>    "111111101100011110010111111111110000001011001111",
(735)=>    "111111101100100001011111111111110000000111011010",
(736)=>    "111111101100100100100110111111110000000011100101",
(737)=>    "111111101100100111101111111111101111111111110001",
(738)=>    "111111101100101010111010111111101111111011111110",
(739)=>    "111111101100101110000011111111101111111000001010",
(740)=>    "111111101100110001001110111111101111110100011001",
(741)=>    "111111101100110100011010111111101111110000101000",
(742)=>    "111111101100110111100110111111101111101100110110",
(743)=>    "111111101100111010110100111111101111101001001000",
(744)=>    "111111101100111110000010111111101111100101010111",
(745)=>    "111111101101000001010001111111101111100001101000",
(746)=>    "111111101101000100100000111111101111011101111010",
(747)=>    "111111101101000111110000111111101111011010001101",
(748)=>    "111111101101001011000000111111101111010110011111",
(749)=>    "111111101101001110010011111111101111010010110100",
(750)=>    "111111101101010001100100111111101111001111001000",
(751)=>    "111111101101010100111000111111101111001011011100",
(752)=>    "111111101101011000001100111111101111000111110010",
(753)=>    "111111101101011011100000111111101111000100001000",
(754)=>    "111111101101011110110100111111101111000000100000",
(755)=>    "111111101101100010001011111111101110111100110111",
(756)=>    "111111101101100101100001111111101110111001010001",
(757)=>    "111111101101101000111000111111101110110101101010",
(758)=>    "111111101101101100010001111111101110110010000011",
(759)=>    "111111101101101111101010111111101110101110011101",
(760)=>    "111111101101110011000010111111101110101010111000",
(761)=>    "111111101101110110011101111111101110100111010011",
(762)=>    "111111101101111001110111111111101110100011101111",
(763)=>    "111111101101111101010011111111101110100000001101",
(764)=>    "111111101110000000101111111111101110011100101011",
(765)=>    "111111101110000100001100111111101110011001001000",
(766)=>    "111111101110000111101010111111101110010101101000",
(767)=>    "111111101110001011001001111111101110010010000111",
(768)=>    "111111101110001110101000111111101110001110101000",
(769)=>    "111111101110010010000111111111101110001011001001",
(770)=>    "111111101110010101101000111111101110000111101010",
(771)=>    "111111101110011001001000111111101110000100001100",
(772)=>    "111111101110011100101011111111101110000000101111",
(773)=>    "111111101110100000001101111111101101111101010011",
(774)=>    "111111101110100011101111111111101101111001110111",
(775)=>    "111111101110100111010011111111101101110110011101",
(776)=>    "111111101110101010111000111111101101110011000010",
(777)=>    "111111101110101110011101111111101101101111101010",
(778)=>    "111111101110110010000011111111101101101100010001",
(779)=>    "111111101110110101101010111111101101101000111000",
(780)=>    "111111101110111001010001111111101101100101100001",
(781)=>    "111111101110111100110111111111101101100010001011",
(782)=>    "111111101111000000100000111111101101011110110100",
(783)=>    "111111101111000100001000111111101101011011100000",
(784)=>    "111111101111000111110010111111101101011000001100",
(785)=>    "111111101111001011011100111111101101010100111000",
(786)=>    "111111101111001111001000111111101101010001100100",
(787)=>    "111111101111010010110100111111101101001110010011",
(788)=>    "111111101111010110011111111111101101001011000000",
(789)=>    "111111101111011010001101111111101101000111110000",
(790)=>    "111111101111011101111010111111101101000100100000",
(791)=>    "111111101111100001101000111111101101000001010001",
(792)=>    "111111101111100101010111111111101100111110000010",
(793)=>    "111111101111101001001000111111101100111010110100",
(794)=>    "111111101111101100110110111111101100110111100110",
(795)=>    "111111101111110000101000111111101100110100011010",
(796)=>    "111111101111110100011001111111101100110001001110",
(797)=>    "111111101111111000001010111111101100101110000011",
(798)=>    "111111101111111011111110111111101100101010111010",
(799)=>    "111111101111111111110001111111101100100111101111",
(800)=>    "111111110000000011100101111111101100100100100110",
(801)=>    "111111110000000111011010111111101100100001011111",
(802)=>    "111111110000001011001111111111101100011110010111",
(803)=>    "111111110000001111000100111111101100011011010001",
(804)=>    "111111110000010010111011111111101100011000001011",
(805)=>    "111111110000010110110001111111101100010101000111",
(806)=>    "111111110000011010101000111111101100010010000011",
(807)=>    "111111110000011110100000111111101100001110111110",
(808)=>    "111111110000100010011010111111101100001011111100",
(809)=>    "111111110000100110010010111111101100001000111010",
(810)=>    "111111110000101010001100111111101100000101111001",
(811)=>    "111111110000101110000111111111101100000010111001",
(812)=>    "111111110000110010000010111111101011111111111010",
(813)=>    "111111110000110101111110111111101011111100111010",
(814)=>    "111111110000111001111001111111101011111001111100",
(815)=>    "111111110000111101110110111111101011110111000000",
(816)=>    "111111110001000001110100111111101011110100000010",
(817)=>    "111111110001000101110001111111101011110001000111",
(818)=>    "111111110001001001110000111111101011101110001100",
(819)=>    "111111110001001101110000111111101011101011010001",
(820)=>    "111111110001010001110000111111101011101000010111",
(821)=>    "111111110001010101110000111111101011100101100000",
(822)=>    "111111110001011001110000111111101011100010101000",
(823)=>    "111111110001011101110010111111101011011111110000",
(824)=>    "111111110001100001110011111111101011011100111010",
(825)=>    "111111110001100101110110111111101011011010000101",
(826)=>    "111111110001101001111010111111101011010111010001",
(827)=>    "111111110001101101111101111111101011010100011100",
(828)=>    "111111110001110010000001111111101011010001101001",
(829)=>    "111111110001110110000110111111101011001110110111",
(830)=>    "111111110001111010001011111111101011001100000110",
(831)=>    "111111110001111110010001111111101011001001010100",
(832)=>    "111111110010000010011000111111101011000110100100",
(833)=>    "111111110010000110011110111111101011000011110110",
(834)=>    "111111110010001010100110111111101011000001001000",
(835)=>    "111111110010001110101110111111101010111110011011",
(836)=>    "111111110010010010110110111111101010111011101110",
(837)=>    "111111110010010110111111111111101010111001000001",
(838)=>    "111111110010011011001001111111101010110110010110",
(839)=>    "111111110010011111010010111111101010110011101100",
(840)=>    "111111110010100011011101111111101010110001000011",
(841)=>    "111111110010100111101000111111101010101110011011",
(842)=>    "111111110010101011110011111111101010101011110011",
(843)=>    "111111110010110000000000111111101010101001001100",
(844)=>    "111111110010110100001100111111101010100110100110",
(845)=>    "111111110010111000011001111111101010100100000001",
(846)=>    "111111110010111100100111111111101010100001011100",
(847)=>    "111111110011000000110101111111101010011110111000",
(848)=>    "111111110011000101000100111111101010011100010101",
(849)=>    "111111110011001001010011111111101010011001110011",
(850)=>    "111111110011001101100011111111101010010111010011",
(851)=>    "111111110011010001110011111111101010010100110011",
(852)=>    "111111110011010110000100111111101010010010010011",
(853)=>    "111111110011011010010100111111101010001111110100",
(854)=>    "111111110011011110100111111111101010001101010111",
(855)=>    "111111110011100010111000111111101010001010111010",
(856)=>    "111111110011100111001011111111101010001000011101",
(857)=>    "111111110011101011011110111111101010000110000011",
(858)=>    "111111110011101111110001111111101010000011100111",
(859)=>    "111111110011110100000101111111101010000001001111",
(860)=>    "111111110011111000011010111111101001111110110101",
(861)=>    "111111110011111100101110111111101001111100011110",
(862)=>    "111111110100000001000100111111101001111010000111",
(863)=>    "111111110100000101011010111111101001110111110001",
(864)=>    "111111110100001001110000111111101001110101011011",
(865)=>    "111111110100001110001000111111101001110011000110",
(866)=>    "111111110100010010011110111111101001110000110010",
(867)=>    "111111110100010110110101111111101001101110100000",
(868)=>    "111111110100011011001111111111101001101100001110",
(869)=>    "111111110100011111100110111111101001101001111110",
(870)=>    "111111110100100011111111111111101001100111101101",
(871)=>    "111111110100101000011001111111101001100101011110",
(872)=>    "111111110100101100110011111111101001100011001111",
(873)=>    "111111110100110001001110111111101001100001000010",
(874)=>    "111111110100110101101001111111101001011110110101",
(875)=>    "111111110100111010000100111111101001011100101001",
(876)=>    "111111110100111110011110111111101001011010011111",
(877)=>    "111111110101000010111011111111101001011000010100",
(878)=>    "111111110101000111010111111111101001010110001100",
(879)=>    "111111110101001011110101111111101001010100000011",
(880)=>    "111111110101010000010001111111101001010001111100",
(881)=>    "111111110101010100101111111111101001001111110101",
(882)=>    "111111110101011001001101111111101001001101101111",
(883)=>    "111111110101011101101100111111101001001011101010",
(884)=>    "111111110101100010001010111111101001001001100110",
(885)=>    "111111110101100110101010111111101001000111100100",
(886)=>    "111111110101101011001001111111101001000101100001",
(887)=>    "111111110101101111101010111111101001000011100000",
(888)=>    "111111110101110100001011111111101001000001100000",
(889)=>    "111111110101111000101100111111101000111111100000",
(890)=>    "111111110101111101001101111111101000111101100001",
(891)=>    "111111110110000001101110111111101000111011100011",
(892)=>    "111111110110000110010001111111101000111001100110",
(893)=>    "111111110110001010110011111111101000110111101011",
(894)=>    "111111110110001111010110111111101000110101101111",
(895)=>    "111111110110010011111001111111101000110011110101",
(896)=>    "111111110110011000011101111111101000110001111100",
(897)=>    "111111110110011101000001111111101000110000000011",
(898)=>    "111111110110100001100101111111101000101110001011",
(899)=>    "111111110110100110001001111111101000101100010110",
(900)=>    "111111110110101010101111111111101000101010100000",
(901)=>    "111111110110101111010101111111101000101000101011",
(902)=>    "111111110110110011111011111111101000100110110111",
(903)=>    "111111110110111000100000111111101000100101000101",
(904)=>    "111111110110111101000110111111101000100011010010",
(905)=>    "111111110111000001101101111111101000100001100001",
(906)=>    "111111110111000110010101111111101000011111110000",
(907)=>    "111111110111001010111100111111101000011110000000",
(908)=>    "111111110111001111100101111111101000011100010010",
(909)=>    "111111110111010100001100111111101000011010100100",
(910)=>    "111111110111011000110101111111101000011000111000",
(911)=>    "111111110111011101011110111111101000010111001011",
(912)=>    "111111110111100010000111111111101000010101100001",
(913)=>    "111111110111100110110000111111101000010011110111",
(914)=>    "111111110111101011011010111111101000010010001110",
(915)=>    "111111110111110000000101111111101000010000100111",
(916)=>    "111111110111110100101111111111101000001110111111",
(917)=>    "111111110111111001011001111111101000001101011001",
(918)=>    "111111110111111110000110111111101000001011110100",
(919)=>    "111111111000000010110000111111101000001010010000",
(920)=>    "111111111000000111011100111111101000001000101011",
(921)=>    "111111111000001100001000111111101000000111001000",
(922)=>    "111111111000010000110100111111101000000101100111",
(923)=>    "111111111000010101100010111111101000000100000111",
(924)=>    "111111111000011010001110111111101000000010100111",
(925)=>    "111111111000011110111011111111101000000001000111",
(926)=>    "111111111000100011101001111111100111111111101001",
(927)=>    "111111111000101000010110111111100111111110001100",
(928)=>    "111111111000101101000100111111100111111100110000",
(929)=>    "111111111000110001110011111111100111111011010101",
(930)=>    "111111111000110110100010111111100111111001111011",
(931)=>    "111111111000111011010000111111100111111000100010",
(932)=>    "111111111000111111111111111111100111110111001010",
(933)=>    "111111111001000100110000111111100111110101110010",
(934)=>    "111111111001001001011111111111100111110100011011",
(935)=>    "111111111001001110010000111111100111110011000101",
(936)=>    "111111111001010010111111111111100111110001110000",
(937)=>    "111111111001010111110000111111100111110000011101",
(938)=>    "111111111001011100100000111111100111101111001010",
(939)=>    "111111111001100001010001111111100111101101111000",
(940)=>    "111111111001100110000011111111100111101100101000",
(941)=>    "111111111001101010110100111111100111101011011000",
(942)=>    "111111111001101111100110111111100111101010000111",
(943)=>    "111111111001110100011001111111100111101000111011",
(944)=>    "111111111001111001001011111111100111100111101110",
(945)=>    "111111111001111101111101111111100111100110100001",
(946)=>    "111111111010000010110000111111100111100101010101",
(947)=>    "111111111010000111100010111111100111100100001011",
(948)=>    "111111111010001100010110111111100111100011000010",
(949)=>    "111111111010010001001010111111100111100001111001",
(950)=>    "111111111010010101111100111111100111100000110001",
(951)=>    "111111111010011010110000111111100111011111101010",
(952)=>    "111111111010011111100100111111100111011110100101",
(953)=>    "111111111010100100011001111111100111011101100000",
(954)=>    "111111111010101001001101111111100111011100011101",
(955)=>    "111111111010101110000011111111100111011011011001",
(956)=>    "111111111010110010110110111111100111011010010111",
(957)=>    "111111111010110111101100111111100111011001010111",
(958)=>    "111111111010111100100001111111100111011000010110",
(959)=>    "111111111011000001010111111111100111010111010111",
(960)=>    "111111111011000110001100111111100111010110011010",
(961)=>    "111111111011001011000010111111100111010101011101",
(962)=>    "111111111011001111111001111111100111010100100001",
(963)=>    "111111111011010100101110111111100111010011100101",
(964)=>    "111111111011011001100101111111100111010010101011",
(965)=>    "111111111011011110011100111111100111010001110001",
(966)=>    "111111111011100011010010111111100111010000111001",
(967)=>    "111111111011101000001001111111100111010000000010",
(968)=>    "111111111011101101000000111111100111001111001011",
(969)=>    "111111111011110001110111111111100111001110010101",
(970)=>    "111111111011110110101111111111100111001101100010",
(971)=>    "111111111011111011100110111111100111001100101110",
(972)=>    "111111111100000000011111111111100111001011111011",
(973)=>    "111111111100000101010110111111100111001011001001",
(974)=>    "111111111100001010001111111111100111001010011000",
(975)=>    "111111111100001111000111111111100111001001101001",
(976)=>    "111111111100010011111110111111100111001000111010",
(977)=>    "111111111100011000110111111111100111001000001101",
(978)=>    "111111111100011101101111111111100111000111011111",
(979)=>    "111111111100100010101000111111100111000110110011",
(980)=>    "111111111100100111100010111111100111000110001001",
(981)=>    "111111111100101100011011111111100111000101011110",
(982)=>    "111111111100110001010011111111100111000100110101",
(983)=>    "111111111100110110001101111111100111000100001101",
(984)=>    "111111111100111011000110111111100111000011100101",
(985)=>    "111111111101000000000000111111100111000011000000",
(986)=>    "111111111101000100111001111111100111000010011010",
(987)=>    "111111111101001001110011111111100111000001110110",
(988)=>    "111111111101001110101101111111100111000001010011",
(989)=>    "111111111101010011100111111111100111000000110001",
(990)=>    "111111111101011000100001111111100111000000010000",
(991)=>    "111111111101011101011100111111100110111111101111",
(992)=>    "111111111101100010010110111111100110111111001111",
(993)=>    "111111111101100111010000111111100110111110110001",
(994)=>    "111111111101101100001010111111100110111110010100",
(995)=>    "111111111101110001000100111111100110111101110111",
(996)=>    "111111111101110110000000111111100110111101011011",
(997)=>    "111111111101111010111010111111100110111101000000",
(998)=>    "111111111101111111110100111111100110111100100111",
(999)=>    "111111111110000100110000111111100110111100001110",
(1000)=>    "111111111110001001101010111111100110111011110111",
(1001)=>    "111111111110001110100110111111100110111011100001",
(1002)=>    "111111111110010011100000111111100110111011001011",
(1003)=>    "111111111110011000011100111111100110111010110101",
(1004)=>    "111111111110011101010111111111100110111010100010",
(1005)=>    "111111111110100010010010111111100110111010001111",
(1006)=>    "111111111110100111001101111111100110111001111100",
(1007)=>    "111111111110101100001001111111100110111001101100",
(1008)=>    "111111111110110001000101111111100110111001011011",
(1009)=>    "111111111110110110000001111111100110111001001101",
(1010)=>    "111111111110111010111011111111100110111000111111",
(1011)=>    "111111111110111111110110111111100110111000110010",
(1012)=>    "111111111111000100110010111111100110111000100110",
(1013)=>    "111111111111001001101110111111100110111000011011",
(1014)=>    "111111111111001110101010111111100110111000010000",
(1015)=>    "111111111111010011100101111111100110111000000110",
(1016)=>    "111111111111011000100001111111100110110111111110",
(1017)=>    "111111111111011101011101111111100110110111111000",
(1018)=>    "111111111111100010011001111111100110110111110010",
(1019)=>    "111111111111100111010100111111100110110111101011",
(1020)=>    "111111111111101100010000111111100110110111100111",
(1021)=>    "111111111111110001001100111111100110110111100100",
(1022)=>    "111111111111110110000111111111100110110111100010",
(1023)=>    "111111111111111011000011111111100110110111100010"

);
end package;
