-- Copyright 2015, J�rgen Defurne
--
-- This file is part of the Experimental Unstable CPU System.
--
-- The Experimental Unstable CPU System Is free software: you can redistribute
-- it and/or modify it under the terms of the GNU Lesser General Public License
-- as published by the Free Software Foundation, either version 3 of the
-- License, or (at your option) any later version.
--
-- The Experimental Unstable CPU System is distributed in the hope that it will
-- be useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU Lesser
-- General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public License
-- along with Experimental Unstable CPU System. If not, see
-- http://www.gnu.org/licenses/lgpl.txt.


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY memory_controller IS
  
  PORT (
    RST  : IN  STD_LOGIC;
    CLK  : IN  STD_LOGIC;
    SEL  : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    EN0  : OUT STD_LOGIC;
    EN1  : OUT STD_LOGIC;
    FULL : OUT STD_LOGIC;
    PULL : IN  STD_LOGIC);

END ENTITY memory_controller;
