module vc_tb ();

dut: vc (
    .
)