-------------------------------------------------------------------------------
-- $Id: t400_por-c.vhd 179 2009-04-01 19:48:38Z arniml $
-------------------------------------------------------------------------------

configuration t400_por_rtl_c0 of t400_por is

  for spartan
  end for;

end t400_por_rtl_c0;
