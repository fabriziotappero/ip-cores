-------------------------------------------------------------------------------
--
-- $Id: t400_mnemonic_pack-p.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2008, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

use work.t400_pack.byte_t;

package t400_mnemonic_pack is

  -- Mnemonics ----------------------------------------------------------------
  type    mnemonic_t is (-- Arithmetic instructions
                         MN_ASC,
                         MN_ADD,
                         MN_ADT,
                         MN_AISC,
                         MN_CASC,
                         MN_CLRA,
                         MN_COMP,
                         MN_NOP,
                         MN_C,
                         MN_XOR,
                         -- Transfer of control instructions
                         MN_JID,
                         MN_JMP,
                         MN_JP_JSRP,
                         MN_JSR,
                         MN_RET,
                         MN_RETSK,
                         -- Memory reference instructions
                         MN_LD,
                         MN_LDD_XAD,
                         MN_LQID,
                         MN_RMB,
                         MN_SMB,
                         MN_STII,
                         MN_X,
                         MN_XDS,
                         MN_XIS,
                         -- Register reference instructions
                         MN_CAB,
                         MN_CBA,
                         MN_LBI,
                         MN_XABR,
                         -- Test instructions
                         MN_SKC,
                         MN_SKE,
                         MN_SKMBZ,
                         MN_SKT,
                         -- Input/output instructions
                         MN_EXT,
                         MN_XAS);

  type mnemonic_rec_t is
    record
      mnemonic   : mnemonic_t;
      multi_byte : boolean;
    end record;

  function decode_opcode_f(opcode   : in byte_t;
                           opt_type : in integer) return
    mnemonic_rec_t;

end t400_mnemonic_pack;


library ieee;
use ieee.std_logic_1164.all;

use work.t400_opt_pack.t400_opt_type_410_c;

package body t400_mnemonic_pack is

  function decode_opcode_f(opcode   : in byte_t;
                           opt_type : in integer) return
    mnemonic_rec_t is
    variable t41x_type_v  : boolean;
    variable mnemonic_v   : mnemonic_t;
    variable multi_byte_v : boolean;
    variable result_v     : mnemonic_rec_t;
  begin
    -- default assignment
    mnemonic_v   := MN_NOP;
    multi_byte_v := false;
    -- determine type
    t41x_type_v  := opt_type = t400_opt_type_410_c;

    case opcode is
      -- Mnemonic ASC----------------------------------------------------------
      when "00110000" =>
        mnemonic_v   := MN_ASC;

      -- Mnemonic ADD ---------------------------------------------------------
      when "00110001" =>
        mnemonic_v   := MN_ADD;

      -- Mnemonic ADT ---------------------------------------------------------
      when "01001010" =>
        if not t41x_type_v then
          mnemonic_v := MN_ADT;
        end if;

      -- Mnemonic AISC --------------------------------------------------------
      when "01010001" | "01010010" | "01010011" |
           "01010100" | "01010101" | "01010110" | "01010111" |
           "01011000" | "01011001" | "01011010" | "01011011" |
           "01011100" | "01011101" | "01011110" | "01011111" =>
        mnemonic_v   := MN_AISC;

      -- Mnemonic CASC --------------------------------------------------------
      when "00010000" =>
        if not t41x_type_v then
          mnemonic_v := MN_CASC;
        end if;

      -- Mnemonic CLRA --------------------------------------------------------
      when "00000000" =>
        mnemonic_v   := MN_CLRA;

      -- Mnemonic COMP --------------------------------------------------------
      when "01000000" =>
        mnemonic_v   := MN_COMP;

      -- Mnemonic NOP ---------------------------------------------------------
      when "01000100" =>
        mnemonic_v   := MN_NOP;

      -- Mnemonic C -----------------------------------------------------------
      when "00110010" |                                         -- RC
           "00100010" =>                                        -- SC
        mnemonic_v   := MN_C;

      -- Mnemonic XOR ---------------------------------------------------------
      when "00000010" =>
        mnemonic_v   := MN_XOR;

      -- Mnemonic JID ---------------------------------------------------------
      when "11111111" =>
        mnemonic_v   := MN_JID;

      -- Mnemonic JMP ---------------------------------------------------------
      when "01100000" | "01100001" | "01100010" | "01100011" =>
        mnemonic_v   := MN_JMP;
        multi_byte_v := true;

      -- Mnemonic JP_JSRP -----------------------------------------------------
      when "10000000" | "10000001" | "10000010" | "10000011" |
           "10000100" | "10000101" | "10000110" | "10000111" |
           "10001000" | "10001001" | "10001010" | "10001011" |
           "10001100" | "10001101" | "10001110" | "10001111" |
           "10010000" | "10010001" | "10010010" | "10010011" |
           "10010100" | "10010101" | "10010110" | "10010111" |
           "10011000" | "10011001" | "10011010" | "10011011" |
           "10011100" | "10011101" | "10011110" | "10011111" |
           "10100000" | "10100001" | "10100010" | "10100011" |
           "10100100" | "10100101" | "10100110" | "10100111" |
           "10101000" | "10101001" | "10101010" | "10101011" |
           "10101100" | "10101101" | "10101110" | "10101111" |
           "10110000" | "10110001" | "10110010" | "10110011" |
           "10110100" | "10110101" | "10110110" | "10110111" |
           "10111000" | "10111001" | "10111010" | "10111011" |
           "10111100" | "10111101" | "10111110" |
           "11000000" | "11000001" | "11000010" | "11000011" |
           "11000100" | "11000101" | "11000110" | "11000111" |
           "11001000" | "11001001" | "11001010" | "11001011" |
           "11001100" | "11001101" | "11001110" | "11001111" |
           "11010000" | "11010001" | "11010010" | "11010011" |
           "11010100" | "11010101" | "11010110" | "11010111" |
           "11011000" | "11011001" | "11011010" | "11011011" |
           "11011100" | "11011101" | "11011110" | "11011111" |
           "11100000" | "11100001" | "11100010" | "11100011" |
           "11100100" | "11100101" | "11100110" | "11100111" |
           "11101000" | "11101001" | "11101010" | "11101011" |
           "11101100" | "11101101" | "11101110" | "11101111" |
           "11110000" | "11110001" | "11110010" | "11110011" |
           "11110100" | "11110101" | "11110110" | "11110111" |
           "11111000" | "11111001" | "11111010" | "11111011" |
           "11111100" | "11111101" | "11111110" =>
        mnemonic_v   := MN_JP_JSRP;

      -- Mnemonic JSR ---------------------------------------------------------
      when "01101000" | "01101001" | "01101010" | "01101011" =>
        mnemonic_v   := MN_JSR;
        multi_byte_v := true;

      -- Mnemonic RET ---------------------------------------------------------
      when "01001000" =>
        mnemonic_v   := MN_RET;

      -- Mnemonic RETSK -------------------------------------------------------
      when "01001001" =>
        mnemonic_v   := MN_RETSK;

      -- Mnemonic LD ----------------------------------------------------------
      when "00000101" | "00010101" | "00100101" | "00110101" =>
        mnemonic_v   := MN_LD;

      -- Mnemonic LDD_XAD -----------------------------------------------------
      when "00100011" =>
        mnemonic_v   := MN_LDD_XAD;
        multi_byte_v := true;

      -- Mnemonic LQID --------------------------------------------------------
      when "10111111" =>
        mnemonic_v   := MN_LQID;

      -- Mnemonic RMB ---------------------------------------------------------
      when "01001100" | "01000101" | "01000010" | "01000011" =>
        mnemonic_v   := MN_RMB;

      -- Mnemonic SMB ---------------------------------------------------------
      when "01001101" | "01000111" | "01000110" | "01001011" =>
        mnemonic_v   := MN_SMB;

      -- Mnemonic STII --------------------------------------------------------
      when "01110000" | "01110001" | "01110010" | "01110011" |
           "01110100" | "01110101" | "01110110" | "01110111" |
           "01111000" | "01111001" | "01111010" | "01111011" |
           "01111100" | "01111101" | "01111110" | "01111111" =>
        mnemonic_v   := MN_STII;

      -- Mnemonic X -----------------------------------------------------------
      when "00000110" | "00010110" | "00100110" | "00110110" =>
        mnemonic_v   := MN_X;

      -- Mnemonic XDS ---------------------------------------------------------
      when "00000111" | "00010111" | "00100111" | "00110111" =>
        mnemonic_v   := MN_XDS;

      -- Mnemonic XIS ---------------------------------------------------------
      when "00000100" | "00010100" | "00100100" | "00110100" =>
        mnemonic_v   := MN_XIS;

      -- Mnemonic CAB ---------------------------------------------------------
      when "01010000" =>
        mnemonic_v   := MN_CAB;

      -- Mnemonic CBA ---------------------------------------------------------
      when "01001110" =>
        mnemonic_v   := MN_CBA;

      -- Mnemonic LBI ---------------------------------------------------------
      when "00001000" | "00001001" | "00001010" | "00001011" |
           "00001100" | "00001101" | "00001110" | "00001111" |
           "00011000" | "00011001" | "00011010" | "00011011" |
           "00011100" | "00011101" | "00011110" | "00011111" |
           "00101000" | "00101001" | "00101010" | "00101011" |
           "00101100" | "00101101" | "00101110" | "00101111" |
           "00111000" | "00111001" | "00111010" | "00111011" |
           "00111100" | "00111101" | "00111110" | "00111111" =>
        mnemonic_v   := MN_LBI;

      -- Mnemonic XABR --------------------------------------------------------
      when "00010010" =>
        if not t41x_type_v then
          mnemonic_v := MN_XABR;
        end if;

      -- Mnemonic SKC ---------------------------------------------------------
      when "00100000" =>
        mnemonic_v   := MN_SKC;

      -- Mnemonic SKE ---------------------------------------------------------
      when "00100001" =>
        mnemonic_v   := MN_SKE;

      -- Mnemonic SKMBZ -------------------------------------------------------
      when "00000001" | "00010001" | "00000011" | "00010011" =>
        mnemonic_v   := MN_SKMBZ;

      -- Mnemonic SKT ---------------------------------------------------------
      when "01000001" =>
        if not t41x_type_v then
          mnemonic_v := MN_SKT;
        end if;

      -- Mnemonic XAS ---------------------------------------------------------
      when "01001111" =>
        mnemonic_v   := MN_XAS;

      -- Mnemonic EXT ---------------------------------------------------------
      when "00110011" =>
        mnemonic_v   := MN_EXT;
        multi_byte_v := true;


      when others =>
        null;
    end case;

    result_v.mnemonic   := mnemonic_v;
    result_v.multi_byte := multi_byte_v;

    return result_v;
  end;

end t400_mnemonic_pack;
