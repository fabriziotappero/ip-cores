`define WB2AXI_AXI_ID_W           4
`define WB2AXI_AXI_ADDR_W         32
`define WB2AXI_AXI_DATA_W         32
`define WB2AXI_AXI_PROT_W         3
`define WB2AXI_AXI_STB_W          4
`define WB2AXI_AXI_LEN_W          4
`define WB2AXI_AXI_SIZE_W         3
`define WB2AXI_AXI_BURST_W        2
`define WB2AXI_AXI_LOCK_W         2
`define WB2AXI_AXI_CACHE_W        4
`define WB2AXI_AXI_RESP_W         2

`define WB2AXI_FIFO_ADDR_DEPTH_W  10
`define WB2AXI_FIFO_ADDR_W        64
`define WB2AXI_FIFO_DATA_DEPTH_W  11
`define WB2AXI_FIFO_DATA_W        64
`define WB2AXI_WB_ADR_W           32
`define WB2AXI_WB_DAT_W           32
`define WB2AXI_WB_TGA_W           8
`define WB2AXI_WB_TGD_W           8
`define WB2AXI_WB_TGC_W           4
`define WB2AXI_WB_SEL_W           4
`define WB2AXI_WB_CTI_W           3
`define WB2AXI_WB_BTE_W           2

