-------------------------------------------------------------------------------
--
-- The Interrupt Controller.
-- It collects the interrupt sources and notifies the decoder.
--
-- $Id: int-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_int_rtl_c0 of t48_int is

  for rtl
  end for;

end t48_int_rtl_c0;
