--------------------------------------------------------------------------------
-- 8-Color 100x37 Textmode Video Controller                                   --
--------------------------------------------------------------------------------
--                                                                            --
-- IMPORTANT NOTICE                                                           --
--                                                                            --
-- Data in reverse order and shifted to the left 2px. Saves LUTs. Use the     --
-- python script <chars.py> to generate your customized character set.        --
--                                                                            --
--------------------------------------------------------------------------------
-- Copyright (C)2011  Mathias H�rtnagl <mathias.hoertnagl@gmail.comt>         --
--                                                                            --
-- This program is free software: you can redistribute it and/or modify       --
-- it under the terms of the GNU General Public License as published by       --
-- the Free Software Foundation, either version 3 of the License, or          --
-- (at your option) any later version.                                        --
--                                                                            --
-- This program is distributed in the hope that it will be useful,            --
-- but WITHOUT ANY WARRANTY; without even the implied warranty of             --
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the              --
-- GNU General Public License for more details.                               --
--                                                                            --
-- You should have received a copy of the GNU General Public License          --
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.      --
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
   port(
      clk      : in  std_logic;
      rom_addr : in  std_logic_vector(11 downto 0);
      rom_word : out std_logic_vector(7 downto 0)
   );
end rom;

architecture rtl of rom is
begin
   chrs : process(clk)
   begin
      if rising_edge(clk) then
         case to_integer(unsigned(rom_addr)) is
            when   18 => rom_word <= "11111001";
            when   19 => rom_word <= "00000110";
            when   20 => rom_word <= "10010110";
            when   21 => rom_word <= "00000110";
            when   22 => rom_word <= "00000110";
            when   23 => rom_word <= "11110110";
            when   24 => rom_word <= "01100110";
            when   25 => rom_word <= "00000110";
            when   26 => rom_word <= "00000110";
            when   27 => rom_word <= "11111001";
            when   34 => rom_word <= "11111001";
            when   35 => rom_word <= "11111111";
            when   36 => rom_word <= "01101111";
            when   37 => rom_word <= "11111111";
            when   38 => rom_word <= "11111111";
            when   39 => rom_word <= "00001111";
            when   40 => rom_word <= "10011111";
            when   41 => rom_word <= "11111111";
            when   42 => rom_word <= "11111111";
            when   43 => rom_word <= "11111001";
            when   52 => rom_word <= "11011000";
            when   53 => rom_word <= "11111101";
            when   54 => rom_word <= "11111101";
            when   55 => rom_word <= "11111101";
            when   56 => rom_word <= "11111101";
            when   57 => rom_word <= "11111000";
            when   58 => rom_word <= "01110000";
            when   59 => rom_word <= "00100000";
            when   68 => rom_word <= "00100000";
            when   69 => rom_word <= "01110000";
            when   70 => rom_word <= "11111000";
            when   71 => rom_word <= "11111101";
            when   72 => rom_word <= "11111000";
            when   73 => rom_word <= "01110000";
            when   74 => rom_word <= "00100000";
            when   83 => rom_word <= "01100000";
            when   84 => rom_word <= "11110000";
            when   85 => rom_word <= "11110000";
            when   86 => rom_word <= "10011111";
            when   87 => rom_word <= "10011111";
            when   88 => rom_word <= "10011111";
            when   89 => rom_word <= "01100000";
            when   90 => rom_word <= "01100000";
            when   91 => rom_word <= "11110000";
            when   99 => rom_word <= "01100000";
            when  100 => rom_word <= "11110000";
            when  101 => rom_word <= "11111001";
            when  102 => rom_word <= "11111111";
            when  103 => rom_word <= "11111111";
            when  104 => rom_word <= "11111001";
            when  105 => rom_word <= "01100000";
            when  106 => rom_word <= "01100000";
            when  107 => rom_word <= "11110000";
            when  118 => rom_word <= "01100000";
            when  119 => rom_word <= "11110000";
            when  120 => rom_word <= "11110000";
            when  121 => rom_word <= "01100000";
            when  128 => rom_word <= "11111111";
            when  129 => rom_word <= "11111111";
            when  130 => rom_word <= "11111111";
            when  131 => rom_word <= "11111111";
            when  132 => rom_word <= "11111111";
            when  133 => rom_word <= "11111111";
            when  134 => rom_word <= "10011111";
            when  135 => rom_word <= "00001111";
            when  136 => rom_word <= "00001111";
            when  137 => rom_word <= "10011111";
            when  138 => rom_word <= "11111111";
            when  139 => rom_word <= "11111111";
            when  140 => rom_word <= "11111111";
            when  141 => rom_word <= "11111111";
            when  142 => rom_word <= "11111111";
            when  143 => rom_word <= "11111111";
            when  149 => rom_word <= "11110000";
            when  150 => rom_word <= "10011001";
            when  151 => rom_word <= "00001001";
            when  152 => rom_word <= "00001001";
            when  153 => rom_word <= "10011001";
            when  154 => rom_word <= "11110000";
            when  160 => rom_word <= "11111111";
            when  161 => rom_word <= "11111111";
            when  162 => rom_word <= "11111111";
            when  163 => rom_word <= "11111111";
            when  164 => rom_word <= "11111111";
            when  165 => rom_word <= "00001111";
            when  166 => rom_word <= "01100110";
            when  167 => rom_word <= "11110110";
            when  168 => rom_word <= "11110110";
            when  169 => rom_word <= "01100110";
            when  170 => rom_word <= "00001111";
            when  171 => rom_word <= "11111111";
            when  172 => rom_word <= "11111111";
            when  173 => rom_word <= "11111111";
            when  174 => rom_word <= "11111111";
            when  175 => rom_word <= "11111111";
            when  178 => rom_word <= "11100001";
            when  179 => rom_word <= "11000001";
            when  180 => rom_word <= "01100001";
            when  181 => rom_word <= "00110001";
            when  182 => rom_word <= "01111000";
            when  183 => rom_word <= "11001100";
            when  184 => rom_word <= "11001100";
            when  185 => rom_word <= "11001100";
            when  186 => rom_word <= "11001100";
            when  187 => rom_word <= "01111000";
            when  194 => rom_word <= "11110000";
            when  195 => rom_word <= "10011001";
            when  196 => rom_word <= "10011001";
            when  197 => rom_word <= "10011001";
            when  198 => rom_word <= "10011001";
            when  199 => rom_word <= "11110000";
            when  200 => rom_word <= "01100000";
            when  201 => rom_word <= "11111001";
            when  202 => rom_word <= "01100000";
            when  203 => rom_word <= "01100000";
            when  210 => rom_word <= "11110011";
            when  211 => rom_word <= "00110011";
            when  212 => rom_word <= "11110011";
            when  213 => rom_word <= "00110000";
            when  214 => rom_word <= "00110000";
            when  215 => rom_word <= "00110000";
            when  216 => rom_word <= "00110000";
            when  217 => rom_word <= "00111000";
            when  218 => rom_word <= "00111100";
            when  219 => rom_word <= "00011100";
            when  226 => rom_word <= "11111011";
            when  227 => rom_word <= "00011011";
            when  228 => rom_word <= "11111011";
            when  229 => rom_word <= "00011011";
            when  230 => rom_word <= "00011011";
            when  231 => rom_word <= "00011011";
            when  232 => rom_word <= "00011011";
            when  233 => rom_word <= "10011011";
            when  234 => rom_word <= "10011111";
            when  235 => rom_word <= "10011101";
            when  236 => rom_word <= "00001100";
            when  243 => rom_word <= "01100000";
            when  244 => rom_word <= "01100000";
            when  245 => rom_word <= "01101111";
            when  246 => rom_word <= "11110000";
            when  247 => rom_word <= "10011111";
            when  248 => rom_word <= "11110000";
            when  249 => rom_word <= "01101111";
            when  250 => rom_word <= "01100000";
            when  251 => rom_word <= "01100000";
            when  257 => rom_word <= "00000100";
            when  258 => rom_word <= "00001100";
            when  259 => rom_word <= "00011100";
            when  260 => rom_word <= "00111100";
            when  261 => rom_word <= "01111100";
            when  262 => rom_word <= "11111101";
            when  263 => rom_word <= "01111100";
            when  264 => rom_word <= "00111100";
            when  265 => rom_word <= "00011100";
            when  266 => rom_word <= "00001100";
            when  267 => rom_word <= "00000100";
            when  273 => rom_word <= "00000001";
            when  274 => rom_word <= "10000001";
            when  275 => rom_word <= "11000001";
            when  276 => rom_word <= "11100001";
            when  277 => rom_word <= "11110001";
            when  278 => rom_word <= "11111101";
            when  279 => rom_word <= "11110001";
            when  280 => rom_word <= "11100001";
            when  281 => rom_word <= "11000001";
            when  282 => rom_word <= "10000001";
            when  283 => rom_word <= "00000001";
            when  290 => rom_word <= "01100000";
            when  291 => rom_word <= "11110000";
            when  292 => rom_word <= "11111001";
            when  293 => rom_word <= "01100000";
            when  294 => rom_word <= "01100000";
            when  295 => rom_word <= "01100000";
            when  296 => rom_word <= "11111001";
            when  297 => rom_word <= "11110000";
            when  298 => rom_word <= "01100000";
            when  306 => rom_word <= "10011001";
            when  307 => rom_word <= "10011001";
            when  308 => rom_word <= "10011001";
            when  309 => rom_word <= "10011001";
            when  310 => rom_word <= "10011001";
            when  311 => rom_word <= "10011001";
            when  312 => rom_word <= "10011001";
            when  314 => rom_word <= "10011001";
            when  315 => rom_word <= "10011001";
            when  322 => rom_word <= "11111011";
            when  323 => rom_word <= "01101111";
            when  324 => rom_word <= "01101111";
            when  325 => rom_word <= "01101111";
            when  326 => rom_word <= "01111011";
            when  327 => rom_word <= "01100011";
            when  328 => rom_word <= "01100011";
            when  329 => rom_word <= "01100011";
            when  330 => rom_word <= "01100011";
            when  331 => rom_word <= "01100011";
            when  337 => rom_word <= "11111000";
            when  338 => rom_word <= "10001101";
            when  339 => rom_word <= "00011000";
            when  340 => rom_word <= "01110000";
            when  341 => rom_word <= "11011000";
            when  342 => rom_word <= "10001101";
            when  343 => rom_word <= "10001101";
            when  344 => rom_word <= "11011000";
            when  345 => rom_word <= "01110000";
            when  346 => rom_word <= "11000000";
            when  347 => rom_word <= "10001101";
            when  348 => rom_word <= "11111000";
            when  360 => rom_word <= "11111101";
            when  361 => rom_word <= "11111101";
            when  362 => rom_word <= "11111101";
            when  363 => rom_word <= "11111101";
            when  370 => rom_word <= "01100000";
            when  371 => rom_word <= "11110000";
            when  372 => rom_word <= "11111001";
            when  373 => rom_word <= "01100000";
            when  374 => rom_word <= "01100000";
            when  375 => rom_word <= "01100000";
            when  376 => rom_word <= "11111001";
            when  377 => rom_word <= "11110000";
            when  378 => rom_word <= "01100000";
            when  379 => rom_word <= "11111001";
            when  386 => rom_word <= "01100000";
            when  387 => rom_word <= "11110000";
            when  388 => rom_word <= "11111001";
            when  389 => rom_word <= "01100000";
            when  390 => rom_word <= "01100000";
            when  391 => rom_word <= "01100000";
            when  392 => rom_word <= "01100000";
            when  393 => rom_word <= "01100000";
            when  394 => rom_word <= "01100000";
            when  395 => rom_word <= "01100000";
            when  402 => rom_word <= "01100000";
            when  403 => rom_word <= "01100000";
            when  404 => rom_word <= "01100000";
            when  405 => rom_word <= "01100000";
            when  406 => rom_word <= "01100000";
            when  407 => rom_word <= "01100000";
            when  408 => rom_word <= "01100000";
            when  409 => rom_word <= "11111001";
            when  410 => rom_word <= "11110000";
            when  411 => rom_word <= "01100000";
            when  421 => rom_word <= "01100000";
            when  422 => rom_word <= "11000000";
            when  423 => rom_word <= "11111101";
            when  424 => rom_word <= "11000000";
            when  425 => rom_word <= "01100000";
            when  437 => rom_word <= "00110000";
            when  438 => rom_word <= "00011000";
            when  439 => rom_word <= "11111101";
            when  440 => rom_word <= "00011000";
            when  441 => rom_word <= "00110000";
            when  454 => rom_word <= "00001100";
            when  455 => rom_word <= "00001100";
            when  456 => rom_word <= "00001100";
            when  457 => rom_word <= "11111101";
            when  469 => rom_word <= "01010000";
            when  470 => rom_word <= "11011000";
            when  471 => rom_word <= "11111101";
            when  472 => rom_word <= "11011000";
            when  473 => rom_word <= "01010000";
            when  484 => rom_word <= "00100000";
            when  485 => rom_word <= "01110000";
            when  486 => rom_word <= "01110000";
            when  487 => rom_word <= "11111000";
            when  488 => rom_word <= "11111000";
            when  489 => rom_word <= "11111101";
            when  490 => rom_word <= "11111101";
            when  500 => rom_word <= "11111101";
            when  501 => rom_word <= "11111101";
            when  502 => rom_word <= "11111000";
            when  503 => rom_word <= "11111000";
            when  504 => rom_word <= "01110000";
            when  505 => rom_word <= "01110000";
            when  506 => rom_word <= "00100000";
            when  530 => rom_word <= "01100000";
            when  531 => rom_word <= "11110000";
            when  532 => rom_word <= "11110000";
            when  533 => rom_word <= "11110000";
            when  534 => rom_word <= "01100000";
            when  535 => rom_word <= "01100000";
            when  536 => rom_word <= "01100000";
            when  538 => rom_word <= "01100000";
            when  539 => rom_word <= "01100000";
            when  545 => rom_word <= "10011001";
            when  546 => rom_word <= "10011001";
            when  547 => rom_word <= "10011001";
            when  548 => rom_word <= "10010000";
            when  563 => rom_word <= "11011000";
            when  564 => rom_word <= "11011000";
            when  565 => rom_word <= "11111101";
            when  566 => rom_word <= "11011000";
            when  567 => rom_word <= "11011000";
            when  568 => rom_word <= "11011000";
            when  569 => rom_word <= "11111101";
            when  570 => rom_word <= "11011000";
            when  571 => rom_word <= "11011000";
            when  576 => rom_word <= "01100000";
            when  577 => rom_word <= "01100000";
            when  578 => rom_word <= "11111000";
            when  579 => rom_word <= "10001101";
            when  580 => rom_word <= "00001101";
            when  581 => rom_word <= "00001100";
            when  582 => rom_word <= "11111000";
            when  583 => rom_word <= "10000001";
            when  584 => rom_word <= "10000001";
            when  585 => rom_word <= "10000101";
            when  586 => rom_word <= "10001101";
            when  587 => rom_word <= "11111000";
            when  588 => rom_word <= "01100000";
            when  589 => rom_word <= "01100000";
            when  596 => rom_word <= "00001101";
            when  597 => rom_word <= "10001101";
            when  598 => rom_word <= "11000000";
            when  599 => rom_word <= "01100000";
            when  600 => rom_word <= "00110000";
            when  601 => rom_word <= "00011000";
            when  602 => rom_word <= "10001101";
            when  603 => rom_word <= "10000101";
            when  610 => rom_word <= "01110000";
            when  611 => rom_word <= "11011000";
            when  612 => rom_word <= "11011000";
            when  613 => rom_word <= "01110000";
            when  614 => rom_word <= "10111001";
            when  615 => rom_word <= "11101100";
            when  616 => rom_word <= "11001100";
            when  617 => rom_word <= "11001100";
            when  618 => rom_word <= "11001100";
            when  619 => rom_word <= "10111001";
            when  625 => rom_word <= "00110000";
            when  626 => rom_word <= "00110000";
            when  627 => rom_word <= "00110000";
            when  628 => rom_word <= "00011000";
            when  642 => rom_word <= "11000000";
            when  643 => rom_word <= "01100000";
            when  644 => rom_word <= "00110000";
            when  645 => rom_word <= "00110000";
            when  646 => rom_word <= "00110000";
            when  647 => rom_word <= "00110000";
            when  648 => rom_word <= "00110000";
            when  649 => rom_word <= "00110000";
            when  650 => rom_word <= "01100000";
            when  651 => rom_word <= "11000000";
            when  658 => rom_word <= "00110000";
            when  659 => rom_word <= "01100000";
            when  660 => rom_word <= "11000000";
            when  661 => rom_word <= "11000000";
            when  662 => rom_word <= "11000000";
            when  663 => rom_word <= "11000000";
            when  664 => rom_word <= "11000000";
            when  665 => rom_word <= "11000000";
            when  666 => rom_word <= "01100000";
            when  667 => rom_word <= "00110000";
            when  677 => rom_word <= "10011001";
            when  678 => rom_word <= "11110000";
            when  679 => rom_word <= "11111111";
            when  680 => rom_word <= "11110000";
            when  681 => rom_word <= "10011001";
            when  693 => rom_word <= "01100000";
            when  694 => rom_word <= "01100000";
            when  695 => rom_word <= "11111001";
            when  696 => rom_word <= "01100000";
            when  697 => rom_word <= "01100000";
            when  713 => rom_word <= "01100000";
            when  714 => rom_word <= "01100000";
            when  715 => rom_word <= "01100000";
            when  716 => rom_word <= "00110000";
            when  727 => rom_word <= "11111101";
            when  746 => rom_word <= "01100000";
            when  747 => rom_word <= "01100000";
            when  756 => rom_word <= "00000001";
            when  757 => rom_word <= "10000001";
            when  758 => rom_word <= "11000000";
            when  759 => rom_word <= "01100000";
            when  760 => rom_word <= "00110000";
            when  761 => rom_word <= "00011000";
            when  762 => rom_word <= "00001100";
            when  763 => rom_word <= "00000100";
            when  770 => rom_word <= "01110000";
            when  771 => rom_word <= "11011000";
            when  772 => rom_word <= "10001101";
            when  773 => rom_word <= "11001101";
            when  774 => rom_word <= "11101101";
            when  775 => rom_word <= "10111101";
            when  776 => rom_word <= "10011101";
            when  777 => rom_word <= "10001101";
            when  778 => rom_word <= "11011000";
            when  779 => rom_word <= "01110000";
            when  786 => rom_word <= "01100000";
            when  787 => rom_word <= "01110000";
            when  788 => rom_word <= "01111000";
            when  789 => rom_word <= "01100000";
            when  790 => rom_word <= "01100000";
            when  791 => rom_word <= "01100000";
            when  792 => rom_word <= "01100000";
            when  793 => rom_word <= "01100000";
            when  794 => rom_word <= "01100000";
            when  795 => rom_word <= "01100000";
            when  802 => rom_word <= "11111000";
            when  803 => rom_word <= "10001101";
            when  804 => rom_word <= "10000001";
            when  805 => rom_word <= "11000000";
            when  806 => rom_word <= "01100000";
            when  807 => rom_word <= "00110000";
            when  808 => rom_word <= "00011000";
            when  809 => rom_word <= "00001100";
            when  810 => rom_word <= "00001100";
            when  811 => rom_word <= "11111101";
            when  818 => rom_word <= "11111000";
            when  819 => rom_word <= "10000101";
            when  820 => rom_word <= "10000001";
            when  821 => rom_word <= "10000001";
            when  822 => rom_word <= "11110000";
            when  823 => rom_word <= "10000001";
            when  824 => rom_word <= "10000001";
            when  825 => rom_word <= "10000001";
            when  826 => rom_word <= "10000101";
            when  827 => rom_word <= "11111000";
            when  834 => rom_word <= "11000000";
            when  835 => rom_word <= "11100000";
            when  836 => rom_word <= "11110000";
            when  837 => rom_word <= "11011000";
            when  838 => rom_word <= "11001100";
            when  839 => rom_word <= "11111101";
            when  840 => rom_word <= "11000000";
            when  841 => rom_word <= "11000000";
            when  842 => rom_word <= "11000000";
            when  843 => rom_word <= "11000000";
            when  850 => rom_word <= "11111101";
            when  851 => rom_word <= "00001100";
            when  852 => rom_word <= "00001100";
            when  853 => rom_word <= "00001100";
            when  854 => rom_word <= "11111100";
            when  855 => rom_word <= "10000001";
            when  856 => rom_word <= "10000001";
            when  857 => rom_word <= "10000001";
            when  858 => rom_word <= "10000101";
            when  859 => rom_word <= "11111000";
            when  866 => rom_word <= "11110000";
            when  867 => rom_word <= "00011000";
            when  868 => rom_word <= "00001100";
            when  869 => rom_word <= "00001100";
            when  870 => rom_word <= "11101100";
            when  871 => rom_word <= "10011101";
            when  872 => rom_word <= "10001101";
            when  873 => rom_word <= "10001101";
            when  874 => rom_word <= "10001101";
            when  875 => rom_word <= "11111000";
            when  882 => rom_word <= "11111101";
            when  883 => rom_word <= "10000001";
            when  884 => rom_word <= "10000001";
            when  885 => rom_word <= "10000001";
            when  886 => rom_word <= "11000000";
            when  887 => rom_word <= "01100000";
            when  888 => rom_word <= "00110000";
            when  889 => rom_word <= "00110000";
            when  890 => rom_word <= "00110000";
            when  891 => rom_word <= "00110000";
            when  898 => rom_word <= "11111000";
            when  899 => rom_word <= "10001101";
            when  900 => rom_word <= "10001101";
            when  901 => rom_word <= "10001101";
            when  902 => rom_word <= "11111000";
            when  903 => rom_word <= "10001101";
            when  904 => rom_word <= "10001101";
            when  905 => rom_word <= "10001101";
            when  906 => rom_word <= "10001101";
            when  907 => rom_word <= "11111000";
            when  914 => rom_word <= "11111000";
            when  915 => rom_word <= "10001101";
            when  916 => rom_word <= "10001101";
            when  917 => rom_word <= "10001101";
            when  918 => rom_word <= "11111001";
            when  919 => rom_word <= "10000001";
            when  920 => rom_word <= "10000001";
            when  921 => rom_word <= "10000001";
            when  922 => rom_word <= "11000100";
            when  923 => rom_word <= "01111000";
            when  932 => rom_word <= "01100000";
            when  933 => rom_word <= "01100000";
            when  937 => rom_word <= "01100000";
            when  938 => rom_word <= "01100000";
            when  948 => rom_word <= "01100000";
            when  949 => rom_word <= "01100000";
            when  953 => rom_word <= "01100000";
            when  954 => rom_word <= "01100000";
            when  955 => rom_word <= "00110000";
            when  963 => rom_word <= "10000001";
            when  964 => rom_word <= "11000000";
            when  965 => rom_word <= "01100000";
            when  966 => rom_word <= "00110000";
            when  967 => rom_word <= "00011000";
            when  968 => rom_word <= "00110000";
            when  969 => rom_word <= "01100000";
            when  970 => rom_word <= "11000000";
            when  971 => rom_word <= "10000001";
            when  981 => rom_word <= "11111001";
            when  984 => rom_word <= "11111001";
            when  995 => rom_word <= "00011000";
            when  996 => rom_word <= "00110000";
            when  997 => rom_word <= "01100000";
            when  998 => rom_word <= "11000000";
            when  999 => rom_word <= "10000001";
            when 1000 => rom_word <= "11000000";
            when 1001 => rom_word <= "01100000";
            when 1002 => rom_word <= "00110000";
            when 1003 => rom_word <= "00011000";
            when 1010 => rom_word <= "11111000";
            when 1011 => rom_word <= "10001101";
            when 1012 => rom_word <= "10001101";
            when 1013 => rom_word <= "11000000";
            when 1014 => rom_word <= "01100000";
            when 1015 => rom_word <= "01100000";
            when 1016 => rom_word <= "01100000";
            when 1018 => rom_word <= "01100000";
            when 1019 => rom_word <= "01100000";
            when 1027 => rom_word <= "11111000";
            when 1028 => rom_word <= "10001101";
            when 1029 => rom_word <= "10001101";
            when 1030 => rom_word <= "11101101";
            when 1031 => rom_word <= "11101101";
            when 1032 => rom_word <= "11101101";
            when 1033 => rom_word <= "11101100";
            when 1034 => rom_word <= "00001100";
            when 1035 => rom_word <= "11111000";
            when 1042 => rom_word <= "00100000";
            when 1043 => rom_word <= "01110000";
            when 1044 => rom_word <= "11011000";
            when 1045 => rom_word <= "10001101";
            when 1046 => rom_word <= "10001101";
            when 1047 => rom_word <= "11111101";
            when 1048 => rom_word <= "10001101";
            when 1049 => rom_word <= "10001101";
            when 1050 => rom_word <= "10001101";
            when 1051 => rom_word <= "10001101";
            when 1058 => rom_word <= "11111100";
            when 1059 => rom_word <= "10001101";
            when 1060 => rom_word <= "10001101";
            when 1061 => rom_word <= "10001101";
            when 1062 => rom_word <= "11111100";
            when 1063 => rom_word <= "10001101";
            when 1064 => rom_word <= "10001101";
            when 1065 => rom_word <= "10001101";
            when 1066 => rom_word <= "10001101";
            when 1067 => rom_word <= "11111100";
            when 1074 => rom_word <= "11110000";
            when 1075 => rom_word <= "10011001";
            when 1076 => rom_word <= "00001101";
            when 1077 => rom_word <= "00001100";
            when 1078 => rom_word <= "00001100";
            when 1079 => rom_word <= "00001100";
            when 1080 => rom_word <= "00001100";
            when 1081 => rom_word <= "00001101";
            when 1082 => rom_word <= "10011001";
            when 1083 => rom_word <= "11110000";
            when 1090 => rom_word <= "01111100";
            when 1091 => rom_word <= "11101100";
            when 1092 => rom_word <= "11001101";
            when 1093 => rom_word <= "10001101";
            when 1094 => rom_word <= "10001101";
            when 1095 => rom_word <= "10001101";
            when 1096 => rom_word <= "10001101";
            when 1097 => rom_word <= "11001101";
            when 1098 => rom_word <= "11101100";
            when 1099 => rom_word <= "01111100";
            when 1106 => rom_word <= "11111100";
            when 1107 => rom_word <= "00001100";
            when 1108 => rom_word <= "00001100";
            when 1109 => rom_word <= "00001100";
            when 1110 => rom_word <= "01111100";
            when 1111 => rom_word <= "00001100";
            when 1112 => rom_word <= "00001100";
            when 1113 => rom_word <= "00001100";
            when 1114 => rom_word <= "00001100";
            when 1115 => rom_word <= "11111100";
            when 1122 => rom_word <= "11111100";
            when 1123 => rom_word <= "00001100";
            when 1124 => rom_word <= "00001100";
            when 1125 => rom_word <= "00001100";
            when 1126 => rom_word <= "01111100";
            when 1127 => rom_word <= "00001100";
            when 1128 => rom_word <= "00001100";
            when 1129 => rom_word <= "00001100";
            when 1130 => rom_word <= "00001100";
            when 1131 => rom_word <= "00001100";
            when 1138 => rom_word <= "11110000";
            when 1139 => rom_word <= "00011001";
            when 1140 => rom_word <= "00001100";
            when 1141 => rom_word <= "00001100";
            when 1142 => rom_word <= "00001100";
            when 1143 => rom_word <= "11101101";
            when 1144 => rom_word <= "10001101";
            when 1145 => rom_word <= "10001101";
            when 1146 => rom_word <= "10011001";
            when 1147 => rom_word <= "11110001";
            when 1154 => rom_word <= "10001101";
            when 1155 => rom_word <= "10001101";
            when 1156 => rom_word <= "10001101";
            when 1157 => rom_word <= "10001101";
            when 1158 => rom_word <= "11111101";
            when 1159 => rom_word <= "10001101";
            when 1160 => rom_word <= "10001101";
            when 1161 => rom_word <= "10001101";
            when 1162 => rom_word <= "10001101";
            when 1163 => rom_word <= "10001101";
            when 1170 => rom_word <= "01100000";
            when 1171 => rom_word <= "01100000";
            when 1172 => rom_word <= "01100000";
            when 1173 => rom_word <= "01100000";
            when 1174 => rom_word <= "01100000";
            when 1175 => rom_word <= "01100000";
            when 1176 => rom_word <= "01100000";
            when 1177 => rom_word <= "01100000";
            when 1178 => rom_word <= "01100000";
            when 1179 => rom_word <= "01100000";
            when 1186 => rom_word <= "11100001";
            when 1187 => rom_word <= "11000000";
            when 1188 => rom_word <= "11000000";
            when 1189 => rom_word <= "11000000";
            when 1190 => rom_word <= "11000000";
            when 1191 => rom_word <= "11000000";
            when 1192 => rom_word <= "11001100";
            when 1193 => rom_word <= "11001100";
            when 1194 => rom_word <= "11001100";
            when 1195 => rom_word <= "01111000";
            when 1202 => rom_word <= "00001101";
            when 1203 => rom_word <= "10001101";
            when 1204 => rom_word <= "11001100";
            when 1205 => rom_word <= "01101100";
            when 1206 => rom_word <= "00111100";
            when 1207 => rom_word <= "00111100";
            when 1208 => rom_word <= "01101100";
            when 1209 => rom_word <= "11001100";
            when 1210 => rom_word <= "10001101";
            when 1211 => rom_word <= "00001101";
            when 1218 => rom_word <= "00001100";
            when 1219 => rom_word <= "00001100";
            when 1220 => rom_word <= "00001100";
            when 1221 => rom_word <= "00001100";
            when 1222 => rom_word <= "00001100";
            when 1223 => rom_word <= "00001100";
            when 1224 => rom_word <= "00001100";
            when 1225 => rom_word <= "00001100";
            when 1226 => rom_word <= "00001100";
            when 1227 => rom_word <= "11111100";
            when 1234 => rom_word <= "10001101";
            when 1235 => rom_word <= "11011101";
            when 1236 => rom_word <= "11111101";
            when 1237 => rom_word <= "11111101";
            when 1238 => rom_word <= "10101101";
            when 1239 => rom_word <= "10001101";
            when 1240 => rom_word <= "10001101";
            when 1241 => rom_word <= "10001101";
            when 1242 => rom_word <= "10001101";
            when 1243 => rom_word <= "10001101";
            when 1250 => rom_word <= "10001101";
            when 1251 => rom_word <= "10011101";
            when 1252 => rom_word <= "10111101";
            when 1253 => rom_word <= "11111101";
            when 1254 => rom_word <= "11101101";
            when 1255 => rom_word <= "11001101";
            when 1256 => rom_word <= "10001101";
            when 1257 => rom_word <= "10001101";
            when 1258 => rom_word <= "10001101";
            when 1259 => rom_word <= "10001101";
            when 1266 => rom_word <= "11111000";
            when 1267 => rom_word <= "10001101";
            when 1268 => rom_word <= "10001101";
            when 1269 => rom_word <= "10001101";
            when 1270 => rom_word <= "10001101";
            when 1271 => rom_word <= "10001101";
            when 1272 => rom_word <= "10001101";
            when 1273 => rom_word <= "10001101";
            when 1274 => rom_word <= "10001101";
            when 1275 => rom_word <= "11111000";
            when 1282 => rom_word <= "11111100";
            when 1283 => rom_word <= "10001101";
            when 1284 => rom_word <= "10001101";
            when 1285 => rom_word <= "10001101";
            when 1286 => rom_word <= "11111100";
            when 1287 => rom_word <= "00001100";
            when 1288 => rom_word <= "00001100";
            when 1289 => rom_word <= "00001100";
            when 1290 => rom_word <= "00001100";
            when 1291 => rom_word <= "00001100";
            when 1298 => rom_word <= "11111000";
            when 1299 => rom_word <= "10001101";
            when 1300 => rom_word <= "10001101";
            when 1301 => rom_word <= "10001101";
            when 1302 => rom_word <= "10001101";
            when 1303 => rom_word <= "10001101";
            when 1304 => rom_word <= "10001101";
            when 1305 => rom_word <= "10101101";
            when 1306 => rom_word <= "11101101";
            when 1307 => rom_word <= "11111000";
            when 1308 => rom_word <= "11000000";
            when 1309 => rom_word <= "10000001";
            when 1314 => rom_word <= "11111100";
            when 1315 => rom_word <= "10001101";
            when 1316 => rom_word <= "10001101";
            when 1317 => rom_word <= "10001101";
            when 1318 => rom_word <= "11111100";
            when 1319 => rom_word <= "01101100";
            when 1320 => rom_word <= "11001100";
            when 1321 => rom_word <= "11001100";
            when 1322 => rom_word <= "10001101";
            when 1323 => rom_word <= "10001101";
            when 1330 => rom_word <= "11111000";
            when 1331 => rom_word <= "00001101";
            when 1332 => rom_word <= "00001100";
            when 1333 => rom_word <= "00011000";
            when 1334 => rom_word <= "01110000";
            when 1335 => rom_word <= "11000000";
            when 1336 => rom_word <= "10000001";
            when 1337 => rom_word <= "10000001";
            when 1338 => rom_word <= "10000101";
            when 1339 => rom_word <= "11111000";
            when 1346 => rom_word <= "11111001";
            when 1347 => rom_word <= "11111001";
            when 1348 => rom_word <= "01100000";
            when 1349 => rom_word <= "01100000";
            when 1350 => rom_word <= "01100000";
            when 1351 => rom_word <= "01100000";
            when 1352 => rom_word <= "01100000";
            when 1353 => rom_word <= "01100000";
            when 1354 => rom_word <= "01100000";
            when 1355 => rom_word <= "01100000";
            when 1362 => rom_word <= "10001101";
            when 1363 => rom_word <= "10001101";
            when 1364 => rom_word <= "10001101";
            when 1365 => rom_word <= "10001101";
            when 1366 => rom_word <= "10001101";
            when 1367 => rom_word <= "10001101";
            when 1368 => rom_word <= "10001101";
            when 1369 => rom_word <= "10001101";
            when 1370 => rom_word <= "10001101";
            when 1371 => rom_word <= "11111000";
            when 1378 => rom_word <= "10001101";
            when 1379 => rom_word <= "10001101";
            when 1380 => rom_word <= "10001101";
            when 1381 => rom_word <= "10001101";
            when 1382 => rom_word <= "10001101";
            when 1383 => rom_word <= "10001101";
            when 1384 => rom_word <= "10001101";
            when 1385 => rom_word <= "11011000";
            when 1386 => rom_word <= "01110000";
            when 1387 => rom_word <= "00100000";
            when 1394 => rom_word <= "10001101";
            when 1395 => rom_word <= "10001101";
            when 1396 => rom_word <= "10001101";
            when 1397 => rom_word <= "10001101";
            when 1398 => rom_word <= "10101101";
            when 1399 => rom_word <= "10101101";
            when 1400 => rom_word <= "10101101";
            when 1401 => rom_word <= "11111101";
            when 1402 => rom_word <= "11011101";
            when 1403 => rom_word <= "11011000";
            when 1410 => rom_word <= "10001101";
            when 1411 => rom_word <= "10001101";
            when 1412 => rom_word <= "11011000";
            when 1413 => rom_word <= "11111000";
            when 1414 => rom_word <= "01110000";
            when 1415 => rom_word <= "01110000";
            when 1416 => rom_word <= "11111000";
            when 1417 => rom_word <= "11011000";
            when 1418 => rom_word <= "10001101";
            when 1419 => rom_word <= "10001101";
            when 1426 => rom_word <= "10011001";
            when 1427 => rom_word <= "10011001";
            when 1428 => rom_word <= "10011001";
            when 1429 => rom_word <= "10011001";
            when 1430 => rom_word <= "11110000";
            when 1431 => rom_word <= "01100000";
            when 1432 => rom_word <= "01100000";
            when 1433 => rom_word <= "01100000";
            when 1434 => rom_word <= "01100000";
            when 1435 => rom_word <= "01100000";
            when 1442 => rom_word <= "11111101";
            when 1443 => rom_word <= "10000001";
            when 1444 => rom_word <= "10000001";
            when 1445 => rom_word <= "11000000";
            when 1446 => rom_word <= "01100000";
            when 1447 => rom_word <= "00110000";
            when 1448 => rom_word <= "00011000";
            when 1449 => rom_word <= "00001100";
            when 1450 => rom_word <= "00001100";
            when 1451 => rom_word <= "11111101";
            when 1458 => rom_word <= "11110000";
            when 1459 => rom_word <= "00110000";
            when 1460 => rom_word <= "00110000";
            when 1461 => rom_word <= "00110000";
            when 1462 => rom_word <= "00110000";
            when 1463 => rom_word <= "00110000";
            when 1464 => rom_word <= "00110000";
            when 1465 => rom_word <= "00110000";
            when 1466 => rom_word <= "00110000";
            when 1467 => rom_word <= "11110000";
            when 1475 => rom_word <= "00000100";
            when 1476 => rom_word <= "00001100";
            when 1477 => rom_word <= "00011100";
            when 1478 => rom_word <= "00111000";
            when 1479 => rom_word <= "01110000";
            when 1480 => rom_word <= "11100000";
            when 1481 => rom_word <= "11000001";
            when 1482 => rom_word <= "10000001";
            when 1483 => rom_word <= "00000001";
            when 1490 => rom_word <= "11110000";
            when 1491 => rom_word <= "11000000";
            when 1492 => rom_word <= "11000000";
            when 1493 => rom_word <= "11000000";
            when 1494 => rom_word <= "11000000";
            when 1495 => rom_word <= "11000000";
            when 1496 => rom_word <= "11000000";
            when 1497 => rom_word <= "11000000";
            when 1498 => rom_word <= "11000000";
            when 1499 => rom_word <= "11110000";
            when 1504 => rom_word <= "00100000";
            when 1505 => rom_word <= "01110000";
            when 1506 => rom_word <= "11011000";
            when 1507 => rom_word <= "10001101";
            when 1533 => rom_word <= "11111111";
            when 1537 => rom_word <= "00110000";
            when 1538 => rom_word <= "01100000";
            when 1539 => rom_word <= "11000000";
            when 1557 => rom_word <= "01111000";
            when 1558 => rom_word <= "11000000";
            when 1559 => rom_word <= "11111000";
            when 1560 => rom_word <= "11001100";
            when 1561 => rom_word <= "11001100";
            when 1562 => rom_word <= "11001100";
            when 1563 => rom_word <= "10111001";
            when 1570 => rom_word <= "00001100";
            when 1571 => rom_word <= "00001100";
            when 1572 => rom_word <= "00001100";
            when 1573 => rom_word <= "01111100";
            when 1574 => rom_word <= "11001100";
            when 1575 => rom_word <= "11001100";
            when 1576 => rom_word <= "11001100";
            when 1577 => rom_word <= "11001100";
            when 1578 => rom_word <= "11001100";
            when 1579 => rom_word <= "01111100";
            when 1589 => rom_word <= "01111000";
            when 1590 => rom_word <= "10001100";
            when 1591 => rom_word <= "00001100";
            when 1592 => rom_word <= "00001100";
            when 1593 => rom_word <= "00001100";
            when 1594 => rom_word <= "10001100";
            when 1595 => rom_word <= "01111000";
            when 1602 => rom_word <= "11000000";
            when 1603 => rom_word <= "11000000";
            when 1604 => rom_word <= "11000000";
            when 1605 => rom_word <= "11111000";
            when 1606 => rom_word <= "11001100";
            when 1607 => rom_word <= "11001100";
            when 1608 => rom_word <= "11001100";
            when 1609 => rom_word <= "11001100";
            when 1610 => rom_word <= "11001100";
            when 1611 => rom_word <= "11111000";
            when 1621 => rom_word <= "11111000";
            when 1622 => rom_word <= "10001101";
            when 1623 => rom_word <= "11111101";
            when 1624 => rom_word <= "00001100";
            when 1625 => rom_word <= "00001100";
            when 1626 => rom_word <= "00001101";
            when 1627 => rom_word <= "11111000";
            when 1634 => rom_word <= "11100000";
            when 1635 => rom_word <= "10110001";
            when 1636 => rom_word <= "00110001";
            when 1637 => rom_word <= "00110000";
            when 1638 => rom_word <= "01111000";
            when 1639 => rom_word <= "00110000";
            when 1640 => rom_word <= "00110000";
            when 1641 => rom_word <= "00110000";
            when 1642 => rom_word <= "00110000";
            when 1643 => rom_word <= "00110000";
            when 1653 => rom_word <= "11111000";
            when 1654 => rom_word <= "11001100";
            when 1655 => rom_word <= "11001100";
            when 1656 => rom_word <= "11001100";
            when 1657 => rom_word <= "11001100";
            when 1658 => rom_word <= "11001100";
            when 1659 => rom_word <= "11111000";
            when 1660 => rom_word <= "11000000";
            when 1661 => rom_word <= "11000100";
            when 1662 => rom_word <= "01111000";
            when 1666 => rom_word <= "00001100";
            when 1667 => rom_word <= "00001100";
            when 1668 => rom_word <= "00001100";
            when 1669 => rom_word <= "01101100";
            when 1670 => rom_word <= "11011100";
            when 1671 => rom_word <= "11001100";
            when 1672 => rom_word <= "11001100";
            when 1673 => rom_word <= "11001100";
            when 1674 => rom_word <= "11001100";
            when 1675 => rom_word <= "11001100";
            when 1682 => rom_word <= "01100000";
            when 1683 => rom_word <= "01100000";
            when 1685 => rom_word <= "01110000";
            when 1686 => rom_word <= "01100000";
            when 1687 => rom_word <= "01100000";
            when 1688 => rom_word <= "01100000";
            when 1689 => rom_word <= "01100000";
            when 1690 => rom_word <= "01100000";
            when 1691 => rom_word <= "01100000";
            when 1698 => rom_word <= "11000000";
            when 1699 => rom_word <= "11000000";
            when 1701 => rom_word <= "11000000";
            when 1702 => rom_word <= "11000000";
            when 1703 => rom_word <= "11000000";
            when 1704 => rom_word <= "11000000";
            when 1705 => rom_word <= "11000000";
            when 1706 => rom_word <= "11000000";
            when 1707 => rom_word <= "11000000";
            when 1708 => rom_word <= "11001100";
            when 1709 => rom_word <= "11001100";
            when 1710 => rom_word <= "01111000";
            when 1714 => rom_word <= "00001100";
            when 1715 => rom_word <= "00001100";
            when 1716 => rom_word <= "00001100";
            when 1717 => rom_word <= "11001100";
            when 1718 => rom_word <= "01101100";
            when 1719 => rom_word <= "00111100";
            when 1720 => rom_word <= "00111100";
            when 1721 => rom_word <= "01101100";
            when 1722 => rom_word <= "11001100";
            when 1723 => rom_word <= "11001100";
            when 1730 => rom_word <= "01110000";
            when 1731 => rom_word <= "01100000";
            when 1732 => rom_word <= "01100000";
            when 1733 => rom_word <= "01100000";
            when 1734 => rom_word <= "01100000";
            when 1735 => rom_word <= "01100000";
            when 1736 => rom_word <= "01100000";
            when 1737 => rom_word <= "01100000";
            when 1738 => rom_word <= "01100000";
            when 1739 => rom_word <= "01100000";
            when 1749 => rom_word <= "11011100";
            when 1750 => rom_word <= "11111101";
            when 1751 => rom_word <= "10101101";
            when 1752 => rom_word <= "10101101";
            when 1753 => rom_word <= "10101101";
            when 1754 => rom_word <= "10101101";
            when 1755 => rom_word <= "10001101";
            when 1765 => rom_word <= "01110100";
            when 1766 => rom_word <= "11001100";
            when 1767 => rom_word <= "11001100";
            when 1768 => rom_word <= "11001100";
            when 1769 => rom_word <= "11001100";
            when 1770 => rom_word <= "11001100";
            when 1771 => rom_word <= "11001100";
            when 1781 => rom_word <= "01111000";
            when 1782 => rom_word <= "11001100";
            when 1783 => rom_word <= "11001100";
            when 1784 => rom_word <= "11001100";
            when 1785 => rom_word <= "11001100";
            when 1786 => rom_word <= "11001100";
            when 1787 => rom_word <= "01111000";
            when 1797 => rom_word <= "01111100";
            when 1798 => rom_word <= "11001100";
            when 1799 => rom_word <= "11001100";
            when 1800 => rom_word <= "11001100";
            when 1801 => rom_word <= "11001100";
            when 1802 => rom_word <= "11001100";
            when 1803 => rom_word <= "01111100";
            when 1804 => rom_word <= "00001100";
            when 1805 => rom_word <= "00001100";
            when 1806 => rom_word <= "00001100";
            when 1813 => rom_word <= "11111000";
            when 1814 => rom_word <= "11001100";
            when 1815 => rom_word <= "11001100";
            when 1816 => rom_word <= "11001100";
            when 1817 => rom_word <= "11001100";
            when 1818 => rom_word <= "11001100";
            when 1819 => rom_word <= "11111000";
            when 1820 => rom_word <= "11000000";
            when 1821 => rom_word <= "11000000";
            when 1822 => rom_word <= "11000000";
            when 1829 => rom_word <= "01110100";
            when 1830 => rom_word <= "11011100";
            when 1831 => rom_word <= "11001100";
            when 1832 => rom_word <= "00001100";
            when 1833 => rom_word <= "00001100";
            when 1834 => rom_word <= "00001100";
            when 1835 => rom_word <= "00001100";
            when 1845 => rom_word <= "11111000";
            when 1846 => rom_word <= "00001101";
            when 1847 => rom_word <= "00111000";
            when 1848 => rom_word <= "11100000";
            when 1849 => rom_word <= "10000001";
            when 1850 => rom_word <= "10000101";
            when 1851 => rom_word <= "11111000";
            when 1858 => rom_word <= "00110000";
            when 1859 => rom_word <= "00110000";
            when 1860 => rom_word <= "00110000";
            when 1861 => rom_word <= "11111100";
            when 1862 => rom_word <= "00110000";
            when 1863 => rom_word <= "00110000";
            when 1864 => rom_word <= "00110000";
            when 1865 => rom_word <= "00110000";
            when 1866 => rom_word <= "00110000";
            when 1867 => rom_word <= "00110000";
            when 1877 => rom_word <= "11001100";
            when 1878 => rom_word <= "11001100";
            when 1879 => rom_word <= "11001100";
            when 1880 => rom_word <= "11001100";
            when 1881 => rom_word <= "11001100";
            when 1882 => rom_word <= "11001100";
            when 1883 => rom_word <= "01111000";
            when 1893 => rom_word <= "10001101";
            when 1894 => rom_word <= "10001101";
            when 1895 => rom_word <= "10001101";
            when 1896 => rom_word <= "10001101";
            when 1897 => rom_word <= "10001101";
            when 1898 => rom_word <= "11011000";
            when 1899 => rom_word <= "00100000";
            when 1909 => rom_word <= "10001101";
            when 1910 => rom_word <= "10001101";
            when 1911 => rom_word <= "10101101";
            when 1912 => rom_word <= "10101101";
            when 1913 => rom_word <= "10101101";
            when 1914 => rom_word <= "11111101";
            when 1915 => rom_word <= "11011000";
            when 1925 => rom_word <= "10001101";
            when 1926 => rom_word <= "11011000";
            when 1927 => rom_word <= "01110000";
            when 1928 => rom_word <= "01110000";
            when 1929 => rom_word <= "01110000";
            when 1930 => rom_word <= "11011000";
            when 1931 => rom_word <= "10001101";
            when 1941 => rom_word <= "10001101";
            when 1942 => rom_word <= "10001101";
            when 1943 => rom_word <= "10001101";
            when 1944 => rom_word <= "10001101";
            when 1945 => rom_word <= "10001101";
            when 1946 => rom_word <= "11001101";
            when 1947 => rom_word <= "10111001";
            when 1948 => rom_word <= "10000001";
            when 1949 => rom_word <= "11000100";
            when 1950 => rom_word <= "01111000";
            when 1957 => rom_word <= "11111101";
            when 1958 => rom_word <= "11000000";
            when 1959 => rom_word <= "01100000";
            when 1960 => rom_word <= "00110000";
            when 1961 => rom_word <= "00011000";
            when 1962 => rom_word <= "00001100";
            when 1963 => rom_word <= "11111101";
            when 1970 => rom_word <= "11000001";
            when 1971 => rom_word <= "01100000";
            when 1972 => rom_word <= "01100000";
            when 1973 => rom_word <= "01100000";
            when 1974 => rom_word <= "00111000";
            when 1975 => rom_word <= "01100000";
            when 1976 => rom_word <= "01100000";
            when 1977 => rom_word <= "01100000";
            when 1978 => rom_word <= "01100000";
            when 1979 => rom_word <= "11000001";
            when 1986 => rom_word <= "01100000";
            when 1987 => rom_word <= "01100000";
            when 1988 => rom_word <= "01100000";
            when 1989 => rom_word <= "01100000";
            when 1990 => rom_word <= "01100000";
            when 1991 => rom_word <= "01100000";
            when 1992 => rom_word <= "01100000";
            when 1993 => rom_word <= "01100000";
            when 1994 => rom_word <= "01100000";
            when 1995 => rom_word <= "01100000";
            when 2002 => rom_word <= "00111000";
            when 2003 => rom_word <= "01100000";
            when 2004 => rom_word <= "01100000";
            when 2005 => rom_word <= "01100000";
            when 2006 => rom_word <= "11000001";
            when 2007 => rom_word <= "01100000";
            when 2008 => rom_word <= "01100000";
            when 2009 => rom_word <= "01100000";
            when 2010 => rom_word <= "01100000";
            when 2011 => rom_word <= "00111000";
            when 2017 => rom_word <= "10111001";
            when 2018 => rom_word <= "11101100";
            when 2036 => rom_word <= "00100000";
            when 2037 => rom_word <= "01110000";
            when 2038 => rom_word <= "11011000";
            when 2039 => rom_word <= "10001101";
            when 2040 => rom_word <= "10001101";
            when 2041 => rom_word <= "10001101";
            when 2042 => rom_word <= "11111101";
            when 2051 => rom_word <= "11110000";
            when 2052 => rom_word <= "10011001";
            when 2053 => rom_word <= "00001100";
            when 2054 => rom_word <= "00001100";
            when 2055 => rom_word <= "00001100";
            when 2056 => rom_word <= "10001101";
            when 2057 => rom_word <= "10011001";
            when 2058 => rom_word <= "11110000";
            when 2059 => rom_word <= "01100000";
            when 2060 => rom_word <= "11001100";
            when 2061 => rom_word <= "01110000";
            when 2066 => rom_word <= "11001100";
            when 2067 => rom_word <= "11001100";
            when 2069 => rom_word <= "11001100";
            when 2070 => rom_word <= "11001100";
            when 2071 => rom_word <= "11001100";
            when 2072 => rom_word <= "11001100";
            when 2073 => rom_word <= "11001100";
            when 2074 => rom_word <= "11001100";
            when 2075 => rom_word <= "01111000";
            when 2081 => rom_word <= "11000000";
            when 2082 => rom_word <= "01100000";
            when 2083 => rom_word <= "00110000";
            when 2085 => rom_word <= "11111000";
            when 2086 => rom_word <= "10001101";
            when 2087 => rom_word <= "11111101";
            when 2088 => rom_word <= "00001100";
            when 2089 => rom_word <= "00001100";
            when 2090 => rom_word <= "00001101";
            when 2091 => rom_word <= "11111000";
            when 2097 => rom_word <= "00100000";
            when 2098 => rom_word <= "01110000";
            when 2099 => rom_word <= "11011000";
            when 2101 => rom_word <= "01111000";
            when 2102 => rom_word <= "11000000";
            when 2103 => rom_word <= "11111000";
            when 2104 => rom_word <= "11001100";
            when 2105 => rom_word <= "11001100";
            when 2106 => rom_word <= "11001100";
            when 2107 => rom_word <= "10111001";
            when 2114 => rom_word <= "11001100";
            when 2117 => rom_word <= "01111000";
            when 2118 => rom_word <= "11000000";
            when 2119 => rom_word <= "11111000";
            when 2120 => rom_word <= "11001100";
            when 2121 => rom_word <= "11001100";
            when 2122 => rom_word <= "11001100";
            when 2123 => rom_word <= "10111001";
            when 2129 => rom_word <= "00011000";
            when 2130 => rom_word <= "00110000";
            when 2131 => rom_word <= "01100000";
            when 2133 => rom_word <= "01111000";
            when 2134 => rom_word <= "11000000";
            when 2135 => rom_word <= "11111000";
            when 2136 => rom_word <= "11001100";
            when 2137 => rom_word <= "11001100";
            when 2138 => rom_word <= "11001100";
            when 2139 => rom_word <= "10111001";
            when 2145 => rom_word <= "01110000";
            when 2146 => rom_word <= "11011000";
            when 2147 => rom_word <= "01110000";
            when 2149 => rom_word <= "01111000";
            when 2150 => rom_word <= "11000000";
            when 2151 => rom_word <= "11111000";
            when 2152 => rom_word <= "11001100";
            when 2153 => rom_word <= "11001100";
            when 2154 => rom_word <= "11001100";
            when 2155 => rom_word <= "10111001";
            when 2165 => rom_word <= "11111000";
            when 2166 => rom_word <= "10001101";
            when 2167 => rom_word <= "00001100";
            when 2168 => rom_word <= "00001100";
            when 2169 => rom_word <= "00001100";
            when 2170 => rom_word <= "10001101";
            when 2171 => rom_word <= "11111000";
            when 2172 => rom_word <= "01100000";
            when 2173 => rom_word <= "00111000";
            when 2177 => rom_word <= "00100000";
            when 2178 => rom_word <= "01110000";
            when 2179 => rom_word <= "11011000";
            when 2181 => rom_word <= "11111000";
            when 2182 => rom_word <= "10001101";
            when 2183 => rom_word <= "11111101";
            when 2184 => rom_word <= "00001100";
            when 2185 => rom_word <= "00001100";
            when 2186 => rom_word <= "00001101";
            when 2187 => rom_word <= "11111000";
            when 2194 => rom_word <= "10001101";
            when 2197 => rom_word <= "11111000";
            when 2198 => rom_word <= "10001101";
            when 2199 => rom_word <= "11111101";
            when 2200 => rom_word <= "00001100";
            when 2201 => rom_word <= "00001100";
            when 2202 => rom_word <= "00001101";
            when 2203 => rom_word <= "11111000";
            when 2209 => rom_word <= "00011000";
            when 2210 => rom_word <= "00110000";
            when 2211 => rom_word <= "01100000";
            when 2213 => rom_word <= "11111000";
            when 2214 => rom_word <= "10001101";
            when 2215 => rom_word <= "11111101";
            when 2216 => rom_word <= "00001100";
            when 2217 => rom_word <= "00001100";
            when 2218 => rom_word <= "00001101";
            when 2219 => rom_word <= "11111000";
            when 2226 => rom_word <= "10011001";
            when 2229 => rom_word <= "01110000";
            when 2230 => rom_word <= "01100000";
            when 2231 => rom_word <= "01100000";
            when 2232 => rom_word <= "01100000";
            when 2233 => rom_word <= "01100000";
            when 2234 => rom_word <= "01100000";
            when 2235 => rom_word <= "01100000";
            when 2241 => rom_word <= "01100000";
            when 2242 => rom_word <= "11110000";
            when 2243 => rom_word <= "10011001";
            when 2245 => rom_word <= "01110000";
            when 2246 => rom_word <= "01100000";
            when 2247 => rom_word <= "01100000";
            when 2248 => rom_word <= "01100000";
            when 2249 => rom_word <= "01100000";
            when 2250 => rom_word <= "01100000";
            when 2251 => rom_word <= "01100000";
            when 2257 => rom_word <= "00011000";
            when 2258 => rom_word <= "00110000";
            when 2259 => rom_word <= "01100000";
            when 2261 => rom_word <= "01110000";
            when 2262 => rom_word <= "01100000";
            when 2263 => rom_word <= "01100000";
            when 2264 => rom_word <= "01100000";
            when 2265 => rom_word <= "01100000";
            when 2266 => rom_word <= "01100000";
            when 2267 => rom_word <= "01100000";
            when 2273 => rom_word <= "10001101";
            when 2275 => rom_word <= "00100000";
            when 2276 => rom_word <= "01110000";
            when 2277 => rom_word <= "11011000";
            when 2278 => rom_word <= "10001101";
            when 2279 => rom_word <= "10001101";
            when 2280 => rom_word <= "11111101";
            when 2281 => rom_word <= "10001101";
            when 2282 => rom_word <= "10001101";
            when 2283 => rom_word <= "10001101";
            when 2288 => rom_word <= "01110000";
            when 2289 => rom_word <= "11011000";
            when 2290 => rom_word <= "01110000";
            when 2291 => rom_word <= "00100000";
            when 2292 => rom_word <= "01110000";
            when 2293 => rom_word <= "11011000";
            when 2294 => rom_word <= "10001101";
            when 2295 => rom_word <= "11111101";
            when 2296 => rom_word <= "10001101";
            when 2297 => rom_word <= "10001101";
            when 2298 => rom_word <= "10001101";
            when 2299 => rom_word <= "10001101";
            when 2304 => rom_word <= "01100000";
            when 2305 => rom_word <= "00110000";
            when 2307 => rom_word <= "11111100";
            when 2308 => rom_word <= "00001100";
            when 2309 => rom_word <= "00001100";
            when 2310 => rom_word <= "00001100";
            when 2311 => rom_word <= "00111100";
            when 2312 => rom_word <= "00001100";
            when 2313 => rom_word <= "00001100";
            when 2314 => rom_word <= "00001100";
            when 2315 => rom_word <= "11111100";
            when 2325 => rom_word <= "11011100";
            when 2326 => rom_word <= "10110001";
            when 2327 => rom_word <= "10110001";
            when 2328 => rom_word <= "11111001";
            when 2329 => rom_word <= "01101100";
            when 2330 => rom_word <= "01101100";
            when 2331 => rom_word <= "11011001";
            when 2338 => rom_word <= "11110001";
            when 2339 => rom_word <= "11011000";
            when 2340 => rom_word <= "11001100";
            when 2341 => rom_word <= "11001100";
            when 2342 => rom_word <= "11111101";
            when 2343 => rom_word <= "11001100";
            when 2344 => rom_word <= "11001100";
            when 2345 => rom_word <= "11001100";
            when 2346 => rom_word <= "11001100";
            when 2347 => rom_word <= "11001101";
            when 2353 => rom_word <= "00100000";
            when 2354 => rom_word <= "01110000";
            when 2355 => rom_word <= "11011000";
            when 2357 => rom_word <= "11111000";
            when 2358 => rom_word <= "10001101";
            when 2359 => rom_word <= "10001101";
            when 2360 => rom_word <= "10001101";
            when 2361 => rom_word <= "10001101";
            when 2362 => rom_word <= "10001101";
            when 2363 => rom_word <= "11111000";
            when 2370 => rom_word <= "10001101";
            when 2373 => rom_word <= "11111000";
            when 2374 => rom_word <= "10001101";
            when 2375 => rom_word <= "10001101";
            when 2376 => rom_word <= "10001101";
            when 2377 => rom_word <= "10001101";
            when 2378 => rom_word <= "10001101";
            when 2379 => rom_word <= "11111000";
            when 2385 => rom_word <= "00011000";
            when 2386 => rom_word <= "00110000";
            when 2387 => rom_word <= "01100000";
            when 2389 => rom_word <= "11111000";
            when 2390 => rom_word <= "10001101";
            when 2391 => rom_word <= "10001101";
            when 2392 => rom_word <= "10001101";
            when 2393 => rom_word <= "10001101";
            when 2394 => rom_word <= "10001101";
            when 2395 => rom_word <= "11111000";
            when 2401 => rom_word <= "00110000";
            when 2402 => rom_word <= "01111000";
            when 2403 => rom_word <= "11001100";
            when 2405 => rom_word <= "11001100";
            when 2406 => rom_word <= "11001100";
            when 2407 => rom_word <= "11001100";
            when 2408 => rom_word <= "11001100";
            when 2409 => rom_word <= "11001100";
            when 2410 => rom_word <= "11001100";
            when 2411 => rom_word <= "01111000";
            when 2417 => rom_word <= "00011000";
            when 2418 => rom_word <= "00110000";
            when 2419 => rom_word <= "01100000";
            when 2421 => rom_word <= "11001100";
            when 2422 => rom_word <= "11001100";
            when 2423 => rom_word <= "11001100";
            when 2424 => rom_word <= "11001100";
            when 2425 => rom_word <= "11001100";
            when 2426 => rom_word <= "11001100";
            when 2427 => rom_word <= "01111000";
            when 2434 => rom_word <= "10001101";
            when 2437 => rom_word <= "10001101";
            when 2438 => rom_word <= "10001101";
            when 2439 => rom_word <= "10001101";
            when 2440 => rom_word <= "10001101";
            when 2441 => rom_word <= "10001101";
            when 2442 => rom_word <= "11001101";
            when 2443 => rom_word <= "10111001";
            when 2444 => rom_word <= "10000001";
            when 2445 => rom_word <= "11000100";
            when 2446 => rom_word <= "01111000";
            when 2449 => rom_word <= "10001101";
            when 2451 => rom_word <= "11111000";
            when 2452 => rom_word <= "10001101";
            when 2453 => rom_word <= "10001101";
            when 2454 => rom_word <= "10001101";
            when 2455 => rom_word <= "10001101";
            when 2456 => rom_word <= "10001101";
            when 2457 => rom_word <= "10001101";
            when 2458 => rom_word <= "10001101";
            when 2459 => rom_word <= "11111000";
            when 2465 => rom_word <= "10001101";
            when 2467 => rom_word <= "10001101";
            when 2468 => rom_word <= "10001101";
            when 2469 => rom_word <= "10001101";
            when 2470 => rom_word <= "10001101";
            when 2471 => rom_word <= "10001101";
            when 2472 => rom_word <= "10001101";
            when 2473 => rom_word <= "10001101";
            when 2474 => rom_word <= "10001101";
            when 2475 => rom_word <= "11111000";
            when 2481 => rom_word <= "01100000";
            when 2482 => rom_word <= "01100000";
            when 2483 => rom_word <= "11111000";
            when 2484 => rom_word <= "10001101";
            when 2485 => rom_word <= "00001100";
            when 2486 => rom_word <= "00001100";
            when 2487 => rom_word <= "00001100";
            when 2488 => rom_word <= "10001101";
            when 2489 => rom_word <= "11111000";
            when 2490 => rom_word <= "01100000";
            when 2491 => rom_word <= "01100000";
            when 2497 => rom_word <= "11110000";
            when 2498 => rom_word <= "00001001";
            when 2499 => rom_word <= "01100110";
            when 2500 => rom_word <= "10010110";
            when 2501 => rom_word <= "10010110";
            when 2502 => rom_word <= "00010110";
            when 2503 => rom_word <= "00010110";
            when 2504 => rom_word <= "10010110";
            when 2505 => rom_word <= "10010110";
            when 2506 => rom_word <= "01110110";
            when 2507 => rom_word <= "00001001";
            when 2508 => rom_word <= "11110000";
            when 2513 => rom_word <= "11110000";
            when 2514 => rom_word <= "00001001";
            when 2515 => rom_word <= "01110110";
            when 2516 => rom_word <= "10010110";
            when 2517 => rom_word <= "10010110";
            when 2518 => rom_word <= "01110110";
            when 2519 => rom_word <= "00110110";
            when 2520 => rom_word <= "01010110";
            when 2521 => rom_word <= "10010110";
            when 2522 => rom_word <= "10010110";
            when 2523 => rom_word <= "00001001";
            when 2524 => rom_word <= "11110000";
            when 2529 => rom_word <= "01111100";
            when 2530 => rom_word <= "11001100";
            when 2531 => rom_word <= "11001100";
            when 2532 => rom_word <= "01111100";
            when 2533 => rom_word <= "10001100";
            when 2534 => rom_word <= "11001100";
            when 2535 => rom_word <= "11101101";
            when 2536 => rom_word <= "11001100";
            when 2537 => rom_word <= "11001100";
            when 2538 => rom_word <= "11001100";
            when 2539 => rom_word <= "10001101";
            when 2545 => rom_word <= "11000001";
            when 2546 => rom_word <= "01100011";
            when 2547 => rom_word <= "01100000";
            when 2548 => rom_word <= "01100000";
            when 2549 => rom_word <= "01100000";
            when 2550 => rom_word <= "11111001";
            when 2551 => rom_word <= "01100000";
            when 2552 => rom_word <= "01100000";
            when 2553 => rom_word <= "01100000";
            when 2554 => rom_word <= "01101100";
            when 2555 => rom_word <= "00111000";
            when 2561 => rom_word <= "01100000";
            when 2562 => rom_word <= "00110000";
            when 2563 => rom_word <= "00011000";
            when 2565 => rom_word <= "01111000";
            when 2566 => rom_word <= "11000000";
            when 2567 => rom_word <= "11111000";
            when 2568 => rom_word <= "11001100";
            when 2569 => rom_word <= "11001100";
            when 2570 => rom_word <= "11001100";
            when 2571 => rom_word <= "10111001";
            when 2577 => rom_word <= "11000000";
            when 2578 => rom_word <= "01100000";
            when 2579 => rom_word <= "00110000";
            when 2581 => rom_word <= "01110000";
            when 2582 => rom_word <= "01100000";
            when 2583 => rom_word <= "01100000";
            when 2584 => rom_word <= "01100000";
            when 2585 => rom_word <= "01100000";
            when 2586 => rom_word <= "01100000";
            when 2587 => rom_word <= "01100000";
            when 2593 => rom_word <= "01100000";
            when 2594 => rom_word <= "00110000";
            when 2595 => rom_word <= "00011000";
            when 2597 => rom_word <= "11111000";
            when 2598 => rom_word <= "10001101";
            when 2599 => rom_word <= "10001101";
            when 2600 => rom_word <= "10001101";
            when 2601 => rom_word <= "10001101";
            when 2602 => rom_word <= "10001101";
            when 2603 => rom_word <= "11111000";
            when 2609 => rom_word <= "01100000";
            when 2610 => rom_word <= "00110000";
            when 2611 => rom_word <= "00011000";
            when 2613 => rom_word <= "11001100";
            when 2614 => rom_word <= "11001100";
            when 2615 => rom_word <= "11001100";
            when 2616 => rom_word <= "11001100";
            when 2617 => rom_word <= "11001100";
            when 2618 => rom_word <= "11001100";
            when 2619 => rom_word <= "01111000";
            when 2626 => rom_word <= "10111001";
            when 2627 => rom_word <= "11101100";
            when 2629 => rom_word <= "11101000";
            when 2630 => rom_word <= "10011001";
            when 2631 => rom_word <= "10011001";
            when 2632 => rom_word <= "10011001";
            when 2633 => rom_word <= "10011001";
            when 2634 => rom_word <= "10011001";
            when 2635 => rom_word <= "10011001";
            when 2640 => rom_word <= "10111001";
            when 2641 => rom_word <= "11101100";
            when 2643 => rom_word <= "10001101";
            when 2644 => rom_word <= "10011101";
            when 2645 => rom_word <= "10111101";
            when 2646 => rom_word <= "11111101";
            when 2647 => rom_word <= "11101101";
            when 2648 => rom_word <= "11001101";
            when 2649 => rom_word <= "10001101";
            when 2650 => rom_word <= "10001101";
            when 2651 => rom_word <= "10001101";
            when 2658 => rom_word <= "11110000";
            when 2659 => rom_word <= "11011000";
            when 2660 => rom_word <= "11011000";
            when 2661 => rom_word <= "11110001";
            when 2663 => rom_word <= "11111001";
            when 2674 => rom_word <= "01110000";
            when 2675 => rom_word <= "11011000";
            when 2676 => rom_word <= "11011000";
            when 2677 => rom_word <= "01110000";
            when 2679 => rom_word <= "11111000";
            when 2690 => rom_word <= "00110000";
            when 2691 => rom_word <= "00110000";
            when 2693 => rom_word <= "00110000";
            when 2694 => rom_word <= "00110000";
            when 2695 => rom_word <= "00011000";
            when 2696 => rom_word <= "00001100";
            when 2697 => rom_word <= "10001101";
            when 2698 => rom_word <= "10001101";
            when 2699 => rom_word <= "11111000";
            when 2710 => rom_word <= "11111101";
            when 2711 => rom_word <= "00001100";
            when 2712 => rom_word <= "00001100";
            when 2713 => rom_word <= "00001100";
            when 2714 => rom_word <= "00001100";
            when 2726 => rom_word <= "11111101";
            when 2727 => rom_word <= "10000001";
            when 2728 => rom_word <= "10000001";
            when 2729 => rom_word <= "10000001";
            when 2730 => rom_word <= "10000001";
            when 2737 => rom_word <= "00011000";
            when 2738 => rom_word <= "00011100";
            when 2739 => rom_word <= "00011001";
            when 2740 => rom_word <= "10011001";
            when 2741 => rom_word <= "11011000";
            when 2742 => rom_word <= "01100000";
            when 2743 => rom_word <= "00110000";
            when 2744 => rom_word <= "00011000";
            when 2745 => rom_word <= "11101100";
            when 2746 => rom_word <= "10000101";
            when 2747 => rom_word <= "11000000";
            when 2748 => rom_word <= "01100000";
            when 2749 => rom_word <= "11110001";
            when 2753 => rom_word <= "00011000";
            when 2754 => rom_word <= "00011100";
            when 2755 => rom_word <= "00011001";
            when 2756 => rom_word <= "10011001";
            when 2757 => rom_word <= "11011000";
            when 2758 => rom_word <= "01100000";
            when 2759 => rom_word <= "00110000";
            when 2760 => rom_word <= "10011001";
            when 2761 => rom_word <= "11001101";
            when 2762 => rom_word <= "01100101";
            when 2763 => rom_word <= "11110011";
            when 2764 => rom_word <= "10000001";
            when 2765 => rom_word <= "10000001";
            when 2770 => rom_word <= "01100000";
            when 2771 => rom_word <= "01100000";
            when 2773 => rom_word <= "01100000";
            when 2774 => rom_word <= "01100000";
            when 2775 => rom_word <= "01100000";
            when 2776 => rom_word <= "11110000";
            when 2777 => rom_word <= "11110000";
            when 2778 => rom_word <= "11110000";
            when 2779 => rom_word <= "01100000";
            when 2789 => rom_word <= "10110001";
            when 2790 => rom_word <= "11011000";
            when 2791 => rom_word <= "01101100";
            when 2792 => rom_word <= "11011000";
            when 2793 => rom_word <= "10110001";
            when 2805 => rom_word <= "01101100";
            when 2806 => rom_word <= "11011000";
            when 2807 => rom_word <= "10110001";
            when 2808 => rom_word <= "11011000";
            when 2809 => rom_word <= "01101100";
            when 2816 => rom_word <= "00100010";
            when 2817 => rom_word <= "10001000";
            when 2818 => rom_word <= "00100010";
            when 2819 => rom_word <= "10001000";
            when 2820 => rom_word <= "00100010";
            when 2821 => rom_word <= "10001000";
            when 2822 => rom_word <= "00100010";
            when 2823 => rom_word <= "10001000";
            when 2824 => rom_word <= "00100010";
            when 2825 => rom_word <= "10001000";
            when 2826 => rom_word <= "00100010";
            when 2827 => rom_word <= "10001000";
            when 2828 => rom_word <= "00100010";
            when 2829 => rom_word <= "10001000";
            when 2830 => rom_word <= "00100010";
            when 2831 => rom_word <= "10001000";
            when 2832 => rom_word <= "10101010";
            when 2833 => rom_word <= "01010101";
            when 2834 => rom_word <= "10101010";
            when 2835 => rom_word <= "01010101";
            when 2836 => rom_word <= "10101010";
            when 2837 => rom_word <= "01010101";
            when 2838 => rom_word <= "10101010";
            when 2839 => rom_word <= "01010101";
            when 2840 => rom_word <= "10101010";
            when 2841 => rom_word <= "01010101";
            when 2842 => rom_word <= "10101010";
            when 2843 => rom_word <= "01010101";
            when 2844 => rom_word <= "10101010";
            when 2845 => rom_word <= "01010101";
            when 2846 => rom_word <= "10101010";
            when 2847 => rom_word <= "01010101";
            when 2848 => rom_word <= "11101110";
            when 2849 => rom_word <= "10111011";
            when 2850 => rom_word <= "11101110";
            when 2851 => rom_word <= "10111011";
            when 2852 => rom_word <= "11101110";
            when 2853 => rom_word <= "10111011";
            when 2854 => rom_word <= "11101110";
            when 2855 => rom_word <= "10111011";
            when 2856 => rom_word <= "11101110";
            when 2857 => rom_word <= "10111011";
            when 2858 => rom_word <= "11101110";
            when 2859 => rom_word <= "10111011";
            when 2860 => rom_word <= "11101110";
            when 2861 => rom_word <= "10111011";
            when 2862 => rom_word <= "11101110";
            when 2863 => rom_word <= "10111011";
            when 2864 => rom_word <= "01100000";
            when 2865 => rom_word <= "01100000";
            when 2866 => rom_word <= "01100000";
            when 2867 => rom_word <= "01100000";
            when 2868 => rom_word <= "01100000";
            when 2869 => rom_word <= "01100000";
            when 2870 => rom_word <= "01100000";
            when 2871 => rom_word <= "01100000";
            when 2872 => rom_word <= "01100000";
            when 2873 => rom_word <= "01100000";
            when 2874 => rom_word <= "01100000";
            when 2875 => rom_word <= "01100000";
            when 2876 => rom_word <= "01100000";
            when 2877 => rom_word <= "01100000";
            when 2878 => rom_word <= "01100000";
            when 2879 => rom_word <= "01100000";
            when 2880 => rom_word <= "01100000";
            when 2881 => rom_word <= "01100000";
            when 2882 => rom_word <= "01100000";
            when 2883 => rom_word <= "01100000";
            when 2884 => rom_word <= "01100000";
            when 2885 => rom_word <= "01100000";
            when 2886 => rom_word <= "01100000";
            when 2887 => rom_word <= "01111100";
            when 2888 => rom_word <= "01100000";
            when 2889 => rom_word <= "01100000";
            when 2890 => rom_word <= "01100000";
            when 2891 => rom_word <= "01100000";
            when 2892 => rom_word <= "01100000";
            when 2893 => rom_word <= "01100000";
            when 2894 => rom_word <= "01100000";
            when 2895 => rom_word <= "01100000";
            when 2896 => rom_word <= "01100000";
            when 2897 => rom_word <= "01100000";
            when 2898 => rom_word <= "01100000";
            when 2899 => rom_word <= "01100000";
            when 2900 => rom_word <= "01100000";
            when 2901 => rom_word <= "01111100";
            when 2902 => rom_word <= "01100000";
            when 2903 => rom_word <= "01111100";
            when 2904 => rom_word <= "01100000";
            when 2905 => rom_word <= "01100000";
            when 2906 => rom_word <= "01100000";
            when 2907 => rom_word <= "01100000";
            when 2908 => rom_word <= "01100000";
            when 2909 => rom_word <= "01100000";
            when 2910 => rom_word <= "01100000";
            when 2911 => rom_word <= "01100000";
            when 2912 => rom_word <= "10110001";
            when 2913 => rom_word <= "10110001";
            when 2914 => rom_word <= "10110001";
            when 2915 => rom_word <= "10110001";
            when 2916 => rom_word <= "10110001";
            when 2917 => rom_word <= "10110001";
            when 2918 => rom_word <= "10110001";
            when 2919 => rom_word <= "10111101";
            when 2920 => rom_word <= "10110001";
            when 2921 => rom_word <= "10110001";
            when 2922 => rom_word <= "10110001";
            when 2923 => rom_word <= "10110001";
            when 2924 => rom_word <= "10110001";
            when 2925 => rom_word <= "10110001";
            when 2926 => rom_word <= "10110001";
            when 2927 => rom_word <= "10110001";
            when 2935 => rom_word <= "11111101";
            when 2936 => rom_word <= "10110001";
            when 2937 => rom_word <= "10110001";
            when 2938 => rom_word <= "10110001";
            when 2939 => rom_word <= "10110001";
            when 2940 => rom_word <= "10110001";
            when 2941 => rom_word <= "10110001";
            when 2942 => rom_word <= "10110001";
            when 2943 => rom_word <= "10110001";
            when 2949 => rom_word <= "01111100";
            when 2950 => rom_word <= "01100000";
            when 2951 => rom_word <= "01111100";
            when 2952 => rom_word <= "01100000";
            when 2953 => rom_word <= "01100000";
            when 2954 => rom_word <= "01100000";
            when 2955 => rom_word <= "01100000";
            when 2956 => rom_word <= "01100000";
            when 2957 => rom_word <= "01100000";
            when 2958 => rom_word <= "01100000";
            when 2959 => rom_word <= "01100000";
            when 2960 => rom_word <= "10110001";
            when 2961 => rom_word <= "10110001";
            when 2962 => rom_word <= "10110001";
            when 2963 => rom_word <= "10110001";
            when 2964 => rom_word <= "10110001";
            when 2965 => rom_word <= "10111101";
            when 2966 => rom_word <= "10000001";
            when 2967 => rom_word <= "10111101";
            when 2968 => rom_word <= "10110001";
            when 2969 => rom_word <= "10110001";
            when 2970 => rom_word <= "10110001";
            when 2971 => rom_word <= "10110001";
            when 2972 => rom_word <= "10110001";
            when 2973 => rom_word <= "10110001";
            when 2974 => rom_word <= "10110001";
            when 2975 => rom_word <= "10110001";
            when 2976 => rom_word <= "10110001";
            when 2977 => rom_word <= "10110001";
            when 2978 => rom_word <= "10110001";
            when 2979 => rom_word <= "10110001";
            when 2980 => rom_word <= "10110001";
            when 2981 => rom_word <= "10110001";
            when 2982 => rom_word <= "10110001";
            when 2983 => rom_word <= "10110001";
            when 2984 => rom_word <= "10110001";
            when 2985 => rom_word <= "10110001";
            when 2986 => rom_word <= "10110001";
            when 2987 => rom_word <= "10110001";
            when 2988 => rom_word <= "10110001";
            when 2989 => rom_word <= "10110001";
            when 2990 => rom_word <= "10110001";
            when 2991 => rom_word <= "10110001";
            when 2997 => rom_word <= "11111101";
            when 2998 => rom_word <= "10000001";
            when 2999 => rom_word <= "10111101";
            when 3000 => rom_word <= "10110001";
            when 3001 => rom_word <= "10110001";
            when 3002 => rom_word <= "10110001";
            when 3003 => rom_word <= "10110001";
            when 3004 => rom_word <= "10110001";
            when 3005 => rom_word <= "10110001";
            when 3006 => rom_word <= "10110001";
            when 3007 => rom_word <= "10110001";
            when 3008 => rom_word <= "10110001";
            when 3009 => rom_word <= "10110001";
            when 3010 => rom_word <= "10110001";
            when 3011 => rom_word <= "10110001";
            when 3012 => rom_word <= "10110001";
            when 3013 => rom_word <= "10111101";
            when 3014 => rom_word <= "10000001";
            when 3015 => rom_word <= "11111101";
            when 3024 => rom_word <= "10110001";
            when 3025 => rom_word <= "10110001";
            when 3026 => rom_word <= "10110001";
            when 3027 => rom_word <= "10110001";
            when 3028 => rom_word <= "10110001";
            when 3029 => rom_word <= "10110001";
            when 3030 => rom_word <= "10110001";
            when 3031 => rom_word <= "11111101";
            when 3040 => rom_word <= "01100000";
            when 3041 => rom_word <= "01100000";
            when 3042 => rom_word <= "01100000";
            when 3043 => rom_word <= "01100000";
            when 3044 => rom_word <= "01100000";
            when 3045 => rom_word <= "01111100";
            when 3046 => rom_word <= "01100000";
            when 3047 => rom_word <= "01111100";
            when 3063 => rom_word <= "01111100";
            when 3064 => rom_word <= "01100000";
            when 3065 => rom_word <= "01100000";
            when 3066 => rom_word <= "01100000";
            when 3067 => rom_word <= "01100000";
            when 3068 => rom_word <= "01100000";
            when 3069 => rom_word <= "01100000";
            when 3070 => rom_word <= "01100000";
            when 3071 => rom_word <= "01100000";
            when 3072 => rom_word <= "01100000";
            when 3073 => rom_word <= "01100000";
            when 3074 => rom_word <= "01100000";
            when 3075 => rom_word <= "01100000";
            when 3076 => rom_word <= "01100000";
            when 3077 => rom_word <= "01100000";
            when 3078 => rom_word <= "01100000";
            when 3079 => rom_word <= "11100011";
            when 3088 => rom_word <= "01100000";
            when 3089 => rom_word <= "01100000";
            when 3090 => rom_word <= "01100000";
            when 3091 => rom_word <= "01100000";
            when 3092 => rom_word <= "01100000";
            when 3093 => rom_word <= "01100000";
            when 3094 => rom_word <= "01100000";
            when 3095 => rom_word <= "11111111";
            when 3111 => rom_word <= "11111111";
            when 3112 => rom_word <= "01100000";
            when 3113 => rom_word <= "01100000";
            when 3114 => rom_word <= "01100000";
            when 3115 => rom_word <= "01100000";
            when 3116 => rom_word <= "01100000";
            when 3117 => rom_word <= "01100000";
            when 3118 => rom_word <= "01100000";
            when 3119 => rom_word <= "01100000";
            when 3120 => rom_word <= "01100000";
            when 3121 => rom_word <= "01100000";
            when 3122 => rom_word <= "01100000";
            when 3123 => rom_word <= "01100000";
            when 3124 => rom_word <= "01100000";
            when 3125 => rom_word <= "01100000";
            when 3126 => rom_word <= "01100000";
            when 3127 => rom_word <= "11100011";
            when 3128 => rom_word <= "01100000";
            when 3129 => rom_word <= "01100000";
            when 3130 => rom_word <= "01100000";
            when 3131 => rom_word <= "01100000";
            when 3132 => rom_word <= "01100000";
            when 3133 => rom_word <= "01100000";
            when 3134 => rom_word <= "01100000";
            when 3135 => rom_word <= "01100000";
            when 3143 => rom_word <= "11111111";
            when 3152 => rom_word <= "01100000";
            when 3153 => rom_word <= "01100000";
            when 3154 => rom_word <= "01100000";
            when 3155 => rom_word <= "01100000";
            when 3156 => rom_word <= "01100000";
            when 3157 => rom_word <= "01100000";
            when 3158 => rom_word <= "01100000";
            when 3159 => rom_word <= "11111111";
            when 3160 => rom_word <= "01100000";
            when 3161 => rom_word <= "01100000";
            when 3162 => rom_word <= "01100000";
            when 3163 => rom_word <= "01100000";
            when 3164 => rom_word <= "01100000";
            when 3165 => rom_word <= "01100000";
            when 3166 => rom_word <= "01100000";
            when 3167 => rom_word <= "01100000";
            when 3168 => rom_word <= "01100000";
            when 3169 => rom_word <= "01100000";
            when 3170 => rom_word <= "01100000";
            when 3171 => rom_word <= "01100000";
            when 3172 => rom_word <= "01100000";
            when 3173 => rom_word <= "11100011";
            when 3174 => rom_word <= "01100000";
            when 3175 => rom_word <= "11100011";
            when 3176 => rom_word <= "01100000";
            when 3177 => rom_word <= "01100000";
            when 3178 => rom_word <= "01100000";
            when 3179 => rom_word <= "01100000";
            when 3180 => rom_word <= "01100000";
            when 3181 => rom_word <= "01100000";
            when 3182 => rom_word <= "01100000";
            when 3183 => rom_word <= "01100000";
            when 3184 => rom_word <= "10110001";
            when 3185 => rom_word <= "10110001";
            when 3186 => rom_word <= "10110001";
            when 3187 => rom_word <= "10110001";
            when 3188 => rom_word <= "10110001";
            when 3189 => rom_word <= "10110001";
            when 3190 => rom_word <= "10110001";
            when 3191 => rom_word <= "10110011";
            when 3192 => rom_word <= "10110001";
            when 3193 => rom_word <= "10110001";
            when 3194 => rom_word <= "10110001";
            when 3195 => rom_word <= "10110001";
            when 3196 => rom_word <= "10110001";
            when 3197 => rom_word <= "10110001";
            when 3198 => rom_word <= "10110001";
            when 3199 => rom_word <= "10110001";
            when 3200 => rom_word <= "10110001";
            when 3201 => rom_word <= "10110001";
            when 3202 => rom_word <= "10110001";
            when 3203 => rom_word <= "10110001";
            when 3204 => rom_word <= "10110001";
            when 3205 => rom_word <= "10110011";
            when 3206 => rom_word <= "00110000";
            when 3207 => rom_word <= "11110011";
            when 3221 => rom_word <= "11110011";
            when 3222 => rom_word <= "00110000";
            when 3223 => rom_word <= "10110011";
            when 3224 => rom_word <= "10110001";
            when 3225 => rom_word <= "10110001";
            when 3226 => rom_word <= "10110001";
            when 3227 => rom_word <= "10110001";
            when 3228 => rom_word <= "10110001";
            when 3229 => rom_word <= "10110001";
            when 3230 => rom_word <= "10110001";
            when 3231 => rom_word <= "10110001";
            when 3232 => rom_word <= "10110001";
            when 3233 => rom_word <= "10110001";
            when 3234 => rom_word <= "10110001";
            when 3235 => rom_word <= "10110001";
            when 3236 => rom_word <= "10110001";
            when 3237 => rom_word <= "10111111";
            when 3239 => rom_word <= "11111111";
            when 3253 => rom_word <= "11111111";
            when 3255 => rom_word <= "10111111";
            when 3256 => rom_word <= "10110001";
            when 3257 => rom_word <= "10110001";
            when 3258 => rom_word <= "10110001";
            when 3259 => rom_word <= "10110001";
            when 3260 => rom_word <= "10110001";
            when 3261 => rom_word <= "10110001";
            when 3262 => rom_word <= "10110001";
            when 3263 => rom_word <= "10110001";
            when 3264 => rom_word <= "10110001";
            when 3265 => rom_word <= "10110001";
            when 3266 => rom_word <= "10110001";
            when 3267 => rom_word <= "10110001";
            when 3268 => rom_word <= "10110001";
            when 3269 => rom_word <= "10110011";
            when 3270 => rom_word <= "00110000";
            when 3271 => rom_word <= "10110011";
            when 3272 => rom_word <= "10110001";
            when 3273 => rom_word <= "10110001";
            when 3274 => rom_word <= "10110001";
            when 3275 => rom_word <= "10110001";
            when 3276 => rom_word <= "10110001";
            when 3277 => rom_word <= "10110001";
            when 3278 => rom_word <= "10110001";
            when 3279 => rom_word <= "10110001";
            when 3285 => rom_word <= "11111111";
            when 3287 => rom_word <= "11111111";
            when 3296 => rom_word <= "10110001";
            when 3297 => rom_word <= "10110001";
            when 3298 => rom_word <= "10110001";
            when 3299 => rom_word <= "10110001";
            when 3300 => rom_word <= "10110001";
            when 3301 => rom_word <= "10111111";
            when 3303 => rom_word <= "10111111";
            when 3304 => rom_word <= "10110001";
            when 3305 => rom_word <= "10110001";
            when 3306 => rom_word <= "10110001";
            when 3307 => rom_word <= "10110001";
            when 3308 => rom_word <= "10110001";
            when 3309 => rom_word <= "10110001";
            when 3310 => rom_word <= "10110001";
            when 3311 => rom_word <= "10110001";
            when 3312 => rom_word <= "01100000";
            when 3313 => rom_word <= "01100000";
            when 3314 => rom_word <= "01100000";
            when 3315 => rom_word <= "01100000";
            when 3316 => rom_word <= "01100000";
            when 3317 => rom_word <= "11111111";
            when 3319 => rom_word <= "11111111";
            when 3328 => rom_word <= "10110001";
            when 3329 => rom_word <= "10110001";
            when 3330 => rom_word <= "10110001";
            when 3331 => rom_word <= "10110001";
            when 3332 => rom_word <= "10110001";
            when 3333 => rom_word <= "10110001";
            when 3334 => rom_word <= "10110001";
            when 3335 => rom_word <= "11111111";
            when 3349 => rom_word <= "11111111";
            when 3351 => rom_word <= "11111111";
            when 3352 => rom_word <= "01100000";
            when 3353 => rom_word <= "01100000";
            when 3354 => rom_word <= "01100000";
            when 3355 => rom_word <= "01100000";
            when 3356 => rom_word <= "01100000";
            when 3357 => rom_word <= "01100000";
            when 3358 => rom_word <= "01100000";
            when 3359 => rom_word <= "01100000";
            when 3367 => rom_word <= "11111111";
            when 3368 => rom_word <= "10110001";
            when 3369 => rom_word <= "10110001";
            when 3370 => rom_word <= "10110001";
            when 3371 => rom_word <= "10110001";
            when 3372 => rom_word <= "10110001";
            when 3373 => rom_word <= "10110001";
            when 3374 => rom_word <= "10110001";
            when 3375 => rom_word <= "10110001";
            when 3376 => rom_word <= "10110001";
            when 3377 => rom_word <= "10110001";
            when 3378 => rom_word <= "10110001";
            when 3379 => rom_word <= "10110001";
            when 3380 => rom_word <= "10110001";
            when 3381 => rom_word <= "10110001";
            when 3382 => rom_word <= "10110001";
            when 3383 => rom_word <= "11110011";
            when 3392 => rom_word <= "01100000";
            when 3393 => rom_word <= "01100000";
            when 3394 => rom_word <= "01100000";
            when 3395 => rom_word <= "01100000";
            when 3396 => rom_word <= "01100000";
            when 3397 => rom_word <= "11100011";
            when 3398 => rom_word <= "01100000";
            when 3399 => rom_word <= "11100011";
            when 3413 => rom_word <= "11100011";
            when 3414 => rom_word <= "01100000";
            when 3415 => rom_word <= "11100011";
            when 3416 => rom_word <= "01100000";
            when 3417 => rom_word <= "01100000";
            when 3418 => rom_word <= "01100000";
            when 3419 => rom_word <= "01100000";
            when 3420 => rom_word <= "01100000";
            when 3421 => rom_word <= "01100000";
            when 3422 => rom_word <= "01100000";
            when 3423 => rom_word <= "01100000";
            when 3431 => rom_word <= "11110011";
            when 3432 => rom_word <= "10110001";
            when 3433 => rom_word <= "10110001";
            when 3434 => rom_word <= "10110001";
            when 3435 => rom_word <= "10110001";
            when 3436 => rom_word <= "10110001";
            when 3437 => rom_word <= "10110001";
            when 3438 => rom_word <= "10110001";
            when 3439 => rom_word <= "10110001";
            when 3440 => rom_word <= "10110001";
            when 3441 => rom_word <= "10110001";
            when 3442 => rom_word <= "10110001";
            when 3443 => rom_word <= "10110001";
            when 3444 => rom_word <= "10110001";
            when 3445 => rom_word <= "10110001";
            when 3446 => rom_word <= "10110001";
            when 3447 => rom_word <= "11111111";
            when 3448 => rom_word <= "10110001";
            when 3449 => rom_word <= "10110001";
            when 3450 => rom_word <= "10110001";
            when 3451 => rom_word <= "10110001";
            when 3452 => rom_word <= "10110001";
            when 3453 => rom_word <= "10110001";
            when 3454 => rom_word <= "10110001";
            when 3455 => rom_word <= "10110001";
            when 3456 => rom_word <= "01100000";
            when 3457 => rom_word <= "01100000";
            when 3458 => rom_word <= "01100000";
            when 3459 => rom_word <= "01100000";
            when 3460 => rom_word <= "01100000";
            when 3461 => rom_word <= "11111111";
            when 3462 => rom_word <= "01100000";
            when 3463 => rom_word <= "11111111";
            when 3464 => rom_word <= "01100000";
            when 3465 => rom_word <= "01100000";
            when 3466 => rom_word <= "01100000";
            when 3467 => rom_word <= "01100000";
            when 3468 => rom_word <= "01100000";
            when 3469 => rom_word <= "01100000";
            when 3470 => rom_word <= "01100000";
            when 3471 => rom_word <= "01100000";
            when 3472 => rom_word <= "01100000";
            when 3473 => rom_word <= "01100000";
            when 3474 => rom_word <= "01100000";
            when 3475 => rom_word <= "01100000";
            when 3476 => rom_word <= "01100000";
            when 3477 => rom_word <= "01100000";
            when 3478 => rom_word <= "01100000";
            when 3479 => rom_word <= "01111100";
            when 3495 => rom_word <= "11100011";
            when 3496 => rom_word <= "01100000";
            when 3497 => rom_word <= "01100000";
            when 3498 => rom_word <= "01100000";
            when 3499 => rom_word <= "01100000";
            when 3500 => rom_word <= "01100000";
            when 3501 => rom_word <= "01100000";
            when 3502 => rom_word <= "01100000";
            when 3503 => rom_word <= "01100000";
            when 3504 => rom_word <= "11111111";
            when 3505 => rom_word <= "11111111";
            when 3506 => rom_word <= "11111111";
            when 3507 => rom_word <= "11111111";
            when 3508 => rom_word <= "11111111";
            when 3509 => rom_word <= "11111111";
            when 3510 => rom_word <= "11111111";
            when 3511 => rom_word <= "11111111";
            when 3512 => rom_word <= "11111111";
            when 3513 => rom_word <= "11111111";
            when 3514 => rom_word <= "11111111";
            when 3515 => rom_word <= "11111111";
            when 3516 => rom_word <= "11111111";
            when 3517 => rom_word <= "11111111";
            when 3518 => rom_word <= "11111111";
            when 3519 => rom_word <= "11111111";
            when 3527 => rom_word <= "11111111";
            when 3528 => rom_word <= "11111111";
            when 3529 => rom_word <= "11111111";
            when 3530 => rom_word <= "11111111";
            when 3531 => rom_word <= "11111111";
            when 3532 => rom_word <= "11111111";
            when 3533 => rom_word <= "11111111";
            when 3534 => rom_word <= "11111111";
            when 3535 => rom_word <= "11111111";
            when 3536 => rom_word <= "00111100";
            when 3537 => rom_word <= "00111100";
            when 3538 => rom_word <= "00111100";
            when 3539 => rom_word <= "00111100";
            when 3540 => rom_word <= "00111100";
            when 3541 => rom_word <= "00111100";
            when 3542 => rom_word <= "00111100";
            when 3543 => rom_word <= "00111100";
            when 3544 => rom_word <= "00111100";
            when 3545 => rom_word <= "00111100";
            when 3546 => rom_word <= "00111100";
            when 3547 => rom_word <= "00111100";
            when 3548 => rom_word <= "00111100";
            when 3549 => rom_word <= "00111100";
            when 3550 => rom_word <= "00111100";
            when 3551 => rom_word <= "00111100";
            when 3552 => rom_word <= "11000011";
            when 3553 => rom_word <= "11000011";
            when 3554 => rom_word <= "11000011";
            when 3555 => rom_word <= "11000011";
            when 3556 => rom_word <= "11000011";
            when 3557 => rom_word <= "11000011";
            when 3558 => rom_word <= "11000011";
            when 3559 => rom_word <= "11000011";
            when 3560 => rom_word <= "11000011";
            when 3561 => rom_word <= "11000011";
            when 3562 => rom_word <= "11000011";
            when 3563 => rom_word <= "11000011";
            when 3564 => rom_word <= "11000011";
            when 3565 => rom_word <= "11000011";
            when 3566 => rom_word <= "11000011";
            when 3567 => rom_word <= "11000011";
            when 3568 => rom_word <= "11111111";
            when 3569 => rom_word <= "11111111";
            when 3570 => rom_word <= "11111111";
            when 3571 => rom_word <= "11111111";
            when 3572 => rom_word <= "11111111";
            when 3573 => rom_word <= "11111111";
            when 3574 => rom_word <= "11111111";
            when 3589 => rom_word <= "10111001";
            when 3590 => rom_word <= "11101100";
            when 3591 => rom_word <= "01101100";
            when 3592 => rom_word <= "01101100";
            when 3593 => rom_word <= "01101100";
            when 3594 => rom_word <= "11101100";
            when 3595 => rom_word <= "10111001";
            when 3602 => rom_word <= "11111000";
            when 3603 => rom_word <= "11001101";
            when 3604 => rom_word <= "10001101";
            when 3605 => rom_word <= "11001101";
            when 3606 => rom_word <= "11101100";
            when 3607 => rom_word <= "01001100";
            when 3608 => rom_word <= "11001100";
            when 3609 => rom_word <= "11001100";
            when 3610 => rom_word <= "11001100";
            when 3611 => rom_word <= "01111100";
            when 3612 => rom_word <= "00001100";
            when 3613 => rom_word <= "00001100";
            when 3618 => rom_word <= "11111101";
            when 3619 => rom_word <= "10001101";
            when 3620 => rom_word <= "10001101";
            when 3621 => rom_word <= "00001100";
            when 3622 => rom_word <= "00001100";
            when 3623 => rom_word <= "00001100";
            when 3624 => rom_word <= "00001100";
            when 3625 => rom_word <= "00001100";
            when 3626 => rom_word <= "00001100";
            when 3627 => rom_word <= "00001100";
            when 3637 => rom_word <= "11111101";
            when 3638 => rom_word <= "11011000";
            when 3639 => rom_word <= "11011000";
            when 3640 => rom_word <= "11011000";
            when 3641 => rom_word <= "11011000";
            when 3642 => rom_word <= "11011000";
            when 3643 => rom_word <= "11011000";
            when 3650 => rom_word <= "11111101";
            when 3651 => rom_word <= "10001101";
            when 3652 => rom_word <= "00011000";
            when 3653 => rom_word <= "00110000";
            when 3654 => rom_word <= "01100000";
            when 3655 => rom_word <= "01100000";
            when 3656 => rom_word <= "00110000";
            when 3657 => rom_word <= "00011000";
            when 3658 => rom_word <= "10001101";
            when 3659 => rom_word <= "11111101";
            when 3669 => rom_word <= "11111001";
            when 3670 => rom_word <= "01101100";
            when 3671 => rom_word <= "01101100";
            when 3672 => rom_word <= "01101100";
            when 3673 => rom_word <= "01101100";
            when 3674 => rom_word <= "01101100";
            when 3675 => rom_word <= "00111000";
            when 3685 => rom_word <= "10011001";
            when 3686 => rom_word <= "10011001";
            when 3687 => rom_word <= "10011001";
            when 3688 => rom_word <= "10011001";
            when 3689 => rom_word <= "10011001";
            when 3690 => rom_word <= "10011001";
            when 3691 => rom_word <= "11111000";
            when 3692 => rom_word <= "00011000";
            when 3693 => rom_word <= "00011000";
            when 3694 => rom_word <= "00001100";
            when 3700 => rom_word <= "10111001";
            when 3701 => rom_word <= "11101100";
            when 3702 => rom_word <= "01100000";
            when 3703 => rom_word <= "01100000";
            when 3704 => rom_word <= "01100000";
            when 3705 => rom_word <= "01100000";
            when 3706 => rom_word <= "01100000";
            when 3707 => rom_word <= "01100000";
            when 3714 => rom_word <= "11111001";
            when 3715 => rom_word <= "01100000";
            when 3716 => rom_word <= "11110000";
            when 3717 => rom_word <= "10011001";
            when 3718 => rom_word <= "10011001";
            when 3719 => rom_word <= "10011001";
            when 3720 => rom_word <= "10011001";
            when 3721 => rom_word <= "11110000";
            when 3722 => rom_word <= "01100000";
            when 3723 => rom_word <= "11111001";
            when 3730 => rom_word <= "01110000";
            when 3731 => rom_word <= "11011000";
            when 3732 => rom_word <= "10001101";
            when 3733 => rom_word <= "10001101";
            when 3734 => rom_word <= "11111101";
            when 3735 => rom_word <= "10001101";
            when 3736 => rom_word <= "10001101";
            when 3737 => rom_word <= "10001101";
            when 3738 => rom_word <= "11011000";
            when 3739 => rom_word <= "01110000";
            when 3746 => rom_word <= "01110000";
            when 3747 => rom_word <= "11011000";
            when 3748 => rom_word <= "10001101";
            when 3749 => rom_word <= "10001101";
            when 3750 => rom_word <= "10001101";
            when 3751 => rom_word <= "11011000";
            when 3752 => rom_word <= "11011000";
            when 3753 => rom_word <= "11011000";
            when 3754 => rom_word <= "11011000";
            when 3755 => rom_word <= "11011101";
            when 3762 => rom_word <= "11100001";
            when 3763 => rom_word <= "00110000";
            when 3764 => rom_word <= "01100000";
            when 3765 => rom_word <= "11000000";
            when 3766 => rom_word <= "11110001";
            when 3767 => rom_word <= "10011001";
            when 3768 => rom_word <= "10011001";
            when 3769 => rom_word <= "10011001";
            when 3770 => rom_word <= "10011001";
            when 3771 => rom_word <= "11110000";
            when 3781 => rom_word <= "11111001";
            when 3782 => rom_word <= "01101111";
            when 3783 => rom_word <= "01101111";
            when 3784 => rom_word <= "01101111";
            when 3785 => rom_word <= "11111001";
            when 3795 => rom_word <= "00000011";
            when 3796 => rom_word <= "10000001";
            when 3797 => rom_word <= "11111001";
            when 3798 => rom_word <= "01101111";
            when 3799 => rom_word <= "01101111";
            when 3800 => rom_word <= "00111111";
            when 3801 => rom_word <= "11111001";
            when 3802 => rom_word <= "00011000";
            when 3803 => rom_word <= "00001100";
            when 3810 => rom_word <= "11100000";
            when 3811 => rom_word <= "00110000";
            when 3812 => rom_word <= "00011000";
            when 3813 => rom_word <= "00011000";
            when 3814 => rom_word <= "11111000";
            when 3815 => rom_word <= "00011000";
            when 3816 => rom_word <= "00011000";
            when 3817 => rom_word <= "00011000";
            when 3818 => rom_word <= "00110000";
            when 3819 => rom_word <= "11100000";
            when 3827 => rom_word <= "11111000";
            when 3828 => rom_word <= "10001101";
            when 3829 => rom_word <= "10001101";
            when 3830 => rom_word <= "10001101";
            when 3831 => rom_word <= "10001101";
            when 3832 => rom_word <= "10001101";
            when 3833 => rom_word <= "10001101";
            when 3834 => rom_word <= "10001101";
            when 3835 => rom_word <= "10001101";
            when 3844 => rom_word <= "11111101";
            when 3847 => rom_word <= "11111101";
            when 3850 => rom_word <= "11111101";
            when 3860 => rom_word <= "01100000";
            when 3861 => rom_word <= "01100000";
            when 3862 => rom_word <= "11111001";
            when 3863 => rom_word <= "01100000";
            when 3864 => rom_word <= "01100000";
            when 3867 => rom_word <= "11111001";
            when 3875 => rom_word <= "00110000";
            when 3876 => rom_word <= "01100000";
            when 3877 => rom_word <= "11000000";
            when 3878 => rom_word <= "10000001";
            when 3879 => rom_word <= "11000000";
            when 3880 => rom_word <= "01100000";
            when 3881 => rom_word <= "00110000";
            when 3883 => rom_word <= "11111001";
            when 3891 => rom_word <= "11000000";
            when 3892 => rom_word <= "01100000";
            when 3893 => rom_word <= "00110000";
            when 3894 => rom_word <= "00011000";
            when 3895 => rom_word <= "00110000";
            when 3896 => rom_word <= "01100000";
            when 3897 => rom_word <= "11000000";
            when 3899 => rom_word <= "11111001";
            when 3906 => rom_word <= "11000001";
            when 3907 => rom_word <= "01100011";
            when 3908 => rom_word <= "01100011";
            when 3909 => rom_word <= "01100000";
            when 3910 => rom_word <= "01100000";
            when 3911 => rom_word <= "01100000";
            when 3912 => rom_word <= "01100000";
            when 3913 => rom_word <= "01100000";
            when 3914 => rom_word <= "01100000";
            when 3915 => rom_word <= "01100000";
            when 3916 => rom_word <= "01100000";
            when 3917 => rom_word <= "01100000";
            when 3918 => rom_word <= "01100000";
            when 3919 => rom_word <= "01100000";
            when 3920 => rom_word <= "01100000";
            when 3921 => rom_word <= "01100000";
            when 3922 => rom_word <= "01100000";
            when 3923 => rom_word <= "01100000";
            when 3924 => rom_word <= "01100000";
            when 3925 => rom_word <= "01100000";
            when 3926 => rom_word <= "01100000";
            when 3927 => rom_word <= "01100000";
            when 3928 => rom_word <= "01100000";
            when 3929 => rom_word <= "01101100";
            when 3930 => rom_word <= "01101100";
            when 3931 => rom_word <= "01101100";
            when 3932 => rom_word <= "00111000";
            when 3941 => rom_word <= "01100000";
            when 3943 => rom_word <= "11111001";
            when 3945 => rom_word <= "01100000";
            when 3957 => rom_word <= "10111001";
            when 3958 => rom_word <= "11101100";
            when 3960 => rom_word <= "10111001";
            when 3961 => rom_word <= "11101100";
            when 3969 => rom_word <= "01110000";
            when 3970 => rom_word <= "11011000";
            when 3971 => rom_word <= "11011000";
            when 3972 => rom_word <= "01110000";
            when 3991 => rom_word <= "01100000";
            when 3992 => rom_word <= "01100000";
            when 4007 => rom_word <= "01100000";
            when 4017 => rom_word <= "11000011";
            when 4018 => rom_word <= "11000000";
            when 4019 => rom_word <= "11000000";
            when 4020 => rom_word <= "11000000";
            when 4021 => rom_word <= "11000000";
            when 4022 => rom_word <= "11000000";
            when 4023 => rom_word <= "11011100";
            when 4024 => rom_word <= "11011000";
            when 4025 => rom_word <= "11011000";
            when 4026 => rom_word <= "11110000";
            when 4027 => rom_word <= "11100000";
            when 4033 => rom_word <= "11011000";
            when 4034 => rom_word <= "10110001";
            when 4035 => rom_word <= "10110001";
            when 4036 => rom_word <= "10110001";
            when 4037 => rom_word <= "10110001";
            when 4038 => rom_word <= "10110001";
            when 4049 => rom_word <= "11110000";
            when 4050 => rom_word <= "10011001";
            when 4051 => rom_word <= "11000000";
            when 4052 => rom_word <= "01100000";
            when 4053 => rom_word <= "00110001";
            when 4054 => rom_word <= "11111001";
            when 4068 => rom_word <= "11111001";
            when 4069 => rom_word <= "11111001";
            when 4070 => rom_word <= "11111001";
            when 4071 => rom_word <= "11111001";
            when 4072 => rom_word <= "11111001";
            when 4073 => rom_word <= "11111001";
            when 4074 => rom_word <= "11111001";
            when others => rom_word <= X"00";
         end case;
      end if;
   end process;
end rtl;