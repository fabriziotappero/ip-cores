-- AC97_OC enable 
  constant CFG_AC97_OC  : integer := CONFIG_AC97_OC_ENABLE;

