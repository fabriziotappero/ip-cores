--Second Order Sections (SOS) automatically generated VHDL package file
--M.Eng. Alexander López Parrado


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package coefs_sos is 


--The number of sections
constant NSECT:integer:=6;

--Number of bits in fractional part of coeffcients
--Fixed point format with 16 bits ([3].[13])
constant Q: integer:=13;

--Gain on each stage
constant GAIN: std_logic_vector(15 downto 0):= std_logic_vector(to_signed(169,16));

--Filter Coefficients ...(b0,b1,b2,a0,a1,a2)_stage1,(b0,b1,b2,a0,a1,a2)_stage0
constant COEFFS: std_logic_vector(575 downto 0):="001000000000000011000000000000000010000000000000001000000000000011000011110101000001111110110000001000000000000011000000000111010001111111100011001000000000000011000100110001100001111110011101001000000000000010111111111000110010000000011101001000000000000011000100011001010001111100101000001000000000000000111111111011100001111111101110001000000000000011000101000110010001111100011001001000000000000001000000000000000010000000000000001000000000000011000101010011000001111010111110001000000000000001000000000100100010000000010010001000000000000011000101001000010001111010011100";

end coefs_sos;
