Paste synthesized model here