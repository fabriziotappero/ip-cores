000000 => x"cafe",
000001 => x"03f7",
000002 => x"929c",
000003 => x"426f",
000004 => x"6f74",
000005 => x"6c6f",
000006 => x"6164",
000007 => x"6572",
000008 => x"bc0e",
000009 => x"bc04",
000010 => x"bc03",
000011 => x"bc02",
000012 => x"bc01",
000013 => x"c000",
000014 => x"cc00",
000015 => x"ec8a",
000016 => x"cc19",
000017 => x"ed0f",
000018 => x"c520",
000019 => x"c907",
000020 => x"be73",
000021 => x"bc00",
000022 => x"ec11",
000023 => x"ec88",
000024 => x"ec8a",
000025 => x"c380",
000026 => x"cff8",
000027 => x"1c07",
000028 => x"2800",
000029 => x"ec08",
000030 => x"ec0b",
000031 => x"ec0d",
000032 => x"ec00",
000033 => x"ed88",
000034 => x"ed8b",
000035 => x"c064",
000036 => x"ed8d",
000037 => x"c901",
000038 => x"ed2f",
000039 => x"ec17",
000040 => x"ec97",
000041 => x"c160",
000042 => x"c909",
000043 => x"c18f",
000044 => x"0923",
000045 => x"29b3",
000046 => x"2a44",
000047 => x"100a",
000048 => x"149b",
000049 => x"9003",
000050 => x"0241",
000051 => x"bdfc",
000052 => x"ed49",
000053 => x"ec22",
000054 => x"d406",
000055 => x"ed0a",
000056 => x"c534",
000057 => x"c905",
000058 => x"be4d",
000059 => x"c12a",
000060 => x"c906",
000061 => x"be4a",
000062 => x"ee11",
000063 => x"be4c",
000064 => x"c13a",
000065 => x"c906",
000066 => x"be45",
000067 => x"ee97",
000068 => x"ee17",
000069 => x"be46",
000070 => x"0250",
000071 => x"be44",
000072 => x"be40",
000073 => x"ec27",
000074 => x"c083",
000075 => x"2001",
000076 => x"c330",
000077 => x"0b60",
000078 => x"bc0f",
000079 => x"c552",
000080 => x"c906",
000081 => x"be36",
000082 => x"c144",
000083 => x"c907",
000084 => x"be33",
000085 => x"c50a",
000086 => x"c907",
000087 => x"be30",
000088 => x"be32",
000089 => x"0300",
000090 => x"0080",
000091 => x"be2e",
000092 => x"be2c",
000093 => x"c0b0",
000094 => x"181e",
000095 => x"81f0",
000096 => x"c0b1",
000097 => x"181e",
000098 => x"8085",
000099 => x"c0b2",
000100 => x"181e",
000101 => x"8052",
000102 => x"c0b3",
000103 => x"181e",
000104 => x"8019",
000105 => x"c0b4",
000106 => x"181e",
000107 => x"8021",
000108 => x"c296",
000109 => x"ca83",
000110 => x"c0f0",
000111 => x"181e",
000112 => x"f705",
000113 => x"c0e4",
000114 => x"181e",
000115 => x"80e1",
000116 => x"c2c8",
000117 => x"ca85",
000118 => x"c0f7",
000119 => x"181e",
000120 => x"f705",
000121 => x"c0f2",
000122 => x"181e",
000123 => x"85da",
000124 => x"2800",
000125 => x"c080",
000126 => x"cc80",
000127 => x"ec99",
000128 => x"3400",
000129 => x"c14a",
000130 => x"c906",
000131 => x"be04",
000132 => x"2800",
000133 => x"2100",
000134 => x"bca0",
000135 => x"bc95",
000136 => x"bc95",
000137 => x"bc95",
000138 => x"bc95",
000139 => x"bc98",
000140 => x"c528",
000141 => x"c906",
000142 => x"be8e",
000143 => x"be96",
000144 => x"edca",
000145 => x"be94",
000146 => x"edc9",
000147 => x"c036",
000148 => x"c805",
000149 => x"3404",
000150 => x"be87",
000151 => x"be8d",
000152 => x"c47e",
000153 => x"cc4a",
000154 => x"180e",
000155 => x"8486",
000156 => x"be88",
000157 => x"3f64",
000158 => x"2066",
000159 => x"be85",
000160 => x"20e6",
000161 => x"be83",
000162 => x"2166",
000163 => x"be81",
000164 => x"21e6",
000165 => x"be7f",
000166 => x"2266",
000167 => x"be7d",
000168 => x"22e6",
000169 => x"be7b",
000170 => x"2366",
000171 => x"c280",
000172 => x"ecda",
000173 => x"ec5e",
000174 => x"be76",
000175 => x"7f5a",
000176 => x"ec06",
000177 => x"2806",
000178 => x"ec0e",
000179 => x"2400",
000180 => x"1858",
000181 => x"85f9",
000182 => x"bc53",
000183 => x"c100",
000184 => x"be28",
000185 => x"c47e",
000186 => x"cc4a",
000187 => x"180d",
000188 => x"8465",
000189 => x"c102",
000190 => x"be22",
000191 => x"2055",
000192 => x"c104",
000193 => x"be1f",
000194 => x"20d5",
000195 => x"c106",
000196 => x"be1c",
000197 => x"2155",
000198 => x"c108",
000199 => x"be19",
000200 => x"21d5",
000201 => x"c10a",
000202 => x"be16",
000203 => x"2255",
000204 => x"c10c",
000205 => x"be13",
000206 => x"22d5",
000207 => x"c10e",
000208 => x"be10",
000209 => x"2355",
000210 => x"c200",
000211 => x"ecca",
000212 => x"ec4e",
000213 => x"c010",
000214 => x"0940",
000215 => x"be09",
000216 => x"7eca",
000217 => x"ec06",
000218 => x"2805",
000219 => x"ec0e",
000220 => x"2400",
000221 => x"1848",
000222 => x"85f7",
000223 => x"bc2a",
000224 => x"0370",
000225 => x"be3f",
000226 => x"3eb0",
000227 => x"0121",
000228 => x"be3c",
000229 => x"26d3",
000230 => x"3460",
000231 => x"c162",
000232 => x"c906",
000233 => x"be33",
000234 => x"be2c",
000235 => x"c47e",
000236 => x"cc4a",
000237 => x"1818",
000238 => x"8433",
000239 => x"be27",
000240 => x"3c94",
000241 => x"2011",
000242 => x"be24",
000243 => x"2091",
000244 => x"be22",
000245 => x"2111",
000246 => x"be20",
000247 => x"2191",
000248 => x"be1e",
000249 => x"2211",
000250 => x"be1c",
000251 => x"2291",
000252 => x"be1a",
000253 => x"2311",
000254 => x"2ad5",
000255 => x"ecda",
000256 => x"ec5e",
000257 => x"be15",
000258 => x"7cda",
000259 => x"ec06",
000260 => x"2801",
000261 => x"ec0e",
000262 => x"2400",
000263 => x"1858",
000264 => x"85f9",
000265 => x"ec11",
000266 => x"ec8a",
000267 => x"c506",
000268 => x"c906",
000269 => x"be0f",
000270 => x"ec06",
000271 => x"2491",
000272 => x"1809",
000273 => x"8015",
000274 => x"c52e",
000275 => x"c907",
000276 => x"be08",
000277 => x"bccf",
000278 => x"0370",
000279 => x"be08",
000280 => x"3c80",
000281 => x"be06",
000282 => x"2490",
000283 => x"3460",
000284 => x"bccb",
000285 => x"bcd3",
000286 => x"bcd7",
000287 => x"bcdb",
000288 => x"bc71",
000289 => x"bcc0",
000290 => x"bd33",
000291 => x"bc6f",
000292 => x"bcc2",
000293 => x"bcda",
000294 => x"c176",
000295 => x"c906",
000296 => x"bebf",
000297 => x"24aa",
000298 => x"8010",
000299 => x"c0a2",
000300 => x"bec9",
000301 => x"24a2",
000302 => x"be20",
000303 => x"24b3",
000304 => x"be1e",
000305 => x"24c4",
000306 => x"be1c",
000307 => x"24d5",
000308 => x"be1a",
000309 => x"24e6",
000310 => x"be18",
000311 => x"c0a2",
000312 => x"bebd",
000313 => x"beb7",
000314 => x"c546",
000315 => x"c906",
000316 => x"beab",
000317 => x"ee06",
000318 => x"bee6",
000319 => x"beb1",
000320 => x"beb0",
000321 => x"beaf",
000322 => x"beae",
000323 => x"c080",
000324 => x"ccc0",
000325 => x"1c01",
000326 => x"2800",
000327 => x"ed0f",
000328 => x"ec88",
000329 => x"ec8b",
000330 => x"ec8c",
000331 => x"ec8a",
000332 => x"ec89",
000333 => x"3400",
000334 => x"0370",
000335 => x"3c90",
000336 => x"bea5",
000337 => x"3c90",
000338 => x"bea3",
000339 => x"3460",
000340 => x"c51a",
000341 => x"c906",
000342 => x"be91",
000343 => x"bea8",
000344 => x"c136",
000345 => x"c905",
000346 => x"3424",
000347 => x"ecca",
000348 => x"be94",
000349 => x"c280",
000350 => x"c00f",
000351 => x"2058",
000352 => x"840e",
000353 => x"be8f",
000354 => x"c0a4",
000355 => x"be92",
000356 => x"ee12",
000357 => x"bebf",
000358 => x"c0ae",
000359 => x"be8e",
000360 => x"0250",
000361 => x"bebb",
000362 => x"c0ba",
000363 => x"be8a",
000364 => x"c0a0",
000365 => x"be88",
000366 => x"7a5a",
000367 => x"c0a0",
000368 => x"be85",
000369 => x"beb3",
000370 => x"c00f",
000371 => x"2058",
000372 => x"8414",
000373 => x"c0a0",
000374 => x"be7f",
000375 => x"be7e",
000376 => x"c010",
000377 => x"1250",
000378 => x"c470",
000379 => x"2240",
000380 => x"c12e",
000381 => x"78c9",
000382 => x"3c90",
000383 => x"c880",
000384 => x"c020",
000385 => x"1818",
000386 => x"f8c2",
000387 => x"be72",
000388 => x"c08f",
000389 => x"2014",
000390 => x"3409",
000391 => x"85f6",
000392 => x"ec20",
000393 => x"dc0f",
000394 => x"b804",
000395 => x"c5fe",
000396 => x"343d",
000397 => x"85d1",
000398 => x"be6c",
000399 => x"2800",
000400 => x"3400",
000401 => x"bc54",
000402 => x"bc92",
000403 => x"c001",
000404 => x"ed0c",
000405 => x"c050",
000406 => x"c83f",
000407 => x"ed0a",
000408 => x"c000",
000409 => x"c801",
000410 => x"bea8",
000411 => x"c154",
000412 => x"c906",
000413 => x"be4a",
000414 => x"c162",
000415 => x"c906",
000416 => x"be47",
000417 => x"be59",
000418 => x"3c80",
000419 => x"be57",
000420 => x"2410",
000421 => x"c4fe",
000422 => x"ccca",
000423 => x"1809",
000424 => x"8439",
000425 => x"c100",
000426 => x"0290",
000427 => x"be2f",
000428 => x"be4e",
000429 => x"3c80",
000430 => x"be4c",
000431 => x"2690",
000432 => x"3ed4",
000433 => x"2055",
000434 => x"c102",
000435 => x"be27",
000436 => x"be46",
000437 => x"3c80",
000438 => x"be44",
000439 => x"2690",
000440 => x"20d5",
000441 => x"c104",
000442 => x"be20",
000443 => x"c106",
000444 => x"be3e",
000445 => x"0180",
000446 => x"be8a",
000447 => x"0121",
000448 => x"c010",
000449 => x"1828",
000450 => x"85fa",
000451 => x"2ad5",
000452 => x"be36",
000453 => x"0180",
000454 => x"be82",
000455 => x"0121",
000456 => x"2400",
000457 => x"02d1",
000458 => x"1858",
000459 => x"85f9",
000460 => x"c001",
000461 => x"ed0c",
000462 => x"c050",
000463 => x"c83f",
000464 => x"ed0a",
000465 => x"c00c",
000466 => x"c801",
000467 => x"be6f",
000468 => x"c506",
000469 => x"c906",
000470 => x"be11",
000471 => x"c68e",
000472 => x"ca80",
000473 => x"3450",
000474 => x"0370",
000475 => x"3dd0",
000476 => x"be6c",
000477 => x"0121",
000478 => x"01d0",
000479 => x"be69",
000480 => x"3460",
000481 => x"c512",
000482 => x"c907",
000483 => x"be04",
000484 => x"bcb9",
000485 => x"bc93",
000486 => x"bca4",
000487 => x"01f0",
000488 => x"78a9",
000489 => x"3c90",
000490 => x"c880",
000491 => x"3419",
000492 => x"8003",
000493 => x"be08",
000494 => x"bdfa",
000495 => x"3430",
000496 => x"0170",
000497 => x"c08d",
000498 => x"be03",
000499 => x"c08a",
000500 => x"03a0",
000501 => x"ec22",
000502 => x"dc05",
000503 => x"b9fe",
000504 => x"ed18",
000505 => x"3470",
000506 => x"ec20",
000507 => x"dc8f",
000508 => x"b9fe",
000509 => x"c800",
000510 => x"3470",
000511 => x"0170",
000512 => x"c200",
000513 => x"c184",
000514 => x"bff8",
000515 => x"c0c7",
000516 => x"1809",
000517 => x"9003",
000518 => x"c0a0",
000519 => x"1001",
000520 => x"c0b0",
000521 => x"1809",
000522 => x"91f8",
000523 => x"c0c6",
000524 => x"1818",
000525 => x"91f5",
000526 => x"c0b9",
000527 => x"1818",
000528 => x"a404",
000529 => x"c0c1",
000530 => x"1809",
000531 => x"a1ef",
000532 => x"0080",
000533 => x"bfe0",
000534 => x"c030",
000535 => x"1090",
000536 => x"c009",
000537 => x"1809",
000538 => x"a402",
000539 => x"0497",
000540 => x"3e42",
000541 => x"3e42",
000542 => x"3e42",
000543 => x"3e42",
000544 => x"2641",
000545 => x"05b9",
000546 => x"85e0",
000547 => x"3420",
000548 => x"0370",
000549 => x"3d42",
000550 => x"3d22",
000551 => x"3d22",
000552 => x"3d22",
000553 => x"be0f",
000554 => x"bfcb",
000555 => x"3d40",
000556 => x"be0c",
000557 => x"bfc8",
000558 => x"3d45",
000559 => x"3d25",
000560 => x"3d25",
000561 => x"3d25",
000562 => x"be06",
000563 => x"bfc2",
000564 => x"0140",
000565 => x"be03",
000566 => x"bfbf",
000567 => x"3460",
000568 => x"c08f",
000569 => x"2121",
000570 => x"c089",
000571 => x"181a",
000572 => x"8803",
000573 => x"c0b0",
000574 => x"bc02",
000575 => x"c0b7",
000576 => x"0892",
000577 => x"3470",
000578 => x"ed0b",
000579 => x"ec22",
000580 => x"dc03",
000581 => x"b9fe",
000582 => x"ec23",
000583 => x"3470",
000584 => x"00f0",
000585 => x"c050",
000586 => x"c837",
000587 => x"ed0a",
000588 => x"c001",
000589 => x"ed0c",
000590 => x"c006",
000591 => x"bff3",
000592 => x"c050",
000593 => x"c83f",
000594 => x"ed0a",
000595 => x"c000",
000596 => x"c805",
000597 => x"bfed",
000598 => x"dc01",
000599 => x"b805",
000600 => x"c53e",
000601 => x"c907",
000602 => x"bf8d",
000603 => x"bc42",
000604 => x"c040",
000605 => x"c83f",
000606 => x"ed0a",
000607 => x"c001",
000608 => x"ed0c",
000609 => x"3c20",
000610 => x"c802",
000611 => x"bfdf",
000612 => x"03a0",
000613 => x"cb80",
000614 => x"3ff0",
000615 => x"0030",
000616 => x"c800",
000617 => x"2407",
000618 => x"bfd8",
000619 => x"2800",
000620 => x"ed0c",
000621 => x"c050",
000622 => x"c83f",
000623 => x"ed0a",
000624 => x"c001",
000625 => x"ed0c",
000626 => x"c000",
000627 => x"c805",
000628 => x"bfce",
000629 => x"dc00",
000630 => x"b9fc",
000631 => x"3410",
000632 => x"00f0",
000633 => x"c040",
000634 => x"c83f",
000635 => x"ed0a",
000636 => x"c001",
000637 => x"ed0c",
000638 => x"3c20",
000639 => x"c803",
000640 => x"bfc2",
000641 => x"0020",
000642 => x"c800",
000643 => x"3c00",
000644 => x"bfbe",
000645 => x"29b3",
000646 => x"ed3c",
000647 => x"0180",
000648 => x"c980",
000649 => x"3410",
000650 => x"e5b0",
000651 => x"ec30",
000652 => x"dc06",
000653 => x"b9fe",
000654 => x"c306",
000655 => x"200e",
000656 => x"840a",
000657 => x"ecb1",
000658 => x"ef32",
000659 => x"2800",
000660 => x"009a",
000661 => x"0f60",
000662 => x"ed99",
000663 => x"edea",
000664 => x"ef34",
000665 => x"3470",
000666 => x"c550",
000667 => x"c907",
000668 => x"bf4b",
000669 => x"c55e",
000670 => x"c907",
000671 => x"bf48",
000672 => x"bf5a",
000673 => x"2800",
000674 => x"3400",
000675 => x"0170",
000676 => x"bf56",
000677 => x"c08d",
000678 => x"1809",
000679 => x"f702",
000680 => x"c088",
000681 => x"1809",
000682 => x"8034",
000683 => x"bdf9",
000684 => x"c528",
000685 => x"c906",
000686 => x"bf39",
000687 => x"bf50",
000688 => x"edca",
000689 => x"bf4e",
000690 => x"edc9",
000691 => x"bff0",
000692 => x"bf3c",
000693 => x"c536",
000694 => x"c906",
000695 => x"bf30",
000696 => x"bf47",
000697 => x"02c0",
000698 => x"bfe9",
000699 => x"bf35",
000700 => x"345d",
000701 => x"8021",
000702 => x"06d1",
000703 => x"bf31",
000704 => x"c0a4",
000705 => x"bf34",
000706 => x"ee32",
000707 => x"bf61",
000708 => x"ee31",
000709 => x"bf5f",
000710 => x"c0ba",
000711 => x"bf2e",
000712 => x"c0a0",
000713 => x"bf2c",
000714 => x"bfc0",
000715 => x"0260",
000716 => x"bf58",
000717 => x"c320",
000718 => x"c1ae",
000719 => x"00e0",
000720 => x"bf25",
000721 => x"3cc0",
000722 => x"c880",
000723 => x"181e",
000724 => x"f8c3",
000725 => x"bf20",
000726 => x"00c0",
000727 => x"c880",
000728 => x"181e",
000729 => x"f8c3",
000730 => x"bf1b",
000731 => x"eca0",
000732 => x"dc9f",
000733 => x"b9df",
000734 => x"bf12",
000735 => x"c69a",
000736 => x"ca80",
000737 => x"3450",
000738 => x"0d0a",
000739 => x"0d0a",
000740 => x"4174",
000741 => x"6c61",
000742 => x"732d",
000743 => x"324b",
000744 => x"2042",
000745 => x"6f6f",
000746 => x"746c",
000747 => x"6f61",
000748 => x"6465",
000749 => x"7220",
000750 => x"2d20",
000751 => x"5632",
000752 => x"3031",
000753 => x"3430",
000754 => x"3531",
000755 => x"360d",
000756 => x"0a62",
000757 => x"7920",
000758 => x"5374",
000759 => x"6570",
000760 => x"6861",
000761 => x"6e20",
000762 => x"4e6f",
000763 => x"6c74",
000764 => x"696e",
000765 => x"672c",
000766 => x"2073",
000767 => x"746e",
000768 => x"6f6c",
000769 => x"7469",
000770 => x"6e67",
000771 => x"4067",
000772 => x"6d61",
000773 => x"696c",
000774 => x"2e63",
000775 => x"6f6d",
000776 => x"0d0a",
000777 => x"7777",
000778 => x"772e",
000779 => x"6f70",
000780 => x"656e",
000781 => x"636f",
000782 => x"7265",
000783 => x"732e",
000784 => x"6f72",
000785 => x"672f",
000786 => x"7072",
000787 => x"6f6a",
000788 => x"6563",
000789 => x"742c",
000790 => x"6174",
000791 => x"6c61",
000792 => x"735f",
000793 => x"636f",
000794 => x"7265",
000795 => x"0d0a",
000796 => x"0000",
000797 => x"0d0a",
000798 => x"426f",
000799 => x"6f74",
000800 => x"2070",
000801 => x"6167",
000802 => x"653a",
000803 => x"2030",
000804 => x"7800",
000805 => x"0d0a",
000806 => x"436c",
000807 => x"6f63",
000808 => x"6b28",
000809 => x"487a",
000810 => x"293a",
000811 => x"2030",
000812 => x"7800",
000813 => x"426f",
000814 => x"6f74",
000815 => x"696e",
000816 => x"670d",
000817 => x"0a00",
000818 => x"4275",
000819 => x"726e",
000820 => x"2045",
000821 => x"4550",
000822 => x"524f",
000823 => x"4d0d",
000824 => x"0a00",
000825 => x"4177",
000826 => x"6169",
000827 => x"7469",
000828 => x"6e67",
000829 => x"2069",
000830 => x"6d61",
000831 => x"6765",
000832 => x"2e2e",
000833 => x"2e0d",
000834 => x"0a00",
000835 => x"5374",
000836 => x"6172",
000837 => x"7469",
000838 => x"6e67",
000839 => x"2069",
000840 => x"6d61",
000841 => x"6765",
000842 => x"2000",
000843 => x"446f",
000844 => x"776e",
000845 => x"6c6f",
000846 => x"6164",
000847 => x"2063",
000848 => x"6f6d",
000849 => x"706c",
000850 => x"6574",
000851 => x"650d",
000852 => x"0a00",
000853 => x"5061",
000854 => x"6765",
000855 => x"2028",
000856 => x"3468",
000857 => x"293a",
000858 => x"2024",
000859 => x"0000",
000860 => x"4164",
000861 => x"6472",
000862 => x"2028",
000863 => x"3868",
000864 => x"293a",
000865 => x"2024",
000866 => x"0000",
000867 => x"2377",
000868 => x"6f72",
000869 => x"6473",
000870 => x"2028",
000871 => x"3468",
000872 => x"293a",
000873 => x"2024",
000874 => x"0000",
000875 => x"4368",
000876 => x"6563",
000877 => x"6b73",
000878 => x"756d",
000879 => x"3a20",
000880 => x"2400",
000881 => x"0d0a",
000882 => x"636d",
000883 => x"642f",
000884 => x"626f",
000885 => x"6f74",
000886 => x"2d73",
000887 => x"7769",
000888 => x"7463",
000889 => x"683a",
000890 => x"0d0a",
000891 => x"2030",
000892 => x"2f27",
000893 => x"3030",
000894 => x"273a",
000895 => x"2028",
000896 => x"5265",
000897 => x"2d29",
000898 => x"5374",
000899 => x"6172",
000900 => x"7420",
000901 => x"636f",
000902 => x"6e73",
000903 => x"6f6c",
000904 => x"650d",
000905 => x"0a20",
000906 => x"312f",
000907 => x"2730",
000908 => x"3127",
000909 => x"3a20",
000910 => x"426f",
000911 => x"6f74",
000912 => x"2055",
000913 => x"4152",
000914 => x"540d",
000915 => x"0a20",
000916 => x"322f",
000917 => x"2731",
000918 => x"3027",
000919 => x"3a20",
000920 => x"426f",
000921 => x"6f74",
000922 => x"2045",
000923 => x"4550",
000924 => x"524f",
000925 => x"4d0d",
000926 => x"0a20",
000927 => x"332f",
000928 => x"2731",
000929 => x"3127",
000930 => x"3a20",
000931 => x"426f",
000932 => x"6f74",
000933 => x"206d",
000934 => x"656d",
000935 => x"6f72",
000936 => x"790d",
000937 => x"0a00",
000938 => x"2034",
000939 => x"3a20",
000940 => x"426f",
000941 => x"6f74",
000942 => x"2057",
000943 => x"420d",
000944 => x"0a20",
000945 => x"703a",
000946 => x"2042",
000947 => x"7572",
000948 => x"6e20",
000949 => x"4545",
000950 => x"5052",
000951 => x"4f4d",
000952 => x"0d0a",
000953 => x"2064",
000954 => x"3a20",
000955 => x"5241",
000956 => x"4d20",
000957 => x"6475",
000958 => x"6d70",
000959 => x"0d0a",
000960 => x"2072",
000961 => x"3a20",
000962 => x"5265",
000963 => x"7365",
000964 => x"740d",
000965 => x"0a20",
000966 => x"773a",
000967 => x"2057",
000968 => x"4220",
000969 => x"6475",
000970 => x"6d70",
000971 => x"0d0a",
000972 => x"0000",
000973 => x"636d",
000974 => x"643a",
000975 => x"3e20",
000976 => x"0000",
000977 => x"494d",
000978 => x"4147",
000979 => x"4520",
000980 => x"4552",
000981 => x"5221",
000982 => x"0d0a",
000983 => x"0000",
000984 => x"0d0a",
000985 => x"4952",
000986 => x"5120",
000987 => x"4552",
000988 => x"5221",
000989 => x"0d0a",
000990 => x"0000",
000991 => x"4348",
000992 => x"4543",
000993 => x"4b53",
000994 => x"554d",
000995 => x"2045",
000996 => x"5252",
000997 => x"210d",
000998 => x"0a00",
000999 => x"5350",
001000 => x"492f",
001001 => x"4545",
001002 => x"5052",
001003 => x"4f4d",
001004 => x"2045",
001005 => x"5252",
001006 => x"210d",
001007 => x"0a00",
001008 => x"5742",
001009 => x"2042",
001010 => x"5553",
001011 => x"2045",
001012 => x"5252",
001013 => x"210d",
001014 => x"0a00",
001015 => x"5072",
001016 => x"6573",
001017 => x"7320",
001018 => x"616e",
001019 => x"7920",
001020 => x"6b65",
001021 => x"790d",
001022 => x"0a00",
others => x"0000"