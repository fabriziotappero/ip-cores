--
----- PACKAGE global -----
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE global IS
	SIGNAL gsrnet: std_logic := 'H';
	SIGNAL purnet: std_logic := 'H';
        SIGNAL tsallnet: std_logic := 'H';
END global;

PACKAGE BODY global IS 
END global;


