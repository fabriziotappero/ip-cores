// megafunction wizard: %ALTDDIO_OUT%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altddio_out 

// ============================================================
// File Name: DDR_O.v
// Megafunction Name(s):
// 			altddio_out
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.0 Build 235 06/17/2009 SP 2 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module DDR_O (
	datain_h,
	datain_l,
	outclock,
	dataout);

	input	[5:0]  datain_h;
	input	[5:0]  datain_l;
	input	  outclock;
	output	[5:0]  dataout;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ARESET_MODE NUMERIC "2"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: EXTEND_OE_DISABLE NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: PRIVATE: OE NUMERIC "0"
// Retrieval info: PRIVATE: OE_REG NUMERIC "0"
// Retrieval info: PRIVATE: POWER_UP_HIGH NUMERIC "0"
// Retrieval info: PRIVATE: SRESET_MODE NUMERIC "2"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIDTH NUMERIC "6"
// Retrieval info: CONSTANT: EXTEND_OE_DISABLE STRING "UNUSED"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altddio_out"
// Retrieval info: CONSTANT: OE_REG STRING "UNUSED"
// Retrieval info: CONSTANT: POWER_UP_HIGH STRING "OFF"
// Retrieval info: CONSTANT: WIDTH NUMERIC "6"
// Retrieval info: USED_PORT: datain_h 0 0 6 0 INPUT NODEFVAL datain_h[5..0]
// Retrieval info: USED_PORT: datain_l 0 0 6 0 INPUT NODEFVAL datain_l[5..0]
// Retrieval info: USED_PORT: dataout 0 0 6 0 OUTPUT NODEFVAL dataout[5..0]
// Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL outclock
// Retrieval info: CONNECT: @datain_h 0 0 6 0 datain_h 0 0 6 0
// Retrieval info: CONNECT: @datain_l 0 0 6 0 datain_l 0 0 6 0
// Retrieval info: CONNECT: dataout 0 0 6 0 @dataout 0 0 6 0
// Retrieval info: CONNECT: @outclock 0 0 0 0 outclock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR_O_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
