// sdram_tb.v

// Generated using ACDS version 13.0 156 at 2013.08.12.18:22:22

`timescale 1 ps / 1 ps
module sdram_tb (
	);

	wire         sdram_inst_clk_bfm_clk_clk;                  // sdram_inst_clk_bfm:clk -> [sdram_inst:clk_clk, sdram_inst_reset_bfm:clk]
	wire         sdram_inst_reset_bfm_reset_reset;            // sdram_inst_reset_bfm:reset -> sdram_inst:reset_reset_n
	wire         sdram_inst_sdram_wire_cs_n;                  // sdram_inst:sdram_wire_cs_n -> sdram_controller_my_partner:zs_cs_n
	wire   [1:0] sdram_inst_sdram_wire_ba;                    // sdram_inst:sdram_wire_ba -> sdram_controller_my_partner:zs_ba
	wire   [3:0] sdram_inst_sdram_wire_dqm;                   // sdram_inst:sdram_wire_dqm -> sdram_controller_my_partner:zs_dqm
	wire         sdram_inst_sdram_wire_cke;                   // sdram_inst:sdram_wire_cke -> sdram_controller_my_partner:zs_cke
	wire  [12:0] sdram_inst_sdram_wire_addr;                  // sdram_inst:sdram_wire_addr -> sdram_controller_my_partner:zs_addr
	wire         sdram_inst_sdram_wire_we_n;                  // sdram_inst:sdram_wire_we_n -> sdram_controller_my_partner:zs_we_n
	wire         sdram_inst_sdram_wire_ras_n;                 // sdram_inst:sdram_wire_ras_n -> sdram_controller_my_partner:zs_ras_n
	wire         sdram_inst_sdram_wire_cas_n;                 // sdram_inst:sdram_wire_cas_n -> sdram_controller_my_partner:zs_cas_n
	wire  [31:0] sdram_controller_my_partner_conduit_dq;      // [] -> [sdram_controller_my_partner:zs_dq, sdram_inst:sdram_wire_dq]
	wire         sdram_controller_my_partner_clk_bfm_clk_clk; // sdram_controller_my_partner_clk_bfm:clk -> sdram_controller_my_partner:clk

	sdram sdram_inst (
		.clk_clk                (sdram_inst_clk_bfm_clk_clk),             //        clk.clk
		.reset_reset_n          (sdram_inst_reset_bfm_reset_reset),       //      reset.reset_n
		.sdram_s1_address       (),                                       //   sdram_s1.address
		.sdram_s1_byteenable_n  (),                                       //           .byteenable_n
		.sdram_s1_chipselect    (),                                       //           .chipselect
		.sdram_s1_writedata     (),                                       //           .writedata
		.sdram_s1_read_n        (),                                       //           .read_n
		.sdram_s1_write_n       (),                                       //           .write_n
		.sdram_s1_readdata      (),                                       //           .readdata
		.sdram_s1_readdatavalid (),                                       //           .readdatavalid
		.sdram_s1_waitrequest   (),                                       //           .waitrequest
		.sdram_wire_addr        (sdram_inst_sdram_wire_addr),             // sdram_wire.addr
		.sdram_wire_ba          (sdram_inst_sdram_wire_ba),               //           .ba
		.sdram_wire_cas_n       (sdram_inst_sdram_wire_cas_n),            //           .cas_n
		.sdram_wire_cke         (sdram_inst_sdram_wire_cke),              //           .cke
		.sdram_wire_cs_n        (sdram_inst_sdram_wire_cs_n),             //           .cs_n
		.sdram_wire_dq          (sdram_controller_my_partner_conduit_dq), //           .dq
		.sdram_wire_dqm         (sdram_inst_sdram_wire_dqm),              //           .dqm
		.sdram_wire_ras_n       (sdram_inst_sdram_wire_ras_n),            //           .ras_n
		.sdram_wire_we_n        (sdram_inst_sdram_wire_we_n),             //           .we_n
		.sdram_clk_clk          ()                                        //  sdram_clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sdram_inst_clk_bfm (
		.clk (sdram_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sdram_inst_reset_bfm (
		.reset (sdram_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sdram_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_sdram_partner_module sdram_controller_my_partner (
		.clk      (sdram_controller_my_partner_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (sdram_controller_my_partner_conduit_dq),      // conduit.dq
		.zs_addr  (sdram_inst_sdram_wire_addr),                  //        .addr
		.zs_ba    (sdram_inst_sdram_wire_ba),                    //        .ba
		.zs_cas_n (sdram_inst_sdram_wire_cas_n),                 //        .cas_n
		.zs_cke   (sdram_inst_sdram_wire_cke),                   //        .cke
		.zs_cs_n  (sdram_inst_sdram_wire_cs_n),                  //        .cs_n
		.zs_dqm   (sdram_inst_sdram_wire_dqm),                   //        .dqm
		.zs_ras_n (sdram_inst_sdram_wire_ras_n),                 //        .ras_n
		.zs_we_n  (sdram_inst_sdram_wire_we_n)                   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sdram_controller_my_partner_clk_bfm (
		.clk (sdram_controller_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
