--------------------------------------------------------------------------------
-- Object        : Package work.package_txt_utilities
-- Last modified : Sun Dec 04 20:16:51 2011.
--------------------------------------------------------------------------------



library ieee, std;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;
---------------------------------------------------------------------------------------------------------------
-- Library declaration
---------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;

---------------------------------------------------------------------------------------------------------------
-- Package declaration
---------------------------------------------------------------------------------------------------------------
package package_txt_utilities is

    -- prints a message to the screen
    procedure fwrite(text: string);

    -- prints the message when active
    -- useful for debug switches
    procedure fwrite(active: boolean; text: string);
    
    --------------------------------------------------
    -- functions to convert strings into data type
    --------------------------------------------------
    -- converts a character into std_logic
    function to_std_logic(c: character) return std_logic; 
    
    -- converts a string into std_logic_vector
    function bin_string_to_std_logic_vector(s: string) return std_logic_vector;    
    function hex_string_to_std_logic_vector(s: string) return std_logic_vector;    

    -------------------------------------------
    -- functions to convert data type to string
    -------------------------------------------
    -- converts std_logic into a character
    function to_char(sl: std_logic) return character;

    -- converts std_logic into a string (1 to 1)
    function to_string(sl: std_logic) return string;

    -- converts std_logic_vector into a string (binary base)
    function to_string(slv: std_logic_vector) return string;

    -- converts boolean into a string
    function to_string(b: boolean) return string;

    -- converts an integer into a single character
    -- (can also be used for hex conversion and other bases)
    function to_char(int: integer) return character;

    -- converts integer into string using specified base
    function to_string(int: integer; base: integer) return string;

    -- converts integer to string, using base 10
    function to_string(int: integer) return string;

    -- convert std_logic_vector into a string in hex format
    function to_hexstring(slv: std_logic_vector) return string;

    -------------------------------------------
    -- functions to manipulate strings
    -------------------------------------------
    -- convert a character to upper case
    function to_upper(c: character) return character;

    -- convert a character to lower case
    function to_lower(c: character) return character;

    -- convert a string to upper case
    function to_upper(s: string) return string;

    -- convert a string to lower case
    function to_lower(s: string) return string;

    --------------------------------------------------
    -- file I/O
    --------------------------------------------------
    -- read variable length string from input file
    procedure fread(file in_file: TEXT; 
                       res_string: out string);
    
    -- print string to a file and start new line
    procedure fwrite(file out_file: TEXT;
                    new_string: in  string);
    
    -- print character to a file and start new line
    procedure fwrite(file out_file: TEXT;
                    char:       in  character);

    -- print string to a file and start new line
    procedure fdebug(level: in integer;
                    threshold: in integer;
                    file out_file: TEXT;
                    new_string: in  string);
end package_txt_utilities;

---------------------------------------------------------------------------------------------------------------
-- Package definitions
---------------------------------------------------------------------------------------------------------------
package body package_txt_utilities is

--=============================================================================================================
-- Process		: print
-- Description	: prints text to the screen
--=============================================================================================================

   procedure fwrite(text: string) is
     variable msg_line: line;
     begin
       write(msg_line, text);
       writeline(output, msg_line);
   end fwrite;

--=============================================================================================================
-- Process		: print
-- Description	: prints text to the screen when active
--=============================================================================================================
procedure fwrite(active: boolean; text: string)  is
     begin
      if active then
         fwrite(text);
      end if;
   end fwrite;

--=============================================================================================================
-- Process		: chr
-- Description	: converts std_logic into a character
--=============================================================================================================
function to_char(sl: std_logic) return character is
    variable c: character;
    begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
    return c;
   end to_char;

--=============================================================================================================
-- Process		: str
-- Description	: converts std_logic into a string (1 to 1)
--=============================================================================================================
function to_string(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
        s(1) := to_char(sl);
        return s;
   end to_string;

--=============================================================================================================
-- Process		: str
-- Description	: converts std_logic_vector into a string (binary base)
--=============================================================================================================
function to_string(slv: std_logic_vector) return string is
     variable result : string (1 to slv'length);
     variable r : integer;
   begin
     r := 1;
     for i in slv'range loop
        result(r) := to_char(slv(i));
        r := r + 1;
     end loop;
     return result;
   end to_string;

--=============================================================================================================
-- Process		: str
-- Description	: 
--=============================================================================================================
function to_string(b: boolean) return string is

    begin
       if b then
          return "true";
      else
        return "false";
       end if;
    end to_string;

--=============================================================================================================
-- Process		: chr
-- Description	: converts an integer into a character 
--=============================================================================================================
function to_char(int: integer) return character is
    variable c: character;
   begin
        case int is
          when  0 => c := '0';
          when  1 => c := '1';
          when  2 => c := '2';
          when  3 => c := '3';
          when  4 => c := '4';
          when  5 => c := '5';
          when  6 => c := '6';
          when  7 => c := '7';
          when  8 => c := '8';
          when  9 => c := '9';
          when 10 => c := 'A';
          when 11 => c := 'B';
          when 12 => c := 'C';
          when 13 => c := 'D';
          when 14 => c := 'E';
          when 15 => c := 'F';
          when 16 => c := 'G';
          when 17 => c := 'H';
          when 18 => c := 'I';
          when 19 => c := 'J';
          when 20 => c := 'K';
          when 21 => c := 'L';
          when 22 => c := 'M';
          when 23 => c := 'N';
          when 24 => c := 'O';
          when 25 => c := 'P';
          when 26 => c := 'Q';
          when 27 => c := 'R';
          when 28 => c := 'S';
          when 29 => c := 'T';
          when 30 => c := 'U';
          when 31 => c := 'V';
          when 32 => c := 'W';
          when 33 => c := 'X';
          when 34 => c := 'Y';
          when 35 => c := 'Z';
          when others => c := '?';
        end case;
        return c;
    end to_char;

--=============================================================================================================
-- Process		: str
-- Description	: convert integer to string using specified base 
--=============================================================================================================
function to_string(int: integer; base: integer) return string is

    variable temp:      string(1 to 10);
    variable num:       integer;
    variable abs_int:   integer;
    variable len:       integer := 1;
    variable power:     integer := 1;

   begin

    -- bug fix for negative numbers
    abs_int := abs(int);

    num     := abs_int;

    while num >= base loop                     -- Determine how many
      len := len + 1;                          -- characters required
      num := num / base;                       -- to represent the
    end loop ;                                 -- number.

    for i in len downto 1 loop                 -- Convert the number to
      temp(i) := to_char(abs_int/power mod base);  -- a string starting
      power := power * base;                   -- with the right hand
    end loop ;                                 -- side.

    -- return result and add sign if required
    if int < 0 then
       return '-'& temp(1 to len);
     else
       return temp(1 to len);
    end if;

   end to_string;

--=============================================================================================================
-- Process		: str
-- Description	: convert integer to string, using base 10
--=============================================================================================================
function to_string(int: integer) return string is

   begin

    return to_string(int, 10) ;

   end to_string;

--=============================================================================================================
-- Process		: hstr
-- Description	: converts a std_logic_vector into a hex string
--=============================================================================================================
function to_hexstring(slv: std_logic_vector) return string is
       variable hexlen: integer;
       variable longslv : std_logic_vector(67 downto 0) := (others => '0');
       variable hex : string(1 to 16);
       variable fourbit : std_logic_vector(3 downto 0);
     begin
       hexlen := (slv'left+1)/4;
       if (slv'left+1) mod 4 /= 0 then
         hexlen := hexlen + 1;
       end if;
       longslv(slv'left downto 0) := slv;
       for i in (hexlen -1) downto 0 loop
         fourbit := longslv(((i*4)+3) downto (i*4));
         case fourbit is
           when "0000" => hex(hexlen -I) := '0';
           when "0001" => hex(hexlen -I) := '1';
           when "0010" => hex(hexlen -I) := '2';
           when "0011" => hex(hexlen -I) := '3';
           when "0100" => hex(hexlen -I) := '4';
           when "0101" => hex(hexlen -I) := '5';
           when "0110" => hex(hexlen -I) := '6';
           when "0111" => hex(hexlen -I) := '7';
           when "1000" => hex(hexlen -I) := '8';
           when "1001" => hex(hexlen -I) := '9';
           when "1010" => hex(hexlen -I) := 'A';
           when "1011" => hex(hexlen -I) := 'B';
           when "1100" => hex(hexlen -I) := 'C';
           when "1101" => hex(hexlen -I) := 'D';
           when "1110" => hex(hexlen -I) := 'E';
           when "1111" => hex(hexlen -I) := 'F';
           when "ZZZZ" => hex(hexlen -I) := 'z';
           when "UUUU" => hex(hexlen -I) := 'u';
           when "XXXX" => hex(hexlen -I) := 'x';
           when others => hex(hexlen -I) := '?';
         end case;
       end loop;
       return hex(1 to hexlen);
     end to_hexstring;

--=============================================================================================================
-- Process		: to_upper
-- Description	: convert a character to upper case
--=============================================================================================================
function to_upper(c: character) return character is

      variable u: character;

    begin

       case c is
        when 'a' => u := 'A';
        when 'b' => u := 'B';
        when 'c' => u := 'C';
        when 'd' => u := 'D';
        when 'e' => u := 'E';
        when 'f' => u := 'F';
        when 'g' => u := 'G';
        when 'h' => u := 'H';
        when 'i' => u := 'I';
        when 'j' => u := 'J';
        when 'k' => u := 'K';
        when 'l' => u := 'L';
        when 'm' => u := 'M';
        when 'n' => u := 'N';
        when 'o' => u := 'O';
        when 'p' => u := 'P';
        when 'q' => u := 'Q';
        when 'r' => u := 'R';
        when 's' => u := 'S';
        when 't' => u := 'T';
        when 'u' => u := 'U';
        when 'v' => u := 'V';
        when 'w' => u := 'W';
        when 'x' => u := 'X';
        when 'y' => u := 'Y';
        when 'z' => u := 'Z';
        when others => u := c;
    end case;

      return u;

   end to_upper;

--=============================================================================================================
-- Process		: to_lower
-- Description	: convert a character to lower case
--=============================================================================================================
function to_lower(c: character) return character is

      variable l: character;

    begin

       case c is
        when 'A' => l := 'a';
        when 'B' => l := 'b';
        when 'C' => l := 'c';
        when 'D' => l := 'd';
        when 'E' => l := 'e';
        when 'F' => l := 'f';
        when 'G' => l := 'g';
        when 'H' => l := 'h';
        when 'I' => l := 'i';
        when 'J' => l := 'j';
        when 'K' => l := 'k';
        when 'L' => l := 'l';
        when 'M' => l := 'm';
        when 'N' => l := 'n';
        when 'O' => l := 'o';
        when 'P' => l := 'p';
        when 'Q' => l := 'q';
        when 'R' => l := 'r';
        when 'S' => l := 's';
        when 'T' => l := 't';
        when 'U' => l := 'u';
        when 'V' => l := 'v';
        when 'W' => l := 'w';
        when 'X' => l := 'x';
        when 'Y' => l := 'y';
        when 'Z' => l := 'z';
        when others => l := c;
    end case;

      return l;

   end to_lower;

--=============================================================================================================
-- Process		: to_upper
-- Description	: convert a string to upper case
--=============================================================================================================
function to_upper(s: string) return string is

     variable uppercase: string (s'range);

   begin

     for i in s'range loop
        uppercase(i):= to_upper(s(i));
     end loop;
     return uppercase;

   end to_upper;

--=============================================================================================================
-- Process		: to_lower
-- Description	: convert a string to lower case
--=============================================================================================================
function to_lower(s: string) return string is

     variable lowercase: string (s'range);

   begin

     for i in s'range loop
        lowercase(i):= to_lower(s(i));
     end loop;
     return lowercase;

   end to_lower;

--=============================================================================================================
-- Process		: to_std_logic
-- Description	: converts a character into a std_logic
--=============================================================================================================
function to_std_logic(c: character) return std_logic is 
    variable sl: std_logic;
    begin
      case c is
        when 'U' => 
           sl := 'U'; 
        when 'X' =>
           sl := 'X';
        when '0' => 
           sl := '0';
        when '1' => 
           sl := '1';
        when 'Z' => 
           sl := 'Z';
        when 'W' => 
           sl := 'W';
        when 'L' => 
           sl := 'L';
        when 'H' => 
           sl := 'H';
        when '-' => 
           sl := '-';
        when others =>
           sl := 'X'; 
    end case;
   return sl;
  end to_std_logic;

--=============================================================================================================
-- Process		: to_std_logic_vector
-- Description	: converts a string into std_logic_vector
--=============================================================================================================
function bin_string_to_std_logic_vector(s: string) return std_logic_vector is 
  variable slv: std_logic_vector(s'high-s'low downto 0);
  variable k: integer;
begin
   k := s'high-s'low;
  for i in s'range loop
     slv(k) := to_std_logic(s(i));
     k      := k - 1;
  end loop;
  return slv;
end bin_string_to_std_logic_vector;                                       

function hex_string_to_std_logic_vector(s: string) return std_logic_vector is 
    variable slv: std_logic_vector(4*s'high-1 downto 0);
begin
    for i in s'range loop
      case s(i) is
        when '0'    =>  slv(4*i-1 downto 4*i-4) := "0000";
        when '1'    =>  slv(4*i-1 downto 4*i-4) := "0001";
        when '2'    =>  slv(4*i-1 downto 4*i-4) := "0010";
        when '3'    =>  slv(4*i-1 downto 4*i-4) := "0011";
        when '4'    =>  slv(4*i-1 downto 4*i-4) := "0100";
        when '5'    =>  slv(4*i-1 downto 4*i-4) := "0101";
        when '6'    =>  slv(4*i-1 downto 4*i-4) := "0110";
        when '7'    =>  slv(4*i-1 downto 4*i-4) := "0111";
        when '8'    =>  slv(4*i-1 downto 4*i-4) := "1000";
        when '9'    =>  slv(4*i-1 downto 4*i-4) := "1001";
        when 'A'    =>  slv(4*i-1 downto 4*i-4) := "1010";
        when 'B'    =>  slv(4*i-1 downto 4*i-4) := "1011";
        when 'C'    =>  slv(4*i-1 downto 4*i-4) := "1100";
        when 'D'    =>  slv(4*i-1 downto 4*i-4) := "1101";
        when 'E'    =>  slv(4*i-1 downto 4*i-4) := "1110";
        when 'F'    =>  slv(4*i-1 downto 4*i-4) := "1111";
        when 'a'    =>  slv(4*i-1 downto 4*i-4) := "1010";
        when 'b'    =>  slv(4*i-1 downto 4*i-4) := "1011";
        when 'c'    =>  slv(4*i-1 downto 4*i-4) := "1100";
        when 'd'    =>  slv(4*i-1 downto 4*i-4) := "1101";
        when 'e'    =>  slv(4*i-1 downto 4*i-4) := "1110";
        when 'f'    =>  slv(4*i-1 downto 4*i-4) := "1111";
        when others =>  slv(4*i-1 downto 4*i-4) := "0000";
      end case;
    end loop;
  return slv;
end hex_string_to_std_logic_vector;   


                                       
--=============================================================================================================
-- Process		: fread
-- Description	: 
--=============================================================================================================
procedure fread(file in_file: TEXT; 
                   res_string: out string) is
       
       variable l:         line;
       variable c:         character;
       variable is_string: boolean;
       
   begin
           
     readline(in_file, l);
     -- clear the contents of the result string
     for i in res_string'range loop
         res_string(i) := ' ';
     end loop;   
     -- read all characters of the line, up to the length  
     -- of the results string
     for i in res_string'range loop
        read(l, c, is_string);
        res_string(i) := c;
        if not is_string then -- found end of line
           exit;
        end if;   
     end loop; 
                     
end fread;

--=============================================================================================================
-- Process		: print
-- Description	: print string to a file
--=============================================================================================================
procedure fwrite(file out_file: TEXT;
                new_string: in  string) is
       
       variable l: line;
       
   begin
      
     write(l, new_string);
     writeline(out_file, l);
                     
end fwrite;

--=============================================================================================================
-- Process		: print
-- Description	: print string to a file
--=============================================================================================================
procedure fdebug(level: in integer;
                 threshold: in integer;
                 file out_file: TEXT;
                 new_string: in  string) is
       
       variable l: line;
       
   begin
    if level <= threshold then
      write(l, new_string);
      writeline(out_file, l);
    end if;
                     
end fdebug;

--=============================================================================================================
-- Process		: print
-- Description	: print character to a file and start new line 
--=============================================================================================================
procedure fwrite(file out_file: TEXT;
                char: in  character) is
       
       variable l: line;
       
   begin
      
     write(l, char);
     writeline(out_file, l);
                     
end fwrite;

--=============================================================================================================
-- Process		: str_write
-- Description	: appends contents of a string to a file until line feed occurs (LF is considered to be the end of the string)
--=============================================================================================================
procedure str_write(file out_file: TEXT; 
                    new_string: in  string) is
 begin
      
   for i in new_string'range loop
      fwrite(out_file, new_string(i));
      if new_string(i) = LF then -- end of string
         exit;
      end if;
   end loop;               

end str_write;
end package_txt_utilities;




