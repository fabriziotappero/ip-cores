//Jul.5.2004 reduce critical path cell
//Apr.5.2005 always @(*)
`include "define.h"
module 
shifter(a,c,shift_func,shift_amount);
	input [31:0] a;
	output [31:0] c;
	input [1:0] shift_func;
	input [4:0] shift_amount;

	 reg [31:0] c;

	always @ (*) begin //
		 if (!shift_func[1]  ) begin
			case (shift_amount[4:0] )
				5'b00000: c=a;
				5'b00001: c={a[30:0],1'b0};
				5'b00010: c={a[29:0],2'b00};
				5'b00011: c={a[28:0],3'b000};
				5'b00100: c={a[27:0],4'b0000};
				5'b00101: c={a[26:0],5'b0_0000};
				5'b00110: c={a[25:0],6'b00_0000};
				5'b00111: c={a[24:0],7'b000_0000};
				5'b01000: c={a[23:0],8'b0000_0000};
				5'b01001: c={a[22:0],9'b0_0000_0000};
				5'b01010: c={a[21:0],10'b00_0000_0000};
				5'b01011: c={a[20:0],11'b000_0000_0000};
				5'b01100: c={a[19:0],12'b0000_0000_0000};
				5'b01101: c={a[18:0],13'b0_0000_0000_0000};
				5'b01110: c={a[17:0],14'b00_0000_0000_0000};
			      5'b01111: c={a[16:0],15'b000_0000_0000_0000};
				5'b10000: c={a[15:0],16'b0000_0000_0000_0000};
				5'b10001: c={a[14:0],16'b0000_0000_0000_0000,1'b0};
				5'b10010: c={a[13:0],16'b0000_0000_0000_0000,2'b00};
				5'b10011: c={a[12:0],16'b0000_0000_0000_0000,3'b000};
				5'b10100: c={a[11:0],16'b0000_0000_0000_0000,4'b0000};
				5'b10101: c={a[10:0],16'b0000_0000_0000_0000,5'b0_0000};
				5'b10110: c={a[9:0],16'b0000_0000_0000_0000,6'b00_0000};
				5'b10111: c={a[8:0],16'b0000_0000_0000_0000,7'b000_0000};
				5'b11000: c={a[7:0],16'b0000_0000_0000_0000,8'b0000_0000};
				5'b11001: c={a[6:0],16'b0000_0000_0000_0000,9'b0_0000_0000};
				5'b11010: c={a[5:0],16'b0000_0000_0000_0000,10'b00_0000_0000};
				5'b11011: c={a[4:0],16'b0000_0000_0000_0000,11'b000_0000_0000};
				5'b11100: c={a[3:0],16'b0000_0000_0000_0000,12'b0000_0000_0000};
				5'b11101: c={a[2:0],16'b0000_0000_0000_0000,13'b0_0000_0000_0000};
				5'b11110: c={a[1:0],16'b0000_0000_0000_0000,14'b00_0000_0000_0000};
			      5'b11111: c={a[0],16'b0000_0000_0000_0000,15'b000_0000_0000_0000};
			endcase
		end else if (shift_func==`SHIFT_RIGHT_UNSIGNED) begin
			case (shift_amount)
				5'b00000: c=a;
				5'b00001: c={1'b0,a[31:1]};
				5'b00010: c={2'b00,a[31:2]};
				5'b00011: c={3'b000,a[31:3]};
				5'b00100: c={4'b0000,a[31:4]};
				5'b00101: c={5'b0_0000,a[31:5]};
				5'b00110: c={6'b00_0000,a[31:6]};
				5'b00111: c={7'b000_0000,a[31:7]};
				5'b01000: c={8'b0000_0000,a[31:8]};
				5'b01001: c={9'b0_0000_0000,a[31:9]};
				5'b01010: c={10'b00_0000_0000,a[31:10]};
				5'b01011: c={11'b000_0000_0000,a[31:11]};			
				5'b01100: c={12'b0000_0000_0000,a[31:12]};
				5'b01101: c={13'b0_0000_0000_0000,a[31:13]};					
				5'b01110: c={14'b00_0000_0000_0000,a[31:14]};
			      5'b01111: c={15'b000_0000_0000_0000,a[31:15]};		
				5'b10000: c={16'b0000_0000_0000_0000,a[31:16]};
				5'b10001: c={16'b0000_0000_0000_0000,1'b0,a[31:17]};
				5'b10010: c={16'b0000_0000_0000_0000,2'b00,a[31:18]};
				5'b10011: c={16'b0000_0000_0000_0000,3'b000,a[31:19]};
				5'b10100: c={16'b0000_0000_0000_0000,4'b0000,a[31:20]};
				5'b10101: c={16'b0000_0000_0000_0000,5'b0_0000,a[31:21]};
				5'b10110: c={16'b0000_0000_0000_0000,6'b00_0000,a[31:22]};
				5'b10111: c={16'b0000_0000_0000_0000,7'b000_0000,a[31:23]};
				5'b11000: c={16'b0000_0000_0000_0000,8'b0000_0000,a[31:24]};
				5'b11001: c={16'b0000_0000_0000_0000,9'b0_0000_0000,a[31:25]};
				5'b11010: c={16'b0000_0000_0000_0000,10'b00_0000_0000,a[31:26]};
				5'b11011: c={16'b0000_0000_0000_0000,11'b000_0000_0000,a[31:27]};			
				5'b11100: c={16'b0000_0000_0000_0000,12'b0000_0000_0000,a[31:28]};
				5'b11101: c={16'b0000_0000_0000_0000,13'b0_0000_0000_0000,a[31:29]};					
				5'b11110: c={16'b0000_0000_0000_0000,14'b00_0000_0000_0000,a[31:30]};
			      5'b11111: c={16'b0000_0000_0000_0000,15'b000_0000_0000_0000,a[31:31]};		
			endcase
		end else begin// SHIFT_RIGHT_SIGNED
			case (shift_amount)	
				5'b00000: c=a;
				5'b00001: c={a[31],a[31:1]};
				5'b00010: c={{2{a[31]}},a[31:2]};
				5'b00011: c={{3{a[31]}},a[31:3]};
				5'b00100: c={{4{a[31]}},a[31:4]};
				5'b00101: c={{5{a[31]}},a[31:5]};
				5'b00110: c={{6{a[31]}},a[31:6]};
				5'b00111: c={{7{a[31]}},a[31:7]};
				5'b01000: c={{8{a[31]}},a[31:8]};
				5'b01001: c={{9{a[31]}},a[31:9]};
				5'b01010: c={{10{a[31]}},a[31:10]};
				5'b01011: c={{11{a[31]}},a[31:11]};			
				5'b01100: c={{12{a[31]}},a[31:12]};
				5'b01101: c={{13{a[31]}},a[31:13]};					
				5'b01110: c={{14{a[31]}},a[31:14]};
			      5'b01111: c={{15{a[31]}},a[31:15]};		
				5'b10000: c={{16{a[31]}},a[31:16]};
				5'b10001: c={{17{a[31]}},a[31:17]};
				5'b10010: c={{18{a[31]}},a[31:18]};
				5'b10011: c={{19{a[31]}},a[31:19]};
				5'b10100: c={{20{a[31]}},a[31:20]};
				5'b10101: c={{21{a[31]}},a[31:21]};
				5'b10110: c={{22{a[31]}},a[31:22]};
				5'b10111: c={{23{a[31]}},a[31:23]};
				5'b11000: c={{24{a[31]}},a[31:24]};
				5'b11001: c={{25{a[31]}},a[31:25]};
				5'b11010: c={{26{a[31]}},a[31:26]};
				5'b11011: c={{27{a[31]}},a[31:27]};			
				5'b11100: c={{28{a[31]}},a[31:28]};
				5'b11101: c={{29{a[31]}},a[31:29]};					
				5'b11110: c={{30{a[31]}},a[31:30]};
			      5'b11111: c={{31{a[31]}},a[31:31]};		
			endcase
		end
	end






endmodule