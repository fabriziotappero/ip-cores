-- SSRAM controller
  constant CFG_SSCTRL  	 : integer := CONFIG_SSCTRL;
  constant CFG_SSCTRLP16 : integer := CONFIG_SSCTRL_PROM16;

