-------------------------------------------------------------------------------
--
-- SD/MMC Bootloader
--
-- $Id: spi_counter-c.vhd 77 2009-04-01 19:53:14Z arniml $
--
-------------------------------------------------------------------------------

configuration spi_counter_rtl_c0 of spi_counter is

  for rtl
  end for;

end spi_counter_rtl_c0;
