module bootrom(clk,adr,romo);
input clk;
input [31:0] adr;
output [15:0] romo;
reg [15:0] romo;
reg [15:0] romout;
always @(adr)
case(adr & 32'hFFFFFFFE)
32'hFFFF1000: romout <= 16'h564C;
32'hFFFF1002: romout <= 16'h4944;
32'hFFFF1004: romout <= 16'h0010;
32'hFFFF1006: romout <= 16'h0000;
32'hFFFF1008: romout <= 16'h0020;
32'hFFFF100A: romout <= 16'h0000;
32'hFFFF100C: romout <= 16'h0000;
32'hFFFF100E: romout <= 16'h0000;
32'hFFFF1010: romout <= 16'h0000;
32'hFFFF1012: romout <= 16'h0000;
32'hFFFF1014: romout <= 16'hFFFF;
32'hFFFF1016: romout <= 16'h1074;
32'hFFFF1018: romout <= 16'hFFFF;
32'hFFFF101A: romout <= 16'h1084;
32'hFFFF101C: romout <= 16'h0000;
32'hFFFF101E: romout <= 16'h0003;
32'hFFFF1020: romout <= 16'hFFFF;
32'hFFFF1022: romout <= 16'h1A5E;
32'hFFFF1024: romout <= 16'h4D4F;
32'hFFFF1026: romout <= 16'h4E49;
32'hFFFF1028: romout <= 16'h544F;
32'hFFFF102A: romout <= 16'h5220;
32'hFFFF102C: romout <= 16'h0000;
32'hFFFF102E: romout <= 16'h0800;
32'hFFFF1030: romout <= 16'h0000;
32'hFFFF1032: romout <= 16'h0000;
32'hFFFF1034: romout <= 16'h0000;
32'hFFFF1036: romout <= 16'h0000;
32'hFFFF1038: romout <= 16'h0000;
32'hFFFF103A: romout <= 16'h0001;
32'hFFFF103C: romout <= 16'hFFFF;
32'hFFFF103E: romout <= 16'h2400;
32'hFFFF1040: romout <= 16'h5449;
32'hFFFF1042: romout <= 16'h4E59;
32'hFFFF1044: romout <= 16'h2042;
32'hFFFF1046: romout <= 16'h4153;
32'hFFFF1048: romout <= 16'h0000;
32'hFFFF104A: romout <= 16'h0800;
32'hFFFF104C: romout <= 16'h0000;
32'hFFFF104E: romout <= 16'h0000;
32'hFFFF1050: romout <= 16'h0000;
32'hFFFF1052: romout <= 16'h0000;
32'hFFFF1054: romout <= 16'h0001;
32'hFFFF1056: romout <= 16'h0002;
32'hFFFF1058: romout <= 16'hFFFF;
32'hFFFF105A: romout <= 16'h12EC;
32'hFFFF105C: romout <= 16'h4944;
32'hFFFF105E: romout <= 16'h4C45;
32'hFFFF1060: romout <= 16'h5441;
32'hFFFF1062: romout <= 16'h534B;
32'hFFFF1064: romout <= 16'h0000;
32'hFFFF1066: romout <= 16'h0400;
32'hFFFF1068: romout <= 16'h0000;
32'hFFFF106A: romout <= 16'h0000;
32'hFFFF106C: romout <= 16'h0000;
32'hFFFF106E: romout <= 16'h0000;
32'hFFFF1070: romout <= 16'h0001;
32'hFFFF1072: romout <= 16'h0003;
32'hFFFF1074: romout <= 16'hFFFF;
32'hFFFF1076: romout <= 16'h16B0;
32'hFFFF1078: romout <= 16'hFFFF;
32'hFFFF107A: romout <= 16'h16D4;
32'hFFFF107C: romout <= 16'hFFFF;
32'hFFFF107E: romout <= 16'h1680;
32'hFFFF1080: romout <= 16'hFFFF;
32'hFFFF1082: romout <= 16'h169A;
32'hFFFF1084: romout <= 16'h0000;
32'hFFFF1086: romout <= 16'h0200;
32'hFFFF1100: romout <= 16'h31FC;
32'hFFFF1102: romout <= 16'h00CE;
32'hFFFF1104: romout <= 16'h0414;
32'hFFFF1106: romout <= 16'h11FC;
32'hFFFF1108: romout <= 16'h0001;
32'hFFFF110A: romout <= 16'h041C;
32'hFFFF110C: romout <= 16'h4EB9;
32'hFFFF110E: romout <= 16'hFFFF;
32'hFFFF1110: romout <= 16'h18E8;
32'hFFFF1112: romout <= 16'h4278;
32'hFFFF1114: romout <= 16'h0418;
32'hFFFF1116: romout <= 16'h4278;
32'hFFFF1118: romout <= 16'h041A;
32'hFFFF111A: romout <= 16'h43F9;
32'hFFFF111C: romout <= 16'hFFFF;
32'hFFFF111E: romout <= 16'h1238;
32'hFFFF1120: romout <= 16'h4EB9;
32'hFFFF1122: romout <= 16'hFFFF;
32'hFFFF1124: romout <= 16'h1858;
32'hFFFF1126: romout <= 16'h47F9;
32'hFFFF1128: romout <= 16'hFFFF;
32'hFFFF112A: romout <= 16'h1132;
32'hFFFF112C: romout <= 16'h4EF9;
32'hFFFF112E: romout <= 16'hFFFF;
32'hFFFF1130: romout <= 16'h1F52;
32'hFFFF1132: romout <= 16'h2079;
32'hFFFF1134: romout <= 16'hFFFF;
32'hFFFF1136: romout <= 16'h2420;
32'hFFFF1138: romout <= 16'h4E60;
32'hFFFF113A: romout <= 16'h31FC;
32'hFFFF113C: romout <= 16'h00CE;
32'hFFFF113E: romout <= 16'h0414;
32'hFFFF1140: romout <= 16'h11FC;
32'hFFFF1142: romout <= 16'h0001;
32'hFFFF1144: romout <= 16'h041C;
32'hFFFF1146: romout <= 16'h4278;
32'hFFFF1148: romout <= 16'h0418;
32'hFFFF114A: romout <= 16'h4278;
32'hFFFF114C: romout <= 16'h041A;
32'hFFFF114E: romout <= 16'h223C;
32'hFFFF1150: romout <= 16'h0000;
32'hFFFF1152: romout <= 16'h8000;
32'hFFFF1154: romout <= 16'h41F9;
32'hFFFF1156: romout <= 16'hFFD8;
32'hFFFF1158: romout <= 16'h0000;
32'hFFFF115A: romout <= 16'h2039;
32'hFFFF115C: romout <= 16'hFFDC;
32'hFFFF115E: romout <= 16'h0C00;
32'hFFFF1160: romout <= 16'h30C0;
32'hFFFF1162: romout <= 16'h5381;
32'hFFFF1164: romout <= 16'h66F4;
32'hFFFF1166: romout <= 16'h41F9;
32'hFFFF1168: romout <= 16'hFFFF;
32'hFFFF116A: romout <= 16'h2022;
32'hFFFF116C: romout <= 16'h21C8;
32'hFFFF116E: romout <= 16'h0008;
32'hFFFF1170: romout <= 16'h41F9;
32'hFFFF1172: romout <= 16'hFFFF;
32'hFFFF1174: romout <= 16'h200C;
32'hFFFF1176: romout <= 16'h21C8;
32'hFFFF1178: romout <= 16'h000C;
32'hFFFF117A: romout <= 16'h41F9;
32'hFFFF117C: romout <= 16'hFFFF;
32'hFFFF117E: romout <= 16'h2038;
32'hFFFF1180: romout <= 16'h21C8;
32'hFFFF1182: romout <= 16'h0010;
32'hFFFF1184: romout <= 16'h41F9;
32'hFFFF1186: romout <= 16'hFFFF;
32'hFFFF1188: romout <= 16'h1298;
32'hFFFF118A: romout <= 16'h21C8;
32'hFFFF118C: romout <= 16'h0078;
32'hFFFF118E: romout <= 16'h41F9;
32'hFFFF1190: romout <= 16'hFFFF;
32'hFFFF1192: romout <= 16'h1250;
32'hFFFF1194: romout <= 16'h21C8;
32'hFFFF1196: romout <= 16'h007C;
32'hFFFF1198: romout <= 16'h41F9;
32'hFFFF119A: romout <= 16'hFFFF;
32'hFFFF119C: romout <= 16'h0800;
32'hFFFF119E: romout <= 16'h21C8;
32'hFFFF11A0: romout <= 16'h0080;
32'hFFFF11A2: romout <= 16'h41F9;
32'hFFFF11A4: romout <= 16'hFFFF;
32'hFFFF11A6: romout <= 16'h0400;
32'hFFFF11A8: romout <= 16'h21C8;
32'hFFFF11AA: romout <= 16'h0084;
32'hFFFF11AC: romout <= 16'h41F9;
32'hFFFF11AE: romout <= 16'hFFFF;
32'hFFFF11B0: romout <= 16'h0C00;
32'hFFFF11B2: romout <= 16'h21C8;
32'hFFFF11B4: romout <= 16'h0088;
32'hFFFF11B6: romout <= 16'h41F9;
32'hFFFF11B8: romout <= 16'hFFFF;
32'hFFFF11BA: romout <= 16'h1312;
32'hFFFF11BC: romout <= 16'h21C8;
32'hFFFF11BE: romout <= 16'h00BC;
32'hFFFF11C0: romout <= 16'h42B8;
32'hFFFF11C2: romout <= 16'h0400;
32'hFFFF11C4: romout <= 16'h027C;
32'hFFFF11C6: romout <= 16'hF000;
32'hFFFF11C8: romout <= 16'h700E;
32'hFFFF11CA: romout <= 16'h43F9;
32'hFFFF11CC: romout <= 16'hFFFF;
32'hFFFF11CE: romout <= 16'h1241;
32'hFFFF11D0: romout <= 16'h4E4F;
32'hFFFF11D2: romout <= 16'h4EF9;
32'hFFFF11D4: romout <= 16'hFFFF;
32'hFFFF11D6: romout <= 16'h2400;
32'hFFFF11D8: romout <= 16'h7005;
32'hFFFF11DA: romout <= 16'h4E4F;
32'hFFFF11DC: romout <= 16'h0C01;
32'hFFFF11DE: romout <= 16'h0078;
32'hFFFF11E0: romout <= 16'h66F0;
32'hFFFF11E2: romout <= 16'h203C;
32'hFFFF11E4: romout <= 16'h0004;
32'hFFFF11E6: romout <= 16'h0000;
32'hFFFF11E8: romout <= 16'h41F9;
32'hFFFF11EA: romout <= 16'h0002;
32'hFFFF11EC: romout <= 16'h0000;
32'hFFFF11EE: romout <= 16'h343C;
32'hFFFF11F0: romout <= 16'h1234;
32'hFFFF11F2: romout <= 16'h30C2;
32'hFFFF11F4: romout <= 16'h5380;
32'hFFFF11F6: romout <= 16'h66FA;
32'hFFFF11F8: romout <= 16'h4EF9;
32'hFFFF11FA: romout <= 16'hFFFF;
32'hFFFF11FC: romout <= 16'h2400;
32'hFFFF11FE: romout <= 16'h4239;
32'hFFFF1200: romout <= 16'hFFDC;
32'hFFFF1202: romout <= 16'h0A07;
32'hFFFF1204: romout <= 16'h45F9;
32'hFFFF1206: romout <= 16'hFFFF;
32'hFFFF1208: romout <= 16'h0000;
32'hFFFF120A: romout <= 16'h121A;
32'hFFFF120C: romout <= 16'h1039;
32'hFFFF120E: romout <= 16'hFFDC;
32'hFFFF1210: romout <= 16'h0A01;
32'hFFFF1212: romout <= 16'h0800;
32'hFFFF1214: romout <= 16'h0005;
32'hFFFF1216: romout <= 16'h67F4;
32'hFFFF1218: romout <= 16'h13C1;
32'hFFFF121A: romout <= 16'hFFDC;
32'hFFFF121C: romout <= 16'h0A00;
32'hFFFF121E: romout <= 16'hB5FC;
32'hFFFF1220: romout <= 16'hFFFF;
32'hFFFF1222: romout <= 16'h0100;
32'hFFFF1224: romout <= 16'h65E4;
32'hFFFF1226: romout <= 16'h60DC;
32'hFFFF1228: romout <= 16'h1039;
32'hFFFF122A: romout <= 16'hFFDD;
32'hFFFF122C: romout <= 16'h0000;
32'hFFFF122E: romout <= 16'h6AF8;
32'hFFFF1230: romout <= 16'h2079;
32'hFFFF1232: romout <= 16'hFFDD;
32'hFFFF1234: romout <= 16'h0004;
32'hFFFF1236: romout <= 16'h4ED0;
32'hFFFF1238: romout <= 16'h5241;
32'hFFFF123A: romout <= 16'h4D20;
32'hFFFF123C: romout <= 16'h5445;
32'hFFFF123E: romout <= 16'h5354;
32'hFFFF1240: romout <= 16'h0042;
32'hFFFF1242: romout <= 16'h4F4F;
32'hFFFF1244: romout <= 16'h5449;
32'hFFFF1246: romout <= 16'h4E47;
32'hFFFF1248: romout <= 16'h2E2E;
32'hFFFF124A: romout <= 16'h2E2E;
32'hFFFF124C: romout <= 16'h00FF;
32'hFFFF124E: romout <= 16'hFFFF;
32'hFFFF1250: romout <= 16'h4EF9;
32'hFFFF1252: romout <= 16'hFFFF;
32'hFFFF1254: romout <= 16'h1100;
32'hFFFF1256: romout <= 16'h4E73;
32'hFFFF1258: romout <= 16'h48E7;
32'hFFFF125A: romout <= 16'hC080;
32'hFFFF125C: romout <= 16'h3238;
32'hFFFF125E: romout <= 16'h0450;
32'hFFFF1260: romout <= 16'h0241;
32'hFFFF1262: romout <= 16'h000F;
32'hFFFF1264: romout <= 16'h41F8;
32'hFFFF1266: romout <= 16'h0440;
32'hFFFF1268: romout <= 16'h3039;
32'hFFFF126A: romout <= 16'hFFDC;
32'hFFFF126C: romout <= 16'h0000;
32'hFFFF126E: romout <= 16'h4279;
32'hFFFF1270: romout <= 16'hFFDC;
32'hFFFF1272: romout <= 16'h0002;
32'hFFFF1274: romout <= 16'h1180;
32'hFFFF1276: romout <= 16'h1000;
32'hFFFF1278: romout <= 16'h5241;
32'hFFFF127A: romout <= 16'h0241;
32'hFFFF127C: romout <= 16'h000F;
32'hFFFF127E: romout <= 16'h31C1;
32'hFFFF1280: romout <= 16'h0450;
32'hFFFF1282: romout <= 16'hB278;
32'hFFFF1284: romout <= 16'h0452;
32'hFFFF1286: romout <= 16'h660A;
32'hFFFF1288: romout <= 16'h5241;
32'hFFFF128A: romout <= 16'h0241;
32'hFFFF128C: romout <= 16'h000F;
32'hFFFF128E: romout <= 16'h31C1;
32'hFFFF1290: romout <= 16'h0452;
32'hFFFF1292: romout <= 16'h4CDF;
32'hFFFF1294: romout <= 16'h0103;
32'hFFFF1296: romout <= 16'h4E73;
32'hFFFF1298: romout <= 16'h2F00;
32'hFFFF129A: romout <= 16'h52B8;
32'hFFFF129C: romout <= 16'h0400;
32'hFFFF129E: romout <= 16'h5279;
32'hFFFF12A0: romout <= 16'hFFD0;
32'hFFFF12A2: romout <= 16'h0066;
32'hFFFF12A4: romout <= 16'h4A39;
32'hFFFF12A6: romout <= 16'hFFFF;
32'hFFFF12A8: romout <= 16'h0000;
32'hFFFF12AA: romout <= 16'h2038;
32'hFFFF12AC: romout <= 16'h0400;
32'hFFFF12AE: romout <= 16'h0200;
32'hFFFF12B0: romout <= 16'h007F;
32'hFFFF12B2: romout <= 16'h0C00;
32'hFFFF12B4: romout <= 16'h0040;
32'hFFFF12B6: romout <= 16'h6604;
32'hFFFF12B8: romout <= 16'h6100;
32'hFFFF12BA: romout <= 16'h0006;
32'hFFFF12BC: romout <= 16'h201F;
32'hFFFF12BE: romout <= 16'h4E73;
32'hFFFF12C0: romout <= 16'h48E7;
32'hFFFF12C2: romout <= 16'hA0C0;
32'hFFFF12C4: romout <= 16'h6100;
32'hFFFF12C6: romout <= 16'h0440;
32'hFFFF12C8: romout <= 16'hD1FC;
32'hFFFF12CA: romout <= 16'h0001;
32'hFFFF12CC: romout <= 16'h0000;
32'hFFFF12CE: romout <= 16'h3010;
32'hFFFF12D0: romout <= 16'hE818;
32'hFFFF12D2: romout <= 16'h3080;
32'hFFFF12D4: romout <= 16'hB1F8;
32'hFFFF12D6: romout <= 16'h0404;
32'hFFFF12D8: romout <= 16'h670C;
32'hFFFF12DA: romout <= 16'h2278;
32'hFFFF12DC: romout <= 16'h0404;
32'hFFFF12DE: romout <= 16'h32B8;
32'hFFFF12E0: romout <= 16'h0414;
32'hFFFF12E2: romout <= 16'h21C8;
32'hFFFF12E4: romout <= 16'h0404;
32'hFFFF12E6: romout <= 16'h4CDF;
32'hFFFF12E8: romout <= 16'h0305;
32'hFFFF12EA: romout <= 16'h4E75;
32'hFFFF12EC: romout <= 16'h4E55;
32'hFFFF12EE: romout <= 16'hFFE8;
32'hFFFF12F0: romout <= 16'h41ED;
32'hFFFF12F2: romout <= 16'hFFFA;
32'hFFFF12F4: romout <= 16'h43ED;
32'hFFFF12F6: romout <= 16'hFFFC;
32'hFFFF12F8: romout <= 16'h3B7C;
32'hFFFF12FA: romout <= 16'h0000;
32'hFFFF12FC: romout <= 16'hFFFA;
32'hFFFF12FE: romout <= 16'h3B7C;
32'hFFFF1300: romout <= 16'h0002;
32'hFFFF1302: romout <= 16'hFFF8;
32'hFFFF1304: romout <= 16'h7048;
32'hFFFF1306: romout <= 16'h4E41;
32'hFFFF1308: romout <= 16'h5279;
32'hFFFF130A: romout <= 16'hFFD0;
32'hFFFF130C: romout <= 16'h0064;
32'hFFFF130E: romout <= 16'h4E40;
32'hFFFF1310: romout <= 16'h60F6;
32'hFFFF1312: romout <= 16'h48E7;
32'hFFFF1314: romout <= 16'h8080;
32'hFFFF1316: romout <= 16'h41F9;
32'hFFFF1318: romout <= 16'hFFFF;
32'hFFFF131A: romout <= 16'h1330;
32'hFFFF131C: romout <= 16'h0280;
32'hFFFF131E: romout <= 16'h0000;
32'hFFFF1320: romout <= 16'h00FF;
32'hFFFF1322: romout <= 16'hE580;
32'hFFFF1324: romout <= 16'h2070;
32'hFFFF1326: romout <= 16'h0000;
32'hFFFF1328: romout <= 16'h4E90;
32'hFFFF132A: romout <= 16'h4CDF;
32'hFFFF132C: romout <= 16'h0101;
32'hFFFF132E: romout <= 16'h4E73;
32'hFFFF1330: romout <= 16'hFFFF;
32'hFFFF1332: romout <= 16'h189A;
32'hFFFF1334: romout <= 16'hFFFF;
32'hFFFF1336: romout <= 16'h187A;
32'hFFFF1338: romout <= 16'hFFFF;
32'hFFFF133A: romout <= 16'h149C;
32'hFFFF133C: romout <= 16'hFFFF;
32'hFFFF133E: romout <= 16'h19A0;
32'hFFFF1340: romout <= 16'hFFFF;
32'hFFFF1342: romout <= 16'h149C;
32'hFFFF1344: romout <= 16'hFFFF;
32'hFFFF1346: romout <= 16'h1658;
32'hFFFF1348: romout <= 16'hFFFF;
32'hFFFF134A: romout <= 16'h1732;
32'hFFFF134C: romout <= 16'hFFFF;
32'hFFFF134E: romout <= 16'h16DA;
32'hFFFF1350: romout <= 16'hFFFF;
32'hFFFF1352: romout <= 16'h149C;
32'hFFFF1354: romout <= 16'hFFFF;
32'hFFFF1356: romout <= 16'h149C;
32'hFFFF1358: romout <= 16'hFFFF;
32'hFFFF135A: romout <= 16'h149C;
32'hFFFF135C: romout <= 16'hFFFF;
32'hFFFF135E: romout <= 16'h18A2;
32'hFFFF1360: romout <= 16'hFFFF;
32'hFFFF1362: romout <= 16'h162C;
32'hFFFF1364: romout <= 16'hFFFF;
32'hFFFF1366: romout <= 16'h1872;
32'hFFFF1368: romout <= 16'hFFFF;
32'hFFFF136A: romout <= 16'h1858;
32'hFFFF136C: romout <= 16'hFFFF;
32'hFFFF136E: romout <= 16'h149C;
32'hFFFF1370: romout <= 16'hFFFF;
32'hFFFF1372: romout <= 16'h149C;
32'hFFFF1374: romout <= 16'hFFFF;
32'hFFFF1376: romout <= 16'h149C;
32'hFFFF1378: romout <= 16'hFFFF;
32'hFFFF137A: romout <= 16'h149C;
32'hFFFF137C: romout <= 16'hFFFF;
32'hFFFF137E: romout <= 16'h149C;
32'hFFFF1380: romout <= 16'hFFFF;
32'hFFFF1382: romout <= 16'h198C;
32'hFFFF1384: romout <= 16'hFFFF;
32'hFFFF1386: romout <= 16'h149C;
32'hFFFF1388: romout <= 16'hFFFF;
32'hFFFF138A: romout <= 16'h149C;
32'hFFFF138C: romout <= 16'hFFFF;
32'hFFFF138E: romout <= 16'h149C;
32'hFFFF1390: romout <= 16'hFFFF;
32'hFFFF1392: romout <= 16'h149C;
32'hFFFF1394: romout <= 16'hFFFF;
32'hFFFF1396: romout <= 16'h149C;
32'hFFFF1398: romout <= 16'hFFFF;
32'hFFFF139A: romout <= 16'h149C;
32'hFFFF139C: romout <= 16'hFFFF;
32'hFFFF139E: romout <= 16'h149C;
32'hFFFF13A0: romout <= 16'hFFFF;
32'hFFFF13A2: romout <= 16'h149C;
32'hFFFF13A4: romout <= 16'hFFFF;
32'hFFFF13A6: romout <= 16'h149C;
32'hFFFF13A8: romout <= 16'hFFFF;
32'hFFFF13AA: romout <= 16'h149C;
32'hFFFF13AC: romout <= 16'hFFFF;
32'hFFFF13AE: romout <= 16'h149C;
32'hFFFF13B0: romout <= 16'hFFFF;
32'hFFFF13B2: romout <= 16'h149C;
32'hFFFF13B4: romout <= 16'hFFFF;
32'hFFFF13B6: romout <= 16'h149C;
32'hFFFF13B8: romout <= 16'hFFFF;
32'hFFFF13BA: romout <= 16'h149C;
32'hFFFF13BC: romout <= 16'hFFFF;
32'hFFFF13BE: romout <= 16'h149C;
32'hFFFF13C0: romout <= 16'hFFFF;
32'hFFFF13C2: romout <= 16'h149C;
32'hFFFF13C4: romout <= 16'hFFFF;
32'hFFFF13C6: romout <= 16'h149C;
32'hFFFF13C8: romout <= 16'hFFFF;
32'hFFFF13CA: romout <= 16'h149C;
32'hFFFF13CC: romout <= 16'hFFFF;
32'hFFFF13CE: romout <= 16'h149C;
32'hFFFF13D0: romout <= 16'hFFFF;
32'hFFFF13D2: romout <= 16'h149C;
32'hFFFF13D4: romout <= 16'hFFFF;
32'hFFFF13D6: romout <= 16'h149C;
32'hFFFF13D8: romout <= 16'hFFFF;
32'hFFFF13DA: romout <= 16'h149C;
32'hFFFF13DC: romout <= 16'hFFFF;
32'hFFFF13DE: romout <= 16'h149C;
32'hFFFF13E0: romout <= 16'hFFFF;
32'hFFFF13E2: romout <= 16'h149C;
32'hFFFF13E4: romout <= 16'hFFFF;
32'hFFFF13E6: romout <= 16'h149C;
32'hFFFF13E8: romout <= 16'hFFFF;
32'hFFFF13EA: romout <= 16'h149C;
32'hFFFF13EC: romout <= 16'hFFFF;
32'hFFFF13EE: romout <= 16'h149C;
32'hFFFF13F0: romout <= 16'hFFFF;
32'hFFFF13F2: romout <= 16'h149C;
32'hFFFF13F4: romout <= 16'hFFFF;
32'hFFFF13F6: romout <= 16'h149C;
32'hFFFF13F8: romout <= 16'hFFFF;
32'hFFFF13FA: romout <= 16'h149C;
32'hFFFF13FC: romout <= 16'hFFFF;
32'hFFFF13FE: romout <= 16'h149C;
32'hFFFF1400: romout <= 16'hFFFF;
32'hFFFF1402: romout <= 16'h149C;
32'hFFFF1404: romout <= 16'hFFFF;
32'hFFFF1406: romout <= 16'h149C;
32'hFFFF1408: romout <= 16'hFFFF;
32'hFFFF140A: romout <= 16'h149C;
32'hFFFF140C: romout <= 16'hFFFF;
32'hFFFF140E: romout <= 16'h149C;
32'hFFFF1410: romout <= 16'hFFFF;
32'hFFFF1412: romout <= 16'h149C;
32'hFFFF1414: romout <= 16'hFFFF;
32'hFFFF1416: romout <= 16'h149C;
32'hFFFF1418: romout <= 16'hFFFF;
32'hFFFF141A: romout <= 16'h149C;
32'hFFFF141C: romout <= 16'hFFFF;
32'hFFFF141E: romout <= 16'h149C;
32'hFFFF1420: romout <= 16'hFFFF;
32'hFFFF1422: romout <= 16'h149C;
32'hFFFF1424: romout <= 16'hFFFF;
32'hFFFF1426: romout <= 16'h149C;
32'hFFFF1428: romout <= 16'hFFFF;
32'hFFFF142A: romout <= 16'h149C;
32'hFFFF142C: romout <= 16'hFFFF;
32'hFFFF142E: romout <= 16'h149C;
32'hFFFF1430: romout <= 16'hFFFF;
32'hFFFF1432: romout <= 16'h149C;
32'hFFFF1434: romout <= 16'hFFFF;
32'hFFFF1436: romout <= 16'h149C;
32'hFFFF1438: romout <= 16'hFFFF;
32'hFFFF143A: romout <= 16'h149C;
32'hFFFF143C: romout <= 16'hFFFF;
32'hFFFF143E: romout <= 16'h149C;
32'hFFFF1440: romout <= 16'hFFFF;
32'hFFFF1442: romout <= 16'h149C;
32'hFFFF1444: romout <= 16'hFFFF;
32'hFFFF1446: romout <= 16'h149C;
32'hFFFF1448: romout <= 16'hFFFF;
32'hFFFF144A: romout <= 16'h149C;
32'hFFFF144C: romout <= 16'hFFFF;
32'hFFFF144E: romout <= 16'h149C;
32'hFFFF1450: romout <= 16'hFFFF;
32'hFFFF1452: romout <= 16'h149C;
32'hFFFF1454: romout <= 16'hFFFF;
32'hFFFF1456: romout <= 16'h149C;
32'hFFFF1458: romout <= 16'hFFFF;
32'hFFFF145A: romout <= 16'h149C;
32'hFFFF145C: romout <= 16'hFFFF;
32'hFFFF145E: romout <= 16'h149C;
32'hFFFF1460: romout <= 16'hFFFF;
32'hFFFF1462: romout <= 16'h149C;
32'hFFFF1464: romout <= 16'hFFFF;
32'hFFFF1466: romout <= 16'h149C;
32'hFFFF1468: romout <= 16'hFFFF;
32'hFFFF146A: romout <= 16'h149C;
32'hFFFF146C: romout <= 16'hFFFF;
32'hFFFF146E: romout <= 16'h149C;
32'hFFFF1470: romout <= 16'hFFFF;
32'hFFFF1472: romout <= 16'h149E;
32'hFFFF1474: romout <= 16'hFFFF;
32'hFFFF1476: romout <= 16'h14B4;
32'hFFFF1478: romout <= 16'hFFFF;
32'hFFFF147A: romout <= 16'h14FE;
32'hFFFF147C: romout <= 16'hFFFF;
32'hFFFF147E: romout <= 16'h149C;
32'hFFFF1480: romout <= 16'hFFFF;
32'hFFFF1482: romout <= 16'h1528;
32'hFFFF1484: romout <= 16'hFFFF;
32'hFFFF1486: romout <= 16'h159A;
32'hFFFF1488: romout <= 16'hFFFF;
32'hFFFF148A: romout <= 16'h15B4;
32'hFFFF148C: romout <= 16'hFFFF;
32'hFFFF148E: romout <= 16'h15FA;
32'hFFFF1490: romout <= 16'hFFFF;
32'hFFFF1492: romout <= 16'h149C;
32'hFFFF1494: romout <= 16'hFFFF;
32'hFFFF1496: romout <= 16'h149C;
32'hFFFF1498: romout <= 16'hFFFF;
32'hFFFF149A: romout <= 16'h15BE;
32'hFFFF149C: romout <= 16'h4E75;
32'hFFFF149E: romout <= 16'h48E7;
32'hFFFF14A0: romout <= 16'hC000;
32'hFFFF14A2: romout <= 16'h21C1;
32'hFFFF14A4: romout <= 16'h0420;
32'hFFFF14A6: romout <= 16'h6100;
32'hFFFF14A8: romout <= 16'h0022;
32'hFFFF14AA: romout <= 16'h11C1;
32'hFFFF14AC: romout <= 16'h0424;
32'hFFFF14AE: romout <= 16'h4CDF;
32'hFFFF14B0: romout <= 16'h0003;
32'hFFFF14B2: romout <= 16'h4E75;
32'hFFFF14B4: romout <= 16'h48E7;
32'hFFFF14B6: romout <= 16'hC000;
32'hFFFF14B8: romout <= 16'h21C1;
32'hFFFF14BA: romout <= 16'h0428;
32'hFFFF14BC: romout <= 16'h6100;
32'hFFFF14BE: romout <= 16'h000C;
32'hFFFF14C0: romout <= 16'h11C1;
32'hFFFF14C2: romout <= 16'h042C;
32'hFFFF14C4: romout <= 16'h4CDF;
32'hFFFF14C6: romout <= 16'h0003;
32'hFFFF14C8: romout <= 16'h4E75;
32'hFFFF14CA: romout <= 16'h48E7;
32'hFFFF14CC: romout <= 16'hA000;
32'hFFFF14CE: romout <= 16'h4282;
32'hFFFF14D0: romout <= 16'hEC99;
32'hFFFF14D2: romout <= 16'h2001;
32'hFFFF14D4: romout <= 16'h0200;
32'hFFFF14D6: romout <= 16'h0003;
32'hFFFF14D8: romout <= 16'h1400;
32'hFFFF14DA: romout <= 16'hE499;
32'hFFFF14DC: romout <= 16'hEA99;
32'hFFFF14DE: romout <= 16'h1001;
32'hFFFF14E0: romout <= 16'h0200;
32'hFFFF14E2: romout <= 16'h0007;
32'hFFFF14E4: romout <= 16'hE540;
32'hFFFF14E6: romout <= 16'h8400;
32'hFFFF14E8: romout <= 16'hE699;
32'hFFFF14EA: romout <= 16'hEA99;
32'hFFFF14EC: romout <= 16'h1001;
32'hFFFF14EE: romout <= 16'h0200;
32'hFFFF14F0: romout <= 16'h0007;
32'hFFFF14F2: romout <= 16'hEB40;
32'hFFFF14F4: romout <= 16'h8400;
32'hFFFF14F6: romout <= 16'h2202;
32'hFFFF14F8: romout <= 16'h4CDF;
32'hFFFF14FA: romout <= 16'h0005;
32'hFFFF14FC: romout <= 16'h4E75;
32'hFFFF14FE: romout <= 16'h48E7;
32'hFFFF1500: romout <= 16'h6080;
32'hFFFF1502: romout <= 16'hC4FC;
32'hFFFF1504: romout <= 16'h00D0;
32'hFFFF1506: romout <= 16'h0282;
32'hFFFF1508: romout <= 16'h0000;
32'hFFFF150A: romout <= 16'hFFFF;
32'hFFFF150C: romout <= 16'hE382;
32'hFFFF150E: romout <= 16'h0281;
32'hFFFF1510: romout <= 16'h0000;
32'hFFFF1512: romout <= 16'h01FF;
32'hFFFF1514: romout <= 16'hD481;
32'hFFFF1516: romout <= 16'h0682;
32'hFFFF1518: romout <= 16'h0002;
32'hFFFF151A: romout <= 16'h0000;
32'hFFFF151C: romout <= 16'h2042;
32'hFFFF151E: romout <= 16'h10B8;
32'hFFFF1520: romout <= 16'h0424;
32'hFFFF1522: romout <= 16'h4CDF;
32'hFFFF1524: romout <= 16'h0106;
32'hFFFF1526: romout <= 16'h4E75;
32'hFFFF1528: romout <= 16'h48E7;
32'hFFFF152A: romout <= 16'hFF30;
32'hFFFF152C: romout <= 16'h0281;
32'hFFFF152E: romout <= 16'h0000;
32'hFFFF1530: romout <= 16'h01FF;
32'hFFFF1532: romout <= 16'h0282;
32'hFFFF1534: romout <= 16'h0000;
32'hFFFF1536: romout <= 16'h01FF;
32'hFFFF1538: romout <= 16'h0283;
32'hFFFF153A: romout <= 16'h0000;
32'hFFFF153C: romout <= 16'h01FF;
32'hFFFF153E: romout <= 16'h0284;
32'hFFFF1540: romout <= 16'h0000;
32'hFFFF1542: romout <= 16'h01FF;
32'hFFFF1544: romout <= 16'h31C3;
32'hFFFF1546: romout <= 16'h0430;
32'hFFFF1548: romout <= 16'h31C4;
32'hFFFF154A: romout <= 16'h0432;
32'hFFFF154C: romout <= 16'h2A01;
32'hFFFF154E: romout <= 16'h9A83;
32'hFFFF1550: romout <= 16'h6A02;
32'hFFFF1552: romout <= 16'h4485;
32'hFFFF1554: romout <= 16'h2C02;
32'hFFFF1556: romout <= 16'h9C84;
32'hFFFF1558: romout <= 16'h6A02;
32'hFFFF155A: romout <= 16'h4486;
32'hFFFF155C: romout <= 16'h7001;
32'hFFFF155E: romout <= 16'h7E01;
32'hFFFF1560: romout <= 16'hB283;
32'hFFFF1562: romout <= 16'h6502;
32'hFFFF1564: romout <= 16'h4480;
32'hFFFF1566: romout <= 16'hB484;
32'hFFFF1568: romout <= 16'h6502;
32'hFFFF156A: romout <= 16'h4487;
32'hFFFF156C: romout <= 16'h2445;
32'hFFFF156E: romout <= 16'h95C6;
32'hFFFF1570: romout <= 16'h4486;
32'hFFFF1572: romout <= 16'h6100;
32'hFFFF1574: romout <= 16'hFF8A;
32'hFFFF1576: romout <= 16'hB681;
32'hFFFF1578: romout <= 16'h6604;
32'hFFFF157A: romout <= 16'hB882;
32'hFFFF157C: romout <= 16'h6716;
32'hFFFF157E: romout <= 16'h264A;
32'hFFFF1580: romout <= 16'hD7CB;
32'hFFFF1582: romout <= 16'hB7C6;
32'hFFFF1584: romout <= 16'h6F04;
32'hFFFF1586: romout <= 16'hD5C6;
32'hFFFF1588: romout <= 16'hD280;
32'hFFFF158A: romout <= 16'hB7C5;
32'hFFFF158C: romout <= 16'h6C04;
32'hFFFF158E: romout <= 16'hD5C5;
32'hFFFF1590: romout <= 16'hD487;
32'hFFFF1592: romout <= 16'h60DE;
32'hFFFF1594: romout <= 16'h4CDF;
32'hFFFF1596: romout <= 16'h0CFF;
32'hFFFF1598: romout <= 16'h4E75;
32'hFFFF159A: romout <= 16'h48E7;
32'hFFFF159C: romout <= 16'h7800;
32'hFFFF159E: romout <= 16'h3601;
32'hFFFF15A0: romout <= 16'h3802;
32'hFFFF15A2: romout <= 16'h3238;
32'hFFFF15A4: romout <= 16'h0430;
32'hFFFF15A6: romout <= 16'h3438;
32'hFFFF15A8: romout <= 16'h0432;
32'hFFFF15AA: romout <= 16'h6100;
32'hFFFF15AC: romout <= 16'hFF7C;
32'hFFFF15AE: romout <= 16'h4CDF;
32'hFFFF15B0: romout <= 16'h001E;
32'hFFFF15B2: romout <= 16'h4E75;
32'hFFFF15B4: romout <= 16'h31C1;
32'hFFFF15B6: romout <= 16'h0430;
32'hFFFF15B8: romout <= 16'h31C2;
32'hFFFF15BA: romout <= 16'h0432;
32'hFFFF15BC: romout <= 16'h4E75;
32'hFFFF15BE: romout <= 16'h48E7;
32'hFFFF15C0: romout <= 16'hFF00;
32'hFFFF15C2: romout <= 16'h3001;
32'hFFFF15C4: romout <= 16'h3E02;
32'hFFFF15C6: romout <= 16'h3A03;
32'hFFFF15C8: romout <= 16'h3C04;
32'hFFFF15CA: romout <= 16'h3802;
32'hFFFF15CC: romout <= 16'h6100;
32'hFFFF15CE: romout <= 16'hFF5A;
32'hFFFF15D0: romout <= 16'h3203;
32'hFFFF15D2: romout <= 16'h3404;
32'hFFFF15D4: romout <= 16'h3605;
32'hFFFF15D6: romout <= 16'h3806;
32'hFFFF15D8: romout <= 16'h6100;
32'hFFFF15DA: romout <= 16'hFF4E;
32'hFFFF15DC: romout <= 16'h3203;
32'hFFFF15DE: romout <= 16'h3404;
32'hFFFF15E0: romout <= 16'h3600;
32'hFFFF15E2: romout <= 16'h3806;
32'hFFFF15E4: romout <= 16'h6100;
32'hFFFF15E6: romout <= 16'hFF42;
32'hFFFF15E8: romout <= 16'h3203;
32'hFFFF15EA: romout <= 16'h3404;
32'hFFFF15EC: romout <= 16'h3600;
32'hFFFF15EE: romout <= 16'h3807;
32'hFFFF15F0: romout <= 16'h6100;
32'hFFFF15F2: romout <= 16'hFF36;
32'hFFFF15F4: romout <= 16'h4CDF;
32'hFFFF15F6: romout <= 16'h00FF;
32'hFFFF15F8: romout <= 16'h4E75;
32'hFFFF15FA: romout <= 16'h48E7;
32'hFFFF15FC: romout <= 16'h7800;
32'hFFFF15FE: romout <= 16'h3F38;
32'hFFFF1600: romout <= 16'h0424;
32'hFFFF1602: romout <= 16'h6100;
32'hFFFF1604: romout <= 16'hFFBA;
32'hFFFF1606: romout <= 16'h31F8;
32'hFFFF1608: romout <= 16'h042C;
32'hFFFF160A: romout <= 16'h0424;
32'hFFFF160C: romout <= 16'hB641;
32'hFFFF160E: romout <= 16'h6504;
32'hFFFF1610: romout <= 16'hB842;
32'hFFFF1612: romout <= 16'h640E;
32'hFFFF1614: romout <= 16'h5241;
32'hFFFF1616: romout <= 16'h5242;
32'hFFFF1618: romout <= 16'h5343;
32'hFFFF161A: romout <= 16'h5344;
32'hFFFF161C: romout <= 16'h6100;
32'hFFFF161E: romout <= 16'hFFA0;
32'hFFFF1620: romout <= 16'h60EA;
32'hFFFF1622: romout <= 16'h31DF;
32'hFFFF1624: romout <= 16'h0424;
32'hFFFF1626: romout <= 16'h4CDF;
32'hFFFF1628: romout <= 16'h001E;
32'hFFFF162A: romout <= 16'h4E75;
32'hFFFF162C: romout <= 16'h11C1;
32'hFFFF162E: romout <= 16'h041C;
32'hFFFF1630: romout <= 16'h4E75;
32'hFFFF1632: romout <= 16'h4E71;
32'hFFFF1634: romout <= 16'h4E71;
32'hFFFF1636: romout <= 16'h4E71;
32'hFFFF1638: romout <= 16'h4E71;
32'hFFFF163A: romout <= 16'h4E71;
32'hFFFF163C: romout <= 16'h4E71;
32'hFFFF163E: romout <= 16'h4E71;
32'hFFFF1640: romout <= 16'h4E71;
32'hFFFF1642: romout <= 16'h4E71;
32'hFFFF1644: romout <= 16'h4E71;
32'hFFFF1646: romout <= 16'h4E71;
32'hFFFF1648: romout <= 16'h4E71;
32'hFFFF164A: romout <= 16'h4E71;
32'hFFFF164C: romout <= 16'h4E71;
32'hFFFF164E: romout <= 16'h4E71;
32'hFFFF1650: romout <= 16'h4E71;
32'hFFFF1652: romout <= 16'h4E71;
32'hFFFF1654: romout <= 16'h4E71;
32'hFFFF1656: romout <= 16'h4E71;
32'hFFFF1658: romout <= 16'h3239;
32'hFFFF165A: romout <= 16'hFFDC;
32'hFFFF165C: romout <= 16'h0000;
32'hFFFF165E: romout <= 16'h6AF8;
32'hFFFF1660: romout <= 16'h4279;
32'hFFFF1662: romout <= 16'hFFDC;
32'hFFFF1664: romout <= 16'h0002;
32'hFFFF1666: romout <= 16'h0241;
32'hFFFF1668: romout <= 16'h00FF;
32'hFFFF166A: romout <= 16'h0C38;
32'hFFFF166C: romout <= 16'h0000;
32'hFFFF166E: romout <= 16'h041C;
32'hFFFF1670: romout <= 16'h670C;
32'hFFFF1672: romout <= 16'h0C01;
32'hFFFF1674: romout <= 16'h000D;
32'hFFFF1676: romout <= 16'h6774;
32'hFFFF1678: romout <= 16'h4EB9;
32'hFFFF167A: romout <= 16'hFFFF;
32'hFFFF167C: romout <= 16'h1732;
32'hFFFF167E: romout <= 16'h4E75;
32'hFFFF1680: romout <= 16'h3F01;
32'hFFFF1682: romout <= 16'h3239;
32'hFFFF1684: romout <= 16'hFFDC;
32'hFFFF1686: romout <= 16'h0000;
32'hFFFF1688: romout <= 16'h6A08;
32'hFFFF168A: romout <= 16'h321F;
32'hFFFF168C: romout <= 16'h003C;
32'hFFFF168E: romout <= 16'h0001;
32'hFFFF1690: romout <= 16'h4E75;
32'hFFFF1692: romout <= 16'h321F;
32'hFFFF1694: romout <= 16'h023C;
32'hFFFF1696: romout <= 16'h00FE;
32'hFFFF1698: romout <= 16'h4E75;
32'hFFFF169A: romout <= 16'h0839;
32'hFFFF169C: romout <= 16'h0000;
32'hFFFF169E: romout <= 16'hFFDC;
32'hFFFF16A0: romout <= 16'h0A01;
32'hFFFF16A2: romout <= 16'h6706;
32'hFFFF16A4: romout <= 16'h003C;
32'hFFFF16A6: romout <= 16'h0001;
32'hFFFF16A8: romout <= 16'h4E75;
32'hFFFF16AA: romout <= 16'h023C;
32'hFFFF16AC: romout <= 16'h00FE;
32'hFFFF16AE: romout <= 16'h4E75;
32'hFFFF16B0: romout <= 16'h4280;
32'hFFFF16B2: romout <= 16'h3039;
32'hFFFF16B4: romout <= 16'hFFDC;
32'hFFFF16B6: romout <= 16'h0000;
32'hFFFF16B8: romout <= 16'h6A12;
32'hFFFF16BA: romout <= 16'h0240;
32'hFFFF16BC: romout <= 16'h00FF;
32'hFFFF16BE: romout <= 16'h4279;
32'hFFFF16C0: romout <= 16'hFFDC;
32'hFFFF16C2: romout <= 16'h0002;
32'hFFFF16C4: romout <= 16'h41F8;
32'hFFFF16C6: romout <= 16'h0460;
32'hFFFF16C8: romout <= 16'h2080;
32'hFFFF16CA: romout <= 16'h4E75;
32'hFFFF16CC: romout <= 16'h41F8;
32'hFFFF16CE: romout <= 16'h0460;
32'hFFFF16D0: romout <= 16'h4290;
32'hFFFF16D2: romout <= 16'h4E75;
32'hFFFF16D4: romout <= 16'h6100;
32'hFFFF16D6: romout <= 16'h005C;
32'hFFFF16D8: romout <= 16'h4E75;
32'hFFFF16DA: romout <= 16'h3239;
32'hFFFF16DC: romout <= 16'hFFDC;
32'hFFFF16DE: romout <= 16'h0000;
32'hFFFF16E0: romout <= 16'h6A06;
32'hFFFF16E2: romout <= 16'h123C;
32'hFFFF16E4: romout <= 16'h0001;
32'hFFFF16E6: romout <= 16'h4E75;
32'hFFFF16E8: romout <= 16'h4201;
32'hFFFF16EA: romout <= 16'h4E75;
32'hFFFF16EC: romout <= 16'h2F01;
32'hFFFF16EE: romout <= 16'h123C;
32'hFFFF16F0: romout <= 16'h000D;
32'hFFFF16F2: romout <= 16'h4EB9;
32'hFFFF16F4: romout <= 16'hFFFF;
32'hFFFF16F6: romout <= 16'h1732;
32'hFFFF16F8: romout <= 16'h123C;
32'hFFFF16FA: romout <= 16'h000A;
32'hFFFF16FC: romout <= 16'h4EB9;
32'hFFFF16FE: romout <= 16'hFFFF;
32'hFFFF1700: romout <= 16'h1732;
32'hFFFF1702: romout <= 16'h221F;
32'hFFFF1704: romout <= 16'h4E75;
32'hFFFF1706: romout <= 16'h3038;
32'hFFFF1708: romout <= 16'h0418;
32'hFFFF170A: romout <= 16'h0240;
32'hFFFF170C: romout <= 16'h007F;
32'hFFFF170E: romout <= 16'hC0F9;
32'hFFFF1710: romout <= 16'hFFDA;
32'hFFFF1712: romout <= 16'h0000;
32'hFFFF1714: romout <= 16'h3438;
32'hFFFF1716: romout <= 16'h041A;
32'hFFFF1718: romout <= 16'h0242;
32'hFFFF171A: romout <= 16'h00FF;
32'hFFFF171C: romout <= 16'hD042;
32'hFFFF171E: romout <= 16'hE340;
32'hFFFF1720: romout <= 16'h0680;
32'hFFFF1722: romout <= 16'hFFD0;
32'hFFFF1724: romout <= 16'h0000;
32'hFFFF1726: romout <= 16'h2040;
32'hFFFF1728: romout <= 16'hE288;
32'hFFFF172A: romout <= 16'h33C0;
32'hFFFF172C: romout <= 16'hFFDA;
32'hFFFF172E: romout <= 16'h0016;
32'hFFFF1730: romout <= 16'h4E75;
32'hFFFF1732: romout <= 16'h0C01;
32'hFFFF1734: romout <= 16'h000D;
32'hFFFF1736: romout <= 16'h6606;
32'hFFFF1738: romout <= 16'h4278;
32'hFFFF173A: romout <= 16'h041A;
32'hFFFF173C: romout <= 16'h4E75;
32'hFFFF173E: romout <= 16'h0C01;
32'hFFFF1740: romout <= 16'h0091;
32'hFFFF1742: romout <= 16'h660E;
32'hFFFF1744: romout <= 16'h0C78;
32'hFFFF1746: romout <= 16'h0033;
32'hFFFF1748: romout <= 16'h041A;
32'hFFFF174A: romout <= 16'h6704;
32'hFFFF174C: romout <= 16'h5278;
32'hFFFF174E: romout <= 16'h041A;
32'hFFFF1750: romout <= 16'h4E75;
32'hFFFF1752: romout <= 16'h0C01;
32'hFFFF1754: romout <= 16'h0090;
32'hFFFF1756: romout <= 16'h660E;
32'hFFFF1758: romout <= 16'h0C78;
32'hFFFF175A: romout <= 16'h0000;
32'hFFFF175C: romout <= 16'h0418;
32'hFFFF175E: romout <= 16'h67F0;
32'hFFFF1760: romout <= 16'h5378;
32'hFFFF1762: romout <= 16'h0418;
32'hFFFF1764: romout <= 16'h4E75;
32'hFFFF1766: romout <= 16'h0C01;
32'hFFFF1768: romout <= 16'h0093;
32'hFFFF176A: romout <= 16'h660E;
32'hFFFF176C: romout <= 16'h0C78;
32'hFFFF176E: romout <= 16'h0000;
32'hFFFF1770: romout <= 16'h041A;
32'hFFFF1772: romout <= 16'h67DC;
32'hFFFF1774: romout <= 16'h5378;
32'hFFFF1776: romout <= 16'h041A;
32'hFFFF1778: romout <= 16'h4E75;
32'hFFFF177A: romout <= 16'h0C01;
32'hFFFF177C: romout <= 16'h0092;
32'hFFFF177E: romout <= 16'h660E;
32'hFFFF1780: romout <= 16'h0C78;
32'hFFFF1782: romout <= 16'h001E;
32'hFFFF1784: romout <= 16'h0418;
32'hFFFF1786: romout <= 16'h67C8;
32'hFFFF1788: romout <= 16'h5278;
32'hFFFF178A: romout <= 16'h0418;
32'hFFFF178C: romout <= 16'h4E75;
32'hFFFF178E: romout <= 16'h0C01;
32'hFFFF1790: romout <= 16'h0094;
32'hFFFF1792: romout <= 16'h6614;
32'hFFFF1794: romout <= 16'h0C78;
32'hFFFF1796: romout <= 16'h0000;
32'hFFFF1798: romout <= 16'h041A;
32'hFFFF179A: romout <= 16'h6706;
32'hFFFF179C: romout <= 16'h4278;
32'hFFFF179E: romout <= 16'h041A;
32'hFFFF17A0: romout <= 16'h4E75;
32'hFFFF17A2: romout <= 16'h4278;
32'hFFFF17A4: romout <= 16'h0418;
32'hFFFF17A6: romout <= 16'h4E75;
32'hFFFF17A8: romout <= 16'h48E7;
32'hFFFF17AA: romout <= 16'hE080;
32'hFFFF17AC: romout <= 16'h0C01;
32'hFFFF17AE: romout <= 16'h0099;
32'hFFFF17B0: romout <= 16'h660A;
32'hFFFF17B2: romout <= 16'h6100;
32'hFFFF17B4: romout <= 16'hFF52;
32'hFFFF17B6: romout <= 16'h3038;
32'hFFFF17B8: romout <= 16'h041A;
32'hFFFF17BA: romout <= 16'h601A;
32'hFFFF17BC: romout <= 16'h0C01;
32'hFFFF17BE: romout <= 16'h0008;
32'hFFFF17C0: romout <= 16'h662C;
32'hFFFF17C2: romout <= 16'h0C78;
32'hFFFF17C4: romout <= 16'h0000;
32'hFFFF17C6: romout <= 16'h041A;
32'hFFFF17C8: romout <= 16'h6742;
32'hFFFF17CA: romout <= 16'h5378;
32'hFFFF17CC: romout <= 16'h041A;
32'hFFFF17CE: romout <= 16'h6100;
32'hFFFF17D0: romout <= 16'hFF36;
32'hFFFF17D2: romout <= 16'h3038;
32'hFFFF17D4: romout <= 16'h041A;
32'hFFFF17D6: romout <= 16'h30E8;
32'hFFFF17D8: romout <= 16'h0002;
32'hFFFF17DA: romout <= 16'h5240;
32'hFFFF17DC: romout <= 16'hB079;
32'hFFFF17DE: romout <= 16'hFFDA;
32'hFFFF17E0: romout <= 16'h0000;
32'hFFFF17E2: romout <= 16'h65F2;
32'hFFFF17E4: romout <= 16'h303C;
32'hFFFF17E6: romout <= 16'h0020;
32'hFFFF17E8: romout <= 16'h3140;
32'hFFFF17EA: romout <= 16'hFFFE;
32'hFFFF17EC: romout <= 16'h601E;
32'hFFFF17EE: romout <= 16'h0C01;
32'hFFFF17F0: romout <= 16'h000A;
32'hFFFF17F2: romout <= 16'h6714;
32'hFFFF17F4: romout <= 16'h6100;
32'hFFFF17F6: romout <= 16'hFF10;
32'hFFFF17F8: romout <= 16'h6100;
32'hFFFF17FA: romout <= 16'h01B8;
32'hFFFF17FC: romout <= 16'h30C1;
32'hFFFF17FE: romout <= 16'h6100;
32'hFFFF1800: romout <= 16'h0012;
32'hFFFF1802: romout <= 16'h4CDF;
32'hFFFF1804: romout <= 16'h0107;
32'hFFFF1806: romout <= 16'h4E75;
32'hFFFF1808: romout <= 16'h6100;
32'hFFFF180A: romout <= 16'h0022;
32'hFFFF180C: romout <= 16'h4CDF;
32'hFFFF180E: romout <= 16'h0107;
32'hFFFF1810: romout <= 16'h4E75;
32'hFFFF1812: romout <= 16'h5279;
32'hFFFF1814: romout <= 16'hFFDA;
32'hFFFF1816: romout <= 16'h0016;
32'hFFFF1818: romout <= 16'h5278;
32'hFFFF181A: romout <= 16'h041A;
32'hFFFF181C: romout <= 16'h3039;
32'hFFFF181E: romout <= 16'hFFDA;
32'hFFFF1820: romout <= 16'h0000;
32'hFFFF1822: romout <= 16'hB078;
32'hFFFF1824: romout <= 16'h041A;
32'hFFFF1826: romout <= 16'h642E;
32'hFFFF1828: romout <= 16'h4278;
32'hFFFF182A: romout <= 16'h041A;
32'hFFFF182C: romout <= 16'h5278;
32'hFFFF182E: romout <= 16'h0418;
32'hFFFF1830: romout <= 16'h3039;
32'hFFFF1832: romout <= 16'hFFDA;
32'hFFFF1834: romout <= 16'h0002;
32'hFFFF1836: romout <= 16'hB078;
32'hFFFF1838: romout <= 16'h0418;
32'hFFFF183A: romout <= 16'h621A;
32'hFFFF183C: romout <= 16'h3039;
32'hFFFF183E: romout <= 16'hFFDA;
32'hFFFF1840: romout <= 16'h0002;
32'hFFFF1842: romout <= 16'h31C0;
32'hFFFF1844: romout <= 16'h0418;
32'hFFFF1846: romout <= 16'h5378;
32'hFFFF1848: romout <= 16'h0418;
32'hFFFF184A: romout <= 16'hE340;
32'hFFFF184C: romout <= 16'h9179;
32'hFFFF184E: romout <= 16'hFFDA;
32'hFFFF1850: romout <= 16'h0016;
32'hFFFF1852: romout <= 16'h6100;
32'hFFFF1854: romout <= 16'h00CE;
32'hFFFF1856: romout <= 16'h4E75;
32'hFFFF1858: romout <= 16'h48E7;
32'hFFFF185A: romout <= 16'hC040;
32'hFFFF185C: romout <= 16'h4281;
32'hFFFF185E: romout <= 16'h1219;
32'hFFFF1860: romout <= 16'h0C01;
32'hFFFF1862: romout <= 16'h0000;
32'hFFFF1864: romout <= 16'h6706;
32'hFFFF1866: romout <= 16'h6100;
32'hFFFF1868: romout <= 16'hFECA;
32'hFFFF186A: romout <= 16'h60F0;
32'hFFFF186C: romout <= 16'h4CDF;
32'hFFFF186E: romout <= 16'h0203;
32'hFFFF1870: romout <= 16'h4E75;
32'hFFFF1872: romout <= 16'h6100;
32'hFFFF1874: romout <= 16'hFFE4;
32'hFFFF1876: romout <= 16'h6000;
32'hFFFF1878: romout <= 16'hFE74;
32'hFFFF187A: romout <= 16'h48E7;
32'hFFFF187C: romout <= 16'hC040;
32'hFFFF187E: romout <= 16'h0241;
32'hFFFF1880: romout <= 16'h00FF;
32'hFFFF1882: romout <= 16'h2001;
32'hFFFF1884: romout <= 16'h1219;
32'hFFFF1886: romout <= 16'h0C01;
32'hFFFF1888: romout <= 16'h0000;
32'hFFFF188A: romout <= 16'h6708;
32'hFFFF188C: romout <= 16'h6100;
32'hFFFF188E: romout <= 16'hFEA4;
32'hFFFF1890: romout <= 16'h57C8;
32'hFFFF1892: romout <= 16'hFFF2;
32'hFFFF1894: romout <= 16'h4CDF;
32'hFFFF1896: romout <= 16'h0203;
32'hFFFF1898: romout <= 16'h4E75;
32'hFFFF189A: romout <= 16'h6100;
32'hFFFF189C: romout <= 16'hFFDE;
32'hFFFF189E: romout <= 16'h6000;
32'hFFFF18A0: romout <= 16'hFE4C;
32'hFFFF18A2: romout <= 16'h0C41;
32'hFFFF18A4: romout <= 16'h00FF;
32'hFFFF18A6: romout <= 16'h670E;
32'hFFFF18A8: romout <= 16'h0C41;
32'hFFFF18AA: romout <= 16'hFF00;
32'hFFFF18AC: romout <= 16'h6714;
32'hFFFF18AE: romout <= 16'h4EB9;
32'hFFFF18B0: romout <= 16'hFFFF;
32'hFFFF18B2: romout <= 16'h18E8;
32'hFFFF18B4: romout <= 16'h4E75;
32'hFFFF18B6: romout <= 16'h3238;
32'hFFFF18B8: romout <= 16'h041A;
32'hFFFF18BA: romout <= 16'hE141;
32'hFFFF18BC: romout <= 16'h1238;
32'hFFFF18BE: romout <= 16'h0418;
32'hFFFF18C0: romout <= 16'h4E75;
32'hFFFF18C2: romout <= 16'h2F01;
32'hFFFF18C4: romout <= 16'h11C1;
32'hFFFF18C6: romout <= 16'h0418;
32'hFFFF18C8: romout <= 16'hE049;
32'hFFFF18CA: romout <= 16'h31C1;
32'hFFFF18CC: romout <= 16'h041A;
32'hFFFF18CE: romout <= 16'h3238;
32'hFFFF18D0: romout <= 16'h0418;
32'hFFFF18D2: romout <= 16'hC2F9;
32'hFFFF18D4: romout <= 16'hFFDA;
32'hFFFF18D6: romout <= 16'h0000;
32'hFFFF18D8: romout <= 16'hD278;
32'hFFFF18DA: romout <= 16'h041A;
32'hFFFF18DC: romout <= 16'hE341;
32'hFFFF18DE: romout <= 16'h33C1;
32'hFFFF18E0: romout <= 16'hFFDA;
32'hFFFF18E2: romout <= 16'h0016;
32'hFFFF18E4: romout <= 16'h221F;
32'hFFFF18E6: romout <= 16'h4E75;
32'hFFFF18E8: romout <= 16'h3239;
32'hFFFF18EA: romout <= 16'hFFDA;
32'hFFFF18EC: romout <= 16'h0000;
32'hFFFF18EE: romout <= 16'hC2F9;
32'hFFFF18F0: romout <= 16'hFFDA;
32'hFFFF18F2: romout <= 16'h0002;
32'hFFFF18F4: romout <= 16'h303C;
32'hFFFF18F6: romout <= 16'h0020;
32'hFFFF18F8: romout <= 16'h207C;
32'hFFFF18FA: romout <= 16'hFFD0;
32'hFFFF18FC: romout <= 16'h0000;
32'hFFFF18FE: romout <= 16'h30C0;
32'hFFFF1900: romout <= 16'h57C9;
32'hFFFF1902: romout <= 16'hFFFC;
32'hFFFF1904: romout <= 16'h3239;
32'hFFFF1906: romout <= 16'hFFDA;
32'hFFFF1908: romout <= 16'h0000;
32'hFFFF190A: romout <= 16'hC2F9;
32'hFFFF190C: romout <= 16'hFFDA;
32'hFFFF190E: romout <= 16'h0002;
32'hFFFF1910: romout <= 16'h3038;
32'hFFFF1912: romout <= 16'h0414;
32'hFFFF1914: romout <= 16'h207C;
32'hFFFF1916: romout <= 16'hFFD1;
32'hFFFF1918: romout <= 16'h0000;
32'hFFFF191A: romout <= 16'h30C0;
32'hFFFF191C: romout <= 16'h57C9;
32'hFFFF191E: romout <= 16'hFFFC;
32'hFFFF1920: romout <= 16'h4E75;
32'hFFFF1922: romout <= 16'h48E7;
32'hFFFF1924: romout <= 16'hE080;
32'hFFFF1926: romout <= 16'h3039;
32'hFFFF1928: romout <= 16'hFFDA;
32'hFFFF192A: romout <= 16'h0000;
32'hFFFF192C: romout <= 16'hC0F9;
32'hFFFF192E: romout <= 16'hFFDA;
32'hFFFF1930: romout <= 16'h0002;
32'hFFFF1932: romout <= 16'h9079;
32'hFFFF1934: romout <= 16'hFFDA;
32'hFFFF1936: romout <= 16'h0000;
32'hFFFF1938: romout <= 16'h41F9;
32'hFFFF193A: romout <= 16'hFFD0;
32'hFFFF193C: romout <= 16'h0000;
32'hFFFF193E: romout <= 16'h3439;
32'hFFFF1940: romout <= 16'hFFDA;
32'hFFFF1942: romout <= 16'h0000;
32'hFFFF1944: romout <= 16'hE342;
32'hFFFF1946: romout <= 16'h30F0;
32'hFFFF1948: romout <= 16'h2000;
32'hFFFF194A: romout <= 16'h57C8;
32'hFFFF194C: romout <= 16'hFFFA;
32'hFFFF194E: romout <= 16'h3239;
32'hFFFF1950: romout <= 16'hFFDA;
32'hFFFF1952: romout <= 16'h0002;
32'hFFFF1954: romout <= 16'h5341;
32'hFFFF1956: romout <= 16'h4EB9;
32'hFFFF1958: romout <= 16'hFFFF;
32'hFFFF195A: romout <= 16'h1962;
32'hFFFF195C: romout <= 16'h4CDF;
32'hFFFF195E: romout <= 16'h0107;
32'hFFFF1960: romout <= 16'h4E75;
32'hFFFF1962: romout <= 16'h48E7;
32'hFFFF1964: romout <= 16'h8080;
32'hFFFF1966: romout <= 16'h3039;
32'hFFFF1968: romout <= 16'hFFDA;
32'hFFFF196A: romout <= 16'h0000;
32'hFFFF196C: romout <= 16'hC0C1;
32'hFFFF196E: romout <= 16'hE340;
32'hFFFF1970: romout <= 16'h0680;
32'hFFFF1972: romout <= 16'hFFD0;
32'hFFFF1974: romout <= 16'h0000;
32'hFFFF1976: romout <= 16'h2040;
32'hFFFF1978: romout <= 16'h3039;
32'hFFFF197A: romout <= 16'hFFDA;
32'hFFFF197C: romout <= 16'h0000;
32'hFFFF197E: romout <= 16'h30FC;
32'hFFFF1980: romout <= 16'h0020;
32'hFFFF1982: romout <= 16'h57C8;
32'hFFFF1984: romout <= 16'hFFFA;
32'hFFFF1986: romout <= 16'h4CDF;
32'hFFFF1988: romout <= 16'h0101;
32'hFFFF198A: romout <= 16'h4E75;
32'hFFFF198C: romout <= 16'h48E7;
32'hFFFF198E: romout <= 16'hF800;
32'hFFFF1990: romout <= 16'h4284;
32'hFFFF1992: romout <= 16'h1802;
32'hFFFF1994: romout <= 16'h4EB9;
32'hFFFF1996: romout <= 16'hFFFF;
32'hFFFF1998: romout <= 16'h2F7A;
32'hFFFF199A: romout <= 16'h4CDF;
32'hFFFF199C: romout <= 16'h001F;
32'hFFFF199E: romout <= 16'h4E75;
32'hFFFF19A0: romout <= 16'h48E7;
32'hFFFF19A2: romout <= 16'hF800;
32'hFFFF19A4: romout <= 16'h4284;
32'hFFFF19A6: romout <= 16'h4EB9;
32'hFFFF19A8: romout <= 16'hFFFF;
32'hFFFF19AA: romout <= 16'h2F7A;
32'hFFFF19AC: romout <= 16'h4CDF;
32'hFFFF19AE: romout <= 16'h001F;
32'hFFFF19B0: romout <= 16'h4E75;
32'hFFFF19B2: romout <= 16'h0241;
32'hFFFF19B4: romout <= 16'h00FF;
32'hFFFF19B6: romout <= 16'h0C01;
32'hFFFF19B8: romout <= 16'h0041;
32'hFFFF19BA: romout <= 16'h6516;
32'hFFFF19BC: romout <= 16'h0C01;
32'hFFFF19BE: romout <= 16'h005A;
32'hFFFF19C0: romout <= 16'h6310;
32'hFFFF19C2: romout <= 16'h0C01;
32'hFFFF19C4: romout <= 16'h007A;
32'hFFFF19C6: romout <= 16'h620A;
32'hFFFF19C8: romout <= 16'h0C01;
32'hFFFF19CA: romout <= 16'h0061;
32'hFFFF19CC: romout <= 16'h6504;
32'hFFFF19CE: romout <= 16'h0401;
32'hFFFF19D0: romout <= 16'h0060;
32'hFFFF19D2: romout <= 16'h0041;
32'hFFFF19D4: romout <= 16'h0100;
32'hFFFF19D6: romout <= 16'h4E75;
32'hFFFF19D8: romout <= 16'h0201;
32'hFFFF19DA: romout <= 16'h00FF;
32'hFFFF19DC: romout <= 16'h0C01;
32'hFFFF19DE: romout <= 16'h001A;
32'hFFFF19E0: romout <= 16'h6204;
32'hFFFF19E2: romout <= 16'h0601;
32'hFFFF19E4: romout <= 16'h0060;
32'hFFFF19E6: romout <= 16'h4E75;
32'hFFFF19E8: romout <= 16'h3F01;
32'hFFFF19EA: romout <= 16'h0201;
32'hFFFF19EC: romout <= 16'h000F;
32'hFFFF19EE: romout <= 16'h0601;
32'hFFFF19F0: romout <= 16'h0030;
32'hFFFF19F2: romout <= 16'h0C01;
32'hFFFF19F4: romout <= 16'h0039;
32'hFFFF19F6: romout <= 16'h6302;
32'hFFFF19F8: romout <= 16'h5E01;
32'hFFFF19FA: romout <= 16'h6100;
32'hFFFF19FC: romout <= 16'hFD36;
32'hFFFF19FE: romout <= 16'h321F;
32'hFFFF1A00: romout <= 16'h4E75;
32'hFFFF1A02: romout <= 16'h3F01;
32'hFFFF1A04: romout <= 16'hE819;
32'hFFFF1A06: romout <= 16'h6100;
32'hFFFF1A08: romout <= 16'hFFE0;
32'hFFFF1A0A: romout <= 16'hE919;
32'hFFFF1A0C: romout <= 16'h6100;
32'hFFFF1A0E: romout <= 16'hFFDA;
32'hFFFF1A10: romout <= 16'h321F;
32'hFFFF1A12: romout <= 16'h4E75;
32'hFFFF1A14: romout <= 16'hE199;
32'hFFFF1A16: romout <= 16'h6100;
32'hFFFF1A18: romout <= 16'hFFEA;
32'hFFFF1A1A: romout <= 16'hE199;
32'hFFFF1A1C: romout <= 16'h6100;
32'hFFFF1A1E: romout <= 16'hFFE4;
32'hFFFF1A20: romout <= 16'hE199;
32'hFFFF1A22: romout <= 16'h6100;
32'hFFFF1A24: romout <= 16'hFFDE;
32'hFFFF1A26: romout <= 16'hE199;
32'hFFFF1A28: romout <= 16'h6100;
32'hFFFF1A2A: romout <= 16'hFFD8;
32'hFFFF1A2C: romout <= 16'h4E75;
32'hFFFF1A2E: romout <= 16'h123C;
32'hFFFF1A30: romout <= 16'h003A;
32'hFFFF1A32: romout <= 16'h4EB9;
32'hFFFF1A34: romout <= 16'hFFFF;
32'hFFFF1A36: romout <= 16'h1732;
32'hFFFF1A38: romout <= 16'h2208;
32'hFFFF1A3A: romout <= 16'h4EB9;
32'hFFFF1A3C: romout <= 16'hFFFF;
32'hFFFF1A3E: romout <= 16'h1A14;
32'hFFFF1A40: romout <= 16'h7407;
32'hFFFF1A42: romout <= 16'h123C;
32'hFFFF1A44: romout <= 16'h0020;
32'hFFFF1A46: romout <= 16'h4EB9;
32'hFFFF1A48: romout <= 16'hFFFF;
32'hFFFF1A4A: romout <= 16'h1732;
32'hFFFF1A4C: romout <= 16'h1218;
32'hFFFF1A4E: romout <= 16'h4EB9;
32'hFFFF1A50: romout <= 16'hFFFF;
32'hFFFF1A52: romout <= 16'h1A02;
32'hFFFF1A54: romout <= 16'h51CA;
32'hFFFF1A56: romout <= 16'hFFEC;
32'hFFFF1A58: romout <= 16'h4EF9;
32'hFFFF1A5A: romout <= 16'hFFFF;
32'hFFFF1A5C: romout <= 16'h16EC;
32'hFFFF1A5E: romout <= 16'h4E55;
32'hFFFF1A60: romout <= 16'hFFE8;
32'hFFFF1A62: romout <= 16'h41ED;
32'hFFFF1A64: romout <= 16'hFFFA;
32'hFFFF1A66: romout <= 16'h43ED;
32'hFFFF1A68: romout <= 16'hFFFC;
32'hFFFF1A6A: romout <= 16'h3B7C;
32'hFFFF1A6C: romout <= 16'h0000;
32'hFFFF1A6E: romout <= 16'hFFFA;
32'hFFFF1A70: romout <= 16'h3B7C;
32'hFFFF1A72: romout <= 16'h0002;
32'hFFFF1A74: romout <= 16'hFFF8;
32'hFFFF1A76: romout <= 16'h7048;
32'hFFFF1A78: romout <= 16'h4E41;
32'hFFFF1A7A: romout <= 16'h4278;
32'hFFFF1A7C: romout <= 16'h041C;
32'hFFFF1A7E: romout <= 16'h6100;
32'hFFFF1A80: romout <= 16'hFC6C;
32'hFFFF1A82: romout <= 16'h123C;
32'hFFFF1A84: romout <= 16'h0024;
32'hFFFF1A86: romout <= 16'h6100;
32'hFFFF1A88: romout <= 16'hFCAA;
32'hFFFF1A8A: romout <= 16'h6100;
32'hFFFF1A8C: romout <= 16'hFBCC;
32'hFFFF1A8E: romout <= 16'h0C01;
32'hFFFF1A90: romout <= 16'h000D;
32'hFFFF1A92: romout <= 16'h6706;
32'hFFFF1A94: romout <= 16'h6100;
32'hFFFF1A96: romout <= 16'hFC9C;
32'hFFFF1A98: romout <= 16'h60F0;
32'hFFFF1A9A: romout <= 16'h4278;
32'hFFFF1A9C: romout <= 16'h041A;
32'hFFFF1A9E: romout <= 16'h6100;
32'hFFFF1AA0: romout <= 16'hFC66;
32'hFFFF1AA2: romout <= 16'h3218;
32'hFFFF1AA4: romout <= 16'h6100;
32'hFFFF1AA6: romout <= 16'hFF32;
32'hFFFF1AA8: romout <= 16'h0C01;
32'hFFFF1AAA: romout <= 16'h0024;
32'hFFFF1AAC: romout <= 16'h6606;
32'hFFFF1AAE: romout <= 16'h3218;
32'hFFFF1AB0: romout <= 16'h6100;
32'hFFFF1AB2: romout <= 16'hFF26;
32'hFFFF1AB4: romout <= 16'h0C01;
32'hFFFF1AB6: romout <= 16'h003A;
32'hFFFF1AB8: romout <= 16'h6700;
32'hFFFF1ABA: romout <= 16'h00FC;
32'hFFFF1ABC: romout <= 16'h0C01;
32'hFFFF1ABE: romout <= 16'h0044;
32'hFFFF1AC0: romout <= 16'h6700;
32'hFFFF1AC2: romout <= 16'h0162;
32'hFFFF1AC4: romout <= 16'h0C01;
32'hFFFF1AC6: romout <= 16'h0042;
32'hFFFF1AC8: romout <= 16'h6700;
32'hFFFF1ACA: romout <= 16'h0936;
32'hFFFF1ACC: romout <= 16'h0C01;
32'hFFFF1ACE: romout <= 16'h004A;
32'hFFFF1AD0: romout <= 16'h6700;
32'hFFFF1AD2: romout <= 16'h0142;
32'hFFFF1AD4: romout <= 16'h0C01;
32'hFFFF1AD6: romout <= 16'h004C;
32'hFFFF1AD8: romout <= 16'h6700;
32'hFFFF1ADA: romout <= 16'h01EE;
32'hFFFF1ADC: romout <= 16'h0C01;
32'hFFFF1ADE: romout <= 16'h003F;
32'hFFFF1AE0: romout <= 16'h672A;
32'hFFFF1AE2: romout <= 16'h0C01;
32'hFFFF1AE4: romout <= 16'h0043;
32'hFFFF1AE6: romout <= 16'h6702;
32'hFFFF1AE8: romout <= 16'h6090;
32'hFFFF1AEA: romout <= 16'h3218;
32'hFFFF1AEC: romout <= 16'h6100;
32'hFFFF1AEE: romout <= 16'hFEEA;
32'hFFFF1AF0: romout <= 16'h0C01;
32'hFFFF1AF2: romout <= 16'h004C;
32'hFFFF1AF4: romout <= 16'h6684;
32'hFFFF1AF6: romout <= 16'h3218;
32'hFFFF1AF8: romout <= 16'h6100;
32'hFFFF1AFA: romout <= 16'hFEDE;
32'hFFFF1AFC: romout <= 16'h0C01;
32'hFFFF1AFE: romout <= 16'h0053;
32'hFFFF1B00: romout <= 16'h6600;
32'hFFFF1B02: romout <= 16'hFF78;
32'hFFFF1B04: romout <= 16'h6100;
32'hFFFF1B06: romout <= 16'hFDE2;
32'hFFFF1B08: romout <= 16'h6000;
32'hFFFF1B0A: romout <= 16'hFF70;
32'hFFFF1B0C: romout <= 16'h43F9;
32'hFFFF1B0E: romout <= 16'hFFFF;
32'hFFFF1B10: romout <= 16'h1B1C;
32'hFFFF1B12: romout <= 16'h4EB9;
32'hFFFF1B14: romout <= 16'hFFFF;
32'hFFFF1B16: romout <= 16'h1858;
32'hFFFF1B18: romout <= 16'h6000;
32'hFFFF1B1A: romout <= 16'hFF60;
32'hFFFF1B1C: romout <= 16'h3F20;
32'hFFFF1B1E: romout <= 16'h3D20;
32'hFFFF1B20: romout <= 16'h4469;
32'hFFFF1B22: romout <= 16'h7370;
32'hFFFF1B24: romout <= 16'h6C61;
32'hFFFF1B26: romout <= 16'h7920;
32'hFFFF1B28: romout <= 16'h6865;
32'hFFFF1B2A: romout <= 16'h6C70;
32'hFFFF1B2C: romout <= 16'h0D0A;
32'hFFFF1B2E: romout <= 16'h434C;
32'hFFFF1B30: romout <= 16'h5320;
32'hFFFF1B32: romout <= 16'h3D20;
32'hFFFF1B34: romout <= 16'h636C;
32'hFFFF1B36: romout <= 16'h6561;
32'hFFFF1B38: romout <= 16'h7220;
32'hFFFF1B3A: romout <= 16'h7363;
32'hFFFF1B3C: romout <= 16'h7265;
32'hFFFF1B3E: romout <= 16'h656E;
32'hFFFF1B40: romout <= 16'h0D0A;
32'hFFFF1B42: romout <= 16'h3A20;
32'hFFFF1B44: romout <= 16'h3D20;
32'hFFFF1B46: romout <= 16'h4564;
32'hFFFF1B48: romout <= 16'h6974;
32'hFFFF1B4A: romout <= 16'h206D;
32'hFFFF1B4C: romout <= 16'h656D;
32'hFFFF1B4E: romout <= 16'h6F72;
32'hFFFF1B50: romout <= 16'h7920;
32'hFFFF1B52: romout <= 16'h6279;
32'hFFFF1B54: romout <= 16'h7465;
32'hFFFF1B56: romout <= 16'h730D;
32'hFFFF1B58: romout <= 16'h0A4C;
32'hFFFF1B5A: romout <= 16'h203D;
32'hFFFF1B5C: romout <= 16'h204C;
32'hFFFF1B5E: romout <= 16'h6F61;
32'hFFFF1B60: romout <= 16'h6420;
32'hFFFF1B62: romout <= 16'h5331;
32'hFFFF1B64: romout <= 16'h3920;
32'hFFFF1B66: romout <= 16'h6669;
32'hFFFF1B68: romout <= 16'h6C65;
32'hFFFF1B6A: romout <= 16'h0D0A;
32'hFFFF1B6C: romout <= 16'h4420;
32'hFFFF1B6E: romout <= 16'h3D20;
32'hFFFF1B70: romout <= 16'h4475;
32'hFFFF1B72: romout <= 16'h6D70;
32'hFFFF1B74: romout <= 16'h206D;
32'hFFFF1B76: romout <= 16'h656D;
32'hFFFF1B78: romout <= 16'h6F72;
32'hFFFF1B7A: romout <= 16'h790D;
32'hFFFF1B7C: romout <= 16'h0A42;
32'hFFFF1B7E: romout <= 16'h203D;
32'hFFFF1B80: romout <= 16'h2073;
32'hFFFF1B82: romout <= 16'h7461;
32'hFFFF1B84: romout <= 16'h7274;
32'hFFFF1B86: romout <= 16'h2074;
32'hFFFF1B88: romout <= 16'h696E;
32'hFFFF1B8A: romout <= 16'h7920;
32'hFFFF1B8C: romout <= 16'h6261;
32'hFFFF1B8E: romout <= 16'h7369;
32'hFFFF1B90: romout <= 16'h630D;
32'hFFFF1B92: romout <= 16'h0A4A;
32'hFFFF1B94: romout <= 16'h203D;
32'hFFFF1B96: romout <= 16'h204A;
32'hFFFF1B98: romout <= 16'h756D;
32'hFFFF1B9A: romout <= 16'h7020;
32'hFFFF1B9C: romout <= 16'h746F;
32'hFFFF1B9E: romout <= 16'h2063;
32'hFFFF1BA0: romout <= 16'h6F64;
32'hFFFF1BA2: romout <= 16'h650D;
32'hFFFF1BA4: romout <= 16'h0A00;
32'hFFFF1BA6: romout <= 16'h3218;
32'hFFFF1BA8: romout <= 16'h6100;
32'hFFFF1BAA: romout <= 16'hFE2E;
32'hFFFF1BAC: romout <= 16'h0C01;
32'hFFFF1BAE: romout <= 16'h0020;
32'hFFFF1BB0: romout <= 16'h67F4;
32'hFFFF1BB2: romout <= 16'h5588;
32'hFFFF1BB4: romout <= 16'h4E75;
32'hFFFF1BB6: romout <= 16'h6100;
32'hFFFF1BB8: romout <= 16'hFFEE;
32'hFFFF1BBA: romout <= 16'h6100;
32'hFFFF1BBC: romout <= 16'h009C;
32'hFFFF1BBE: romout <= 16'h2241;
32'hFFFF1BC0: romout <= 16'h6100;
32'hFFFF1BC2: romout <= 16'hFFE4;
32'hFFFF1BC4: romout <= 16'h6100;
32'hFFFF1BC6: romout <= 16'h0092;
32'hFFFF1BC8: romout <= 16'h12C1;
32'hFFFF1BCA: romout <= 16'h6100;
32'hFFFF1BCC: romout <= 16'hFFDA;
32'hFFFF1BCE: romout <= 16'h6100;
32'hFFFF1BD0: romout <= 16'h0088;
32'hFFFF1BD2: romout <= 16'h12C1;
32'hFFFF1BD4: romout <= 16'h6100;
32'hFFFF1BD6: romout <= 16'hFFD0;
32'hFFFF1BD8: romout <= 16'h6100;
32'hFFFF1BDA: romout <= 16'h007E;
32'hFFFF1BDC: romout <= 16'h12C1;
32'hFFFF1BDE: romout <= 16'h6100;
32'hFFFF1BE0: romout <= 16'hFFC6;
32'hFFFF1BE2: romout <= 16'h6100;
32'hFFFF1BE4: romout <= 16'h0074;
32'hFFFF1BE6: romout <= 16'h12C1;
32'hFFFF1BE8: romout <= 16'h6100;
32'hFFFF1BEA: romout <= 16'hFFBC;
32'hFFFF1BEC: romout <= 16'h6100;
32'hFFFF1BEE: romout <= 16'h006A;
32'hFFFF1BF0: romout <= 16'h12C1;
32'hFFFF1BF2: romout <= 16'h6100;
32'hFFFF1BF4: romout <= 16'hFFB2;
32'hFFFF1BF6: romout <= 16'h6100;
32'hFFFF1BF8: romout <= 16'h0060;
32'hFFFF1BFA: romout <= 16'h12C1;
32'hFFFF1BFC: romout <= 16'h6100;
32'hFFFF1BFE: romout <= 16'hFFA8;
32'hFFFF1C00: romout <= 16'h6100;
32'hFFFF1C02: romout <= 16'h0056;
32'hFFFF1C04: romout <= 16'h12C1;
32'hFFFF1C06: romout <= 16'h6100;
32'hFFFF1C08: romout <= 16'hFF9E;
32'hFFFF1C0A: romout <= 16'h6100;
32'hFFFF1C0C: romout <= 16'h004C;
32'hFFFF1C0E: romout <= 16'h12C1;
32'hFFFF1C10: romout <= 16'h6000;
32'hFFFF1C12: romout <= 16'hFE68;
32'hFFFF1C14: romout <= 16'h6100;
32'hFFFF1C16: romout <= 16'hFF90;
32'hFFFF1C18: romout <= 16'h6100;
32'hFFFF1C1A: romout <= 16'h003E;
32'hFFFF1C1C: romout <= 16'h2041;
32'hFFFF1C1E: romout <= 16'h4E90;
32'hFFFF1C20: romout <= 16'h6000;
32'hFFFF1C22: romout <= 16'hFE58;
32'hFFFF1C24: romout <= 16'h6100;
32'hFFFF1C26: romout <= 16'hFF80;
32'hFFFF1C28: romout <= 16'h6100;
32'hFFFF1C2A: romout <= 16'h002E;
32'hFFFF1C2C: romout <= 16'h2041;
32'hFFFF1C2E: romout <= 16'h4EB9;
32'hFFFF1C30: romout <= 16'hFFFF;
32'hFFFF1C32: romout <= 16'h16EC;
32'hFFFF1C34: romout <= 16'h6100;
32'hFFFF1C36: romout <= 16'hFDF8;
32'hFFFF1C38: romout <= 16'h6100;
32'hFFFF1C3A: romout <= 16'hFDF4;
32'hFFFF1C3C: romout <= 16'h6100;
32'hFFFF1C3E: romout <= 16'hFDF0;
32'hFFFF1C40: romout <= 16'h6100;
32'hFFFF1C42: romout <= 16'hFDEC;
32'hFFFF1C44: romout <= 16'h6100;
32'hFFFF1C46: romout <= 16'hFDE8;
32'hFFFF1C48: romout <= 16'h6100;
32'hFFFF1C4A: romout <= 16'hFDE4;
32'hFFFF1C4C: romout <= 16'h6100;
32'hFFFF1C4E: romout <= 16'hFDE0;
32'hFFFF1C50: romout <= 16'h6100;
32'hFFFF1C52: romout <= 16'hFDDC;
32'hFFFF1C54: romout <= 16'h6000;
32'hFFFF1C56: romout <= 16'hFE24;
32'hFFFF1C58: romout <= 16'h48E7;
32'hFFFF1C5A: romout <= 16'hA000;
32'hFFFF1C5C: romout <= 16'h4282;
32'hFFFF1C5E: romout <= 16'h7007;
32'hFFFF1C60: romout <= 16'h3218;
32'hFFFF1C62: romout <= 16'h6100;
32'hFFFF1C64: romout <= 16'hFD74;
32'hFFFF1C66: romout <= 16'h6100;
32'hFFFF1C68: romout <= 16'h001E;
32'hFFFF1C6A: romout <= 16'hB23C;
32'hFFFF1C6C: romout <= 16'h00FF;
32'hFFFF1C6E: romout <= 16'h670E;
32'hFFFF1C70: romout <= 16'hE98A;
32'hFFFF1C72: romout <= 16'h0281;
32'hFFFF1C74: romout <= 16'h0000;
32'hFFFF1C76: romout <= 16'h000F;
32'hFFFF1C78: romout <= 16'h8481;
32'hFFFF1C7A: romout <= 16'h51C8;
32'hFFFF1C7C: romout <= 16'hFFE4;
32'hFFFF1C7E: romout <= 16'h2202;
32'hFFFF1C80: romout <= 16'h4CDF;
32'hFFFF1C82: romout <= 16'h0005;
32'hFFFF1C84: romout <= 16'h4E75;
32'hFFFF1C86: romout <= 16'h0C01;
32'hFFFF1C88: romout <= 16'h0030;
32'hFFFF1C8A: romout <= 16'h6538;
32'hFFFF1C8C: romout <= 16'h0C01;
32'hFFFF1C8E: romout <= 16'h0039;
32'hFFFF1C90: romout <= 16'h6206;
32'hFFFF1C92: romout <= 16'h0401;
32'hFFFF1C94: romout <= 16'h0030;
32'hFFFF1C96: romout <= 16'h4E75;
32'hFFFF1C98: romout <= 16'h0C01;
32'hFFFF1C9A: romout <= 16'h0041;
32'hFFFF1C9C: romout <= 16'h6526;
32'hFFFF1C9E: romout <= 16'h0C01;
32'hFFFF1CA0: romout <= 16'h0046;
32'hFFFF1CA2: romout <= 16'h620A;
32'hFFFF1CA4: romout <= 16'h0401;
32'hFFFF1CA6: romout <= 16'h0041;
32'hFFFF1CA8: romout <= 16'h0601;
32'hFFFF1CAA: romout <= 16'h000A;
32'hFFFF1CAC: romout <= 16'h4E75;
32'hFFFF1CAE: romout <= 16'h0C01;
32'hFFFF1CB0: romout <= 16'h0061;
32'hFFFF1CB2: romout <= 16'h6510;
32'hFFFF1CB4: romout <= 16'h0C01;
32'hFFFF1CB6: romout <= 16'h0066;
32'hFFFF1CB8: romout <= 16'h620A;
32'hFFFF1CBA: romout <= 16'h0401;
32'hFFFF1CBC: romout <= 16'h0061;
32'hFFFF1CBE: romout <= 16'h0601;
32'hFFFF1CC0: romout <= 16'h000A;
32'hFFFF1CC2: romout <= 16'h4E75;
32'hFFFF1CC4: romout <= 16'h72FF;
32'hFFFF1CC6: romout <= 16'h4E75;
32'hFFFF1CC8: romout <= 16'h600A;
32'hFFFF1CCA: romout <= 16'h6100;
32'hFFFF1CCC: romout <= 16'h0174;
32'hFFFF1CCE: romout <= 16'h0C00;
32'hFFFF1CD0: romout <= 16'h000A;
32'hFFFF1CD2: romout <= 16'h66F6;
32'hFFFF1CD4: romout <= 16'h6100;
32'hFFFF1CD6: romout <= 16'h016A;
32'hFFFF1CD8: romout <= 16'h1800;
32'hFFFF1CDA: romout <= 16'h0C04;
32'hFFFF1CDC: romout <= 16'h001A;
32'hFFFF1CDE: romout <= 16'h6700;
32'hFFFF1CE0: romout <= 16'hFD9A;
32'hFFFF1CE2: romout <= 16'h0C04;
32'hFFFF1CE4: romout <= 16'h0053;
32'hFFFF1CE6: romout <= 16'h66E2;
32'hFFFF1CE8: romout <= 16'h6100;
32'hFFFF1CEA: romout <= 16'h0156;
32'hFFFF1CEC: romout <= 16'h1800;
32'hFFFF1CEE: romout <= 16'h0C04;
32'hFFFF1CF0: romout <= 16'h0030;
32'hFFFF1CF2: romout <= 16'h65D6;
32'hFFFF1CF4: romout <= 16'h0C04;
32'hFFFF1CF6: romout <= 16'h0039;
32'hFFFF1CF8: romout <= 16'h62D0;
32'hFFFF1CFA: romout <= 16'h6100;
32'hFFFF1CFC: romout <= 16'h0144;
32'hFFFF1CFE: romout <= 16'h6100;
32'hFFFF1D00: romout <= 16'hFF86;
32'hFFFF1D02: romout <= 16'h1401;
32'hFFFF1D04: romout <= 16'h6100;
32'hFFFF1D06: romout <= 16'h013A;
32'hFFFF1D08: romout <= 16'h6100;
32'hFFFF1D0A: romout <= 16'hFF7C;
32'hFFFF1D0C: romout <= 16'hE90A;
32'hFFFF1D0E: romout <= 16'h8202;
32'hFFFF1D10: romout <= 16'h1601;
32'hFFFF1D12: romout <= 16'h0C04;
32'hFFFF1D14: romout <= 16'h0030;
32'hFFFF1D16: romout <= 16'h67B2;
32'hFFFF1D18: romout <= 16'h0C04;
32'hFFFF1D1A: romout <= 16'h0031;
32'hFFFF1D1C: romout <= 16'h676A;
32'hFFFF1D1E: romout <= 16'h0C04;
32'hFFFF1D20: romout <= 16'h0032;
32'hFFFF1D22: romout <= 16'h676A;
32'hFFFF1D24: romout <= 16'h0C04;
32'hFFFF1D26: romout <= 16'h0033;
32'hFFFF1D28: romout <= 16'h676A;
32'hFFFF1D2A: romout <= 16'h0C04;
32'hFFFF1D2C: romout <= 16'h0035;
32'hFFFF1D2E: romout <= 16'h679A;
32'hFFFF1D30: romout <= 16'h0C04;
32'hFFFF1D32: romout <= 16'h0037;
32'hFFFF1D34: romout <= 16'h6764;
32'hFFFF1D36: romout <= 16'h0C04;
32'hFFFF1D38: romout <= 16'h0038;
32'hFFFF1D3A: romout <= 16'h676A;
32'hFFFF1D3C: romout <= 16'h0C04;
32'hFFFF1D3E: romout <= 16'h0039;
32'hFFFF1D40: romout <= 16'h6770;
32'hFFFF1D42: romout <= 16'h6086;
32'hFFFF1D44: romout <= 16'h0243;
32'hFFFF1D46: romout <= 16'h00FF;
32'hFFFF1D48: romout <= 16'h5343;
32'hFFFF1D4A: romout <= 16'h4282;
32'hFFFF1D4C: romout <= 16'h6100;
32'hFFFF1D4E: romout <= 16'h00F2;
32'hFFFF1D50: romout <= 16'h6100;
32'hFFFF1D52: romout <= 16'hFF34;
32'hFFFF1D54: romout <= 16'hE98A;
32'hFFFF1D56: romout <= 16'h8401;
32'hFFFF1D58: romout <= 16'h6100;
32'hFFFF1D5A: romout <= 16'h00E6;
32'hFFFF1D5C: romout <= 16'h6100;
32'hFFFF1D5E: romout <= 16'hFF28;
32'hFFFF1D60: romout <= 16'hE98A;
32'hFFFF1D62: romout <= 16'h8401;
32'hFFFF1D64: romout <= 16'h12C2;
32'hFFFF1D66: romout <= 16'h51CB;
32'hFFFF1D68: romout <= 16'hFFE2;
32'hFFFF1D6A: romout <= 16'h4282;
32'hFFFF1D6C: romout <= 16'h6100;
32'hFFFF1D6E: romout <= 16'h00D2;
32'hFFFF1D70: romout <= 16'h6100;
32'hFFFF1D72: romout <= 16'hFF14;
32'hFFFF1D74: romout <= 16'hE98A;
32'hFFFF1D76: romout <= 16'h8401;
32'hFFFF1D78: romout <= 16'h6100;
32'hFFFF1D7A: romout <= 16'h00C6;
32'hFFFF1D7C: romout <= 16'h6100;
32'hFFFF1D7E: romout <= 16'hFF08;
32'hFFFF1D80: romout <= 16'hE98A;
32'hFFFF1D82: romout <= 16'h8401;
32'hFFFF1D84: romout <= 16'h6000;
32'hFFFF1D86: romout <= 16'hFF44;
32'hFFFF1D88: romout <= 16'h6100;
32'hFFFF1D8A: romout <= 16'h0034;
32'hFFFF1D8C: romout <= 16'h60B6;
32'hFFFF1D8E: romout <= 16'h6100;
32'hFFFF1D90: romout <= 16'h003C;
32'hFFFF1D92: romout <= 16'h60B0;
32'hFFFF1D94: romout <= 16'h6100;
32'hFFFF1D96: romout <= 16'h0044;
32'hFFFF1D98: romout <= 16'h60AA;
32'hFFFF1D9A: romout <= 16'h6100;
32'hFFFF1D9C: romout <= 16'h003E;
32'hFFFF1D9E: romout <= 16'h21C9;
32'hFFFF1DA0: romout <= 16'h0800;
32'hFFFF1DA2: romout <= 16'h6000;
32'hFFFF1DA4: romout <= 16'hFCD6;
32'hFFFF1DA6: romout <= 16'h6100;
32'hFFFF1DA8: romout <= 16'h0024;
32'hFFFF1DAA: romout <= 16'h21C9;
32'hFFFF1DAC: romout <= 16'h0800;
32'hFFFF1DAE: romout <= 16'h6000;
32'hFFFF1DB0: romout <= 16'hFCCA;
32'hFFFF1DB2: romout <= 16'h6100;
32'hFFFF1DB4: romout <= 16'h000A;
32'hFFFF1DB6: romout <= 16'h21C9;
32'hFFFF1DB8: romout <= 16'h0800;
32'hFFFF1DBA: romout <= 16'h6000;
32'hFFFF1DBC: romout <= 16'hFCBE;
32'hFFFF1DBE: romout <= 16'h4282;
32'hFFFF1DC0: romout <= 16'h6100;
32'hFFFF1DC2: romout <= 16'h007E;
32'hFFFF1DC4: romout <= 16'h6100;
32'hFFFF1DC6: romout <= 16'hFEC0;
32'hFFFF1DC8: romout <= 16'h1401;
32'hFFFF1DCA: romout <= 16'h604A;
32'hFFFF1DCC: romout <= 16'h4282;
32'hFFFF1DCE: romout <= 16'h6100;
32'hFFFF1DD0: romout <= 16'h0070;
32'hFFFF1DD2: romout <= 16'h6100;
32'hFFFF1DD4: romout <= 16'hFEB2;
32'hFFFF1DD6: romout <= 16'h1401;
32'hFFFF1DD8: romout <= 16'h6024;
32'hFFFF1DDA: romout <= 16'h4282;
32'hFFFF1DDC: romout <= 16'h6100;
32'hFFFF1DDE: romout <= 16'h0062;
32'hFFFF1DE0: romout <= 16'h6100;
32'hFFFF1DE2: romout <= 16'hFEA4;
32'hFFFF1DE4: romout <= 16'h1401;
32'hFFFF1DE6: romout <= 16'h6100;
32'hFFFF1DE8: romout <= 16'h0058;
32'hFFFF1DEA: romout <= 16'h6100;
32'hFFFF1DEC: romout <= 16'hFE9A;
32'hFFFF1DEE: romout <= 16'hE98A;
32'hFFFF1DF0: romout <= 16'h8401;
32'hFFFF1DF2: romout <= 16'h6100;
32'hFFFF1DF4: romout <= 16'h004C;
32'hFFFF1DF6: romout <= 16'h6100;
32'hFFFF1DF8: romout <= 16'hFE8E;
32'hFFFF1DFA: romout <= 16'hE98A;
32'hFFFF1DFC: romout <= 16'h8401;
32'hFFFF1DFE: romout <= 16'h6100;
32'hFFFF1E00: romout <= 16'h0040;
32'hFFFF1E02: romout <= 16'h6100;
32'hFFFF1E04: romout <= 16'hFE82;
32'hFFFF1E06: romout <= 16'hE98A;
32'hFFFF1E08: romout <= 16'h8401;
32'hFFFF1E0A: romout <= 16'h6100;
32'hFFFF1E0C: romout <= 16'h0034;
32'hFFFF1E0E: romout <= 16'h6100;
32'hFFFF1E10: romout <= 16'hFE76;
32'hFFFF1E12: romout <= 16'hE98A;
32'hFFFF1E14: romout <= 16'h8401;
32'hFFFF1E16: romout <= 16'h6100;
32'hFFFF1E18: romout <= 16'h0028;
32'hFFFF1E1A: romout <= 16'h6100;
32'hFFFF1E1C: romout <= 16'hFE6A;
32'hFFFF1E1E: romout <= 16'hE98A;
32'hFFFF1E20: romout <= 16'h8401;
32'hFFFF1E22: romout <= 16'h6100;
32'hFFFF1E24: romout <= 16'h001C;
32'hFFFF1E26: romout <= 16'h6100;
32'hFFFF1E28: romout <= 16'hFE5E;
32'hFFFF1E2A: romout <= 16'hE98A;
32'hFFFF1E2C: romout <= 16'h8401;
32'hFFFF1E2E: romout <= 16'h6100;
32'hFFFF1E30: romout <= 16'h0010;
32'hFFFF1E32: romout <= 16'h6100;
32'hFFFF1E34: romout <= 16'hFE52;
32'hFFFF1E36: romout <= 16'hE98A;
32'hFFFF1E38: romout <= 16'h8401;
32'hFFFF1E3A: romout <= 16'h4284;
32'hFFFF1E3C: romout <= 16'h2242;
32'hFFFF1E3E: romout <= 16'h4E75;
32'hFFFF1E40: romout <= 16'h6100;
32'hFFFF1E42: romout <= 16'hF898;
32'hFFFF1E44: romout <= 16'h670C;
32'hFFFF1E46: romout <= 16'h6100;
32'hFFFF1E48: romout <= 16'hF810;
32'hFFFF1E4A: romout <= 16'h0C01;
32'hFFFF1E4C: romout <= 16'h0003;
32'hFFFF1E4E: romout <= 16'h6700;
32'hFFFF1E50: romout <= 16'hFC2A;
32'hFFFF1E52: romout <= 16'h6100;
32'hFFFF1E54: romout <= 16'h1288;
32'hFFFF1E56: romout <= 16'h67E8;
32'hFFFF1E58: romout <= 16'h1200;
32'hFFFF1E5A: romout <= 16'h4E75;
32'hFFFF1E5C: romout <= 16'h33FC;
32'hFFFF1E5E: romout <= 16'h000F;
32'hFFFF1E60: romout <= 16'hFFD4;
32'hFFFF1E62: romout <= 16'h0040;
32'hFFFF1E64: romout <= 16'h33FC;
32'hFFFF1E66: romout <= 16'h411B;
32'hFFFF1E68: romout <= 16'hFFD4;
32'hFFFF1E6A: romout <= 16'h0000;
32'hFFFF1E6C: romout <= 16'h4279;
32'hFFFF1E6E: romout <= 16'hFFD4;
32'hFFFF1E70: romout <= 16'h0002;
32'hFFFF1E72: romout <= 16'h4279;
32'hFFFF1E74: romout <= 16'hFFD4;
32'hFFFF1E76: romout <= 16'h0008;
32'hFFFF1E78: romout <= 16'h4279;
32'hFFFF1E7A: romout <= 16'hFFD4;
32'hFFFF1E7C: romout <= 16'h000A;
32'hFFFF1E7E: romout <= 16'h33FC;
32'hFFFF1E80: romout <= 16'h00FF;
32'hFFFF1E82: romout <= 16'hFFD4;
32'hFFFF1E84: romout <= 16'h000C;
32'hFFFF1E86: romout <= 16'h4279;
32'hFFFF1E88: romout <= 16'hFFD4;
32'hFFFF1E8A: romout <= 16'h000E;
32'hFFFF1E8C: romout <= 16'h33FC;
32'hFFFF1E8E: romout <= 16'h1104;
32'hFFFF1E90: romout <= 16'hFFD4;
32'hFFFF1E92: romout <= 16'h0004;
32'hFFFF1E94: romout <= 16'h203C;
32'hFFFF1E96: romout <= 16'h007A;
32'hFFFF1E98: romout <= 16'h1200;
32'hFFFF1E9A: romout <= 16'h5380;
32'hFFFF1E9C: romout <= 16'h66FC;
32'hFFFF1E9E: romout <= 16'h4279;
32'hFFFF1EA0: romout <= 16'hFFD4;
32'hFFFF1EA2: romout <= 16'h0004;
32'hFFFF1EA4: romout <= 16'h33FC;
32'hFFFF1EA6: romout <= 16'h0000;
32'hFFFF1EA8: romout <= 16'hFFD4;
32'hFFFF1EAA: romout <= 16'h0040;
32'hFFFF1EAC: romout <= 16'h4E75;
32'hFFFF1EAE: romout <= 16'h303C;
32'hFFFF1EB0: romout <= 16'h5151;
32'hFFFF1EB2: romout <= 16'h33C0;
32'hFFFF1EB4: romout <= 16'hFFDC;
32'hFFFF1EB6: romout <= 16'h0300;
32'hFFFF1EB8: romout <= 16'h0839;
32'hFFFF1EBA: romout <= 16'h0007;
32'hFFFF1EBC: romout <= 16'hFFDC;
32'hFFFF1EBE: romout <= 16'h0303;
32'hFFFF1EC0: romout <= 16'h66F6;
32'hFFFF1EC2: romout <= 16'h203C;
32'hFFFF1EC4: romout <= 16'h007A;
32'hFFFF1EC6: romout <= 16'h1200;
32'hFFFF1EC8: romout <= 16'h5380;
32'hFFFF1ECA: romout <= 16'h66FC;
32'hFFFF1ECC: romout <= 16'h303C;
32'hFFFF1ECE: romout <= 16'hACAC;
32'hFFFF1ED0: romout <= 16'h33C0;
32'hFFFF1ED2: romout <= 16'hFFDC;
32'hFFFF1ED4: romout <= 16'h0300;
32'hFFFF1ED6: romout <= 16'h0839;
32'hFFFF1ED8: romout <= 16'h0007;
32'hFFFF1EDA: romout <= 16'hFFDC;
32'hFFFF1EDC: romout <= 16'h0303;
32'hFFFF1EDE: romout <= 16'h66F6;
32'hFFFF1EE0: romout <= 16'h3039;
32'hFFFF1EE2: romout <= 16'hFFDC;
32'hFFFF1EE4: romout <= 16'h0302;
32'hFFFF1EE6: romout <= 16'h4840;
32'hFFFF1EE8: romout <= 16'h303C;
32'hFFFF1EEA: romout <= 16'hAAAA;
32'hFFFF1EEC: romout <= 16'h33C0;
32'hFFFF1EEE: romout <= 16'hFFDC;
32'hFFFF1EF0: romout <= 16'h0300;
32'hFFFF1EF2: romout <= 16'h0839;
32'hFFFF1EF4: romout <= 16'h0007;
32'hFFFF1EF6: romout <= 16'hFFDC;
32'hFFFF1EF8: romout <= 16'h0303;
32'hFFFF1EFA: romout <= 16'h66F6;
32'hFFFF1EFC: romout <= 16'h3039;
32'hFFFF1EFE: romout <= 16'hFFDC;
32'hFFFF1F00: romout <= 16'h0302;
32'hFFFF1F02: romout <= 16'h4E75;
32'hFFFF1F04: romout <= 16'h48E7;
32'hFFFF1F06: romout <= 16'hC044;
32'hFFFF1F08: romout <= 16'h2A7C;
32'hFFFF1F0A: romout <= 16'h0000;
32'hFFFF1F0C: romout <= 16'h0700;
32'hFFFF1F0E: romout <= 16'h2001;
32'hFFFF1F10: romout <= 16'h6100;
32'hFFFF1F12: romout <= 16'h122C;
32'hFFFF1F14: romout <= 16'h227C;
32'hFFFF1F16: romout <= 16'h0000;
32'hFFFF1F18: romout <= 16'h0700;
32'hFFFF1F1A: romout <= 16'h6100;
32'hFFFF1F1C: romout <= 16'hF93C;
32'hFFFF1F1E: romout <= 16'h4CDF;
32'hFFFF1F20: romout <= 16'h2203;
32'hFFFF1F22: romout <= 16'h4E75;
32'hFFFF1F24: romout <= 16'h48E7;
32'hFFFF1F26: romout <= 16'hB000;
32'hFFFF1F28: romout <= 16'h343C;
32'hFFFF1F2A: romout <= 16'h0007;
32'hFFFF1F2C: romout <= 16'h1001;
32'hFFFF1F2E: romout <= 16'h0240;
32'hFFFF1F30: romout <= 16'h000F;
32'hFFFF1F32: romout <= 16'h0C40;
32'hFFFF1F34: romout <= 16'h0009;
32'hFFFF1F36: romout <= 16'h6302;
32'hFFFF1F38: romout <= 16'h5E40;
32'hFFFF1F3A: romout <= 16'h0640;
32'hFFFF1F3C: romout <= 16'h0130;
32'hFFFF1F3E: romout <= 16'h3602;
32'hFFFF1F40: romout <= 16'hE343;
32'hFFFF1F42: romout <= 16'h3380;
32'hFFFF1F44: romout <= 16'h3000;
32'hFFFF1F46: romout <= 16'hE899;
32'hFFFF1F48: romout <= 16'h57CA;
32'hFFFF1F4A: romout <= 16'hFFE2;
32'hFFFF1F4C: romout <= 16'h4CDF;
32'hFFFF1F4E: romout <= 16'h000D;
32'hFFFF1F50: romout <= 16'h4E75;
32'hFFFF1F52: romout <= 16'h207C;
32'hFFFF1F54: romout <= 16'h0000;
32'hFFFF1F56: romout <= 16'h0008;
32'hFFFF1F58: romout <= 16'h203C;
32'hFFFF1F5A: romout <= 16'hAAAA;
32'hFFFF1F5C: romout <= 16'h5555;
32'hFFFF1F5E: romout <= 16'h43F9;
32'hFFFF1F60: romout <= 16'hFFD0;
32'hFFFF1F62: romout <= 16'h0014;
32'hFFFF1F64: romout <= 16'h2080;
32'hFFFF1F66: romout <= 16'hB098;
32'hFFFF1F68: romout <= 16'h6614;
32'hFFFF1F6A: romout <= 16'h2208;
32'hFFFF1F6C: romout <= 16'h4A41;
32'hFFFF1F6E: romout <= 16'h6606;
32'hFFFF1F70: romout <= 16'h4EB9;
32'hFFFF1F72: romout <= 16'hFFFF;
32'hFFFF1F74: romout <= 16'h1F24;
32'hFFFF1F76: romout <= 16'hB1FC;
32'hFFFF1F78: romout <= 16'h00FF;
32'hFFFF1F7A: romout <= 16'hFFFC;
32'hFFFF1F7C: romout <= 16'h65E6;
32'hFFFF1F7E: romout <= 16'h2448;
32'hFFFF1F80: romout <= 16'h207C;
32'hFFFF1F82: romout <= 16'h0000;
32'hFFFF1F84: romout <= 16'h0008;
32'hFFFF1F86: romout <= 16'h2018;
32'hFFFF1F88: romout <= 16'h2208;
32'hFFFF1F8A: romout <= 16'h4A41;
32'hFFFF1F8C: romout <= 16'h6606;
32'hFFFF1F8E: romout <= 16'h4EB9;
32'hFFFF1F90: romout <= 16'hFFFF;
32'hFFFF1F92: romout <= 16'h1F24;
32'hFFFF1F94: romout <= 16'h0C80;
32'hFFFF1F96: romout <= 16'hAAAA;
32'hFFFF1F98: romout <= 16'h5555;
32'hFFFF1F9A: romout <= 16'h67EA;
32'hFFFF1F9C: romout <= 16'hB5C8;
32'hFFFF1F9E: romout <= 16'h6668;
32'hFFFF1FA0: romout <= 16'h207C;
32'hFFFF1FA2: romout <= 16'h0000;
32'hFFFF1FA4: romout <= 16'h0008;
32'hFFFF1FA6: romout <= 16'h203C;
32'hFFFF1FA8: romout <= 16'h5555;
32'hFFFF1FAA: romout <= 16'hAAAA;
32'hFFFF1FAC: romout <= 16'h2080;
32'hFFFF1FAE: romout <= 16'hB098;
32'hFFFF1FB0: romout <= 16'h6614;
32'hFFFF1FB2: romout <= 16'h2208;
32'hFFFF1FB4: romout <= 16'h4A41;
32'hFFFF1FB6: romout <= 16'h6606;
32'hFFFF1FB8: romout <= 16'h4EB9;
32'hFFFF1FBA: romout <= 16'hFFFF;
32'hFFFF1FBC: romout <= 16'h1F24;
32'hFFFF1FBE: romout <= 16'hB1FC;
32'hFFFF1FC0: romout <= 16'h00FF;
32'hFFFF1FC2: romout <= 16'hFFFC;
32'hFFFF1FC4: romout <= 16'h65E6;
32'hFFFF1FC6: romout <= 16'h2448;
32'hFFFF1FC8: romout <= 16'h207C;
32'hFFFF1FCA: romout <= 16'h0000;
32'hFFFF1FCC: romout <= 16'h0008;
32'hFFFF1FCE: romout <= 16'h2018;
32'hFFFF1FD0: romout <= 16'h2208;
32'hFFFF1FD2: romout <= 16'h4A41;
32'hFFFF1FD4: romout <= 16'h6606;
32'hFFFF1FD6: romout <= 16'h4EB9;
32'hFFFF1FD8: romout <= 16'hFFFF;
32'hFFFF1FDA: romout <= 16'h1F24;
32'hFFFF1FDC: romout <= 16'h0C80;
32'hFFFF1FDE: romout <= 16'h5555;
32'hFFFF1FE0: romout <= 16'hAAAA;
32'hFFFF1FE2: romout <= 16'h67EA;
32'hFFFF1FE4: romout <= 16'hB5C8;
32'hFFFF1FE6: romout <= 16'h6620;
32'hFFFF1FE8: romout <= 16'h21C8;
32'hFFFF1FEA: romout <= 16'h0500;
32'hFFFF1FEC: romout <= 16'h91FC;
32'hFFFF1FEE: romout <= 16'h0000;
32'hFFFF1FF0: romout <= 16'h000C;
32'hFFFF1FF2: romout <= 16'h21C8;
32'hFFFF1FF4: romout <= 16'h0404;
32'hFFFF1FF6: romout <= 16'h21FC;
32'hFFFF1FF8: romout <= 16'h4652;
32'hFFFF1FFA: romout <= 16'h4545;
32'hFFFF1FFC: romout <= 16'h0400;
32'hFFFF1FFE: romout <= 16'h21FC;
32'hFFFF2000: romout <= 16'h0000;
32'hFFFF2002: romout <= 16'h0408;
32'hFFFF2004: romout <= 16'h0408;
32'hFFFF2006: romout <= 16'h4ED3;
32'hFFFF2008: romout <= 16'h4ED3;
32'hFFFF200A: romout <= 16'h60FC;
32'hFFFF200C: romout <= 16'h48E7;
32'hFFFF200E: romout <= 16'hF0C0;
32'hFFFF2010: romout <= 16'h43F9;
32'hFFFF2012: romout <= 16'hFFFF;
32'hFFFF2014: romout <= 16'h204E;
32'hFFFF2016: romout <= 16'h4EB9;
32'hFFFF2018: romout <= 16'hFFFF;
32'hFFFF201A: romout <= 16'h1858;
32'hFFFF201C: romout <= 16'h4CDF;
32'hFFFF201E: romout <= 16'h030F;
32'hFFFF2020: romout <= 16'h4E73;
32'hFFFF2022: romout <= 16'h48E7;
32'hFFFF2024: romout <= 16'hF0C0;
32'hFFFF2026: romout <= 16'h43F9;
32'hFFFF2028: romout <= 16'hFFFF;
32'hFFFF202A: romout <= 16'h205C;
32'hFFFF202C: romout <= 16'h4EB9;
32'hFFFF202E: romout <= 16'hFFFF;
32'hFFFF2030: romout <= 16'h1858;
32'hFFFF2032: romout <= 16'h4CDF;
32'hFFFF2034: romout <= 16'h030F;
32'hFFFF2036: romout <= 16'h4E73;
32'hFFFF2038: romout <= 16'h48E7;
32'hFFFF203A: romout <= 16'hF0C0;
32'hFFFF203C: romout <= 16'h43F9;
32'hFFFF203E: romout <= 16'hFFFF;
32'hFFFF2040: romout <= 16'h2066;
32'hFFFF2042: romout <= 16'h4EB9;
32'hFFFF2044: romout <= 16'hFFFF;
32'hFFFF2046: romout <= 16'h1858;
32'hFFFF2048: romout <= 16'h4CDF;
32'hFFFF204A: romout <= 16'h030F;
32'hFFFF204C: romout <= 16'h4E73;
32'hFFFF204E: romout <= 16'h4164;
32'hFFFF2050: romout <= 16'h6472;
32'hFFFF2052: romout <= 16'h6573;
32'hFFFF2054: romout <= 16'h7320;
32'hFFFF2056: romout <= 16'h6572;
32'hFFFF2058: romout <= 16'h726F;
32'hFFFF205A: romout <= 16'h7200;
32'hFFFF205C: romout <= 16'h4275;
32'hFFFF205E: romout <= 16'h7320;
32'hFFFF2060: romout <= 16'h6572;
32'hFFFF2062: romout <= 16'h726F;
32'hFFFF2064: romout <= 16'h7200;
32'hFFFF2066: romout <= 16'h496C;
32'hFFFF2068: romout <= 16'h6C65;
32'hFFFF206A: romout <= 16'h6761;
32'hFFFF206C: romout <= 16'h6C20;
32'hFFFF206E: romout <= 16'h696E;
32'hFFFF2070: romout <= 16'h7374;
32'hFFFF2072: romout <= 16'h7275;
32'hFFFF2074: romout <= 16'h6374;
32'hFFFF2076: romout <= 16'h696F;
32'hFFFF2078: romout <= 16'h6E00;
32'hFFFF207A: romout <= 16'h4469;
32'hFFFF207C: romout <= 16'h7669;
32'hFFFF207E: romout <= 16'h6465;
32'hFFFF2080: romout <= 16'h2062;
32'hFFFF2082: romout <= 16'h7920;
32'hFFFF2084: romout <= 16'h7A65;
32'hFFFF2086: romout <= 16'h726F;
32'hFFFF2400: romout <= 16'h6000;
32'hFFFF2402: romout <= 16'h0022;
32'hFFFF2404: romout <= 16'h6000;
32'hFFFF2406: romout <= 16'h005A;
32'hFFFF2408: romout <= 16'h6000;
32'hFFFF240A: romout <= 16'h0C96;
32'hFFFF240C: romout <= 16'h6000;
32'hFFFF240E: romout <= 16'h0CA4;
32'hFFFF2410: romout <= 16'h6000;
32'hFFFF2412: romout <= 16'h0CB8;
32'hFFFF2414: romout <= 16'h6000;
32'hFFFF2416: romout <= 16'h0CC6;
32'hFFFF2418: romout <= 16'h6000;
32'hFFFF241A: romout <= 16'h0CD8;
32'hFFFF241C: romout <= 16'h00C0;
32'hFFFF241E: romout <= 16'h0000;
32'hFFFF2420: romout <= 16'h00F0;
32'hFFFF2422: romout <= 16'h0000;
32'hFFFF2424: romout <= 16'h41F9;
32'hFFFF2426: romout <= 16'hFFFF;
32'hFFFF2428: romout <= 16'h2400;
32'hFFFF242A: romout <= 16'h21C8;
32'hFFFF242C: romout <= 16'h0600;
32'hFFFF242E: romout <= 16'h2E79;
32'hFFFF2430: romout <= 16'hFFFF;
32'hFFFF2432: romout <= 16'h2420;
32'hFFFF2434: romout <= 16'h4DF9;
32'hFFFF2436: romout <= 16'hFFFF;
32'hFFFF2438: romout <= 16'h30F8;
32'hFFFF243A: romout <= 16'h6100;
32'hFFFF243C: romout <= 16'h0C58;
32'hFFFF243E: romout <= 16'h21F9;
32'hFFFF2440: romout <= 16'hFFFF;
32'hFFFF2442: romout <= 16'h241C;
32'hFFFF2444: romout <= 16'h0624;
32'hFFFF2446: romout <= 16'h2039;
32'hFFFF2448: romout <= 16'hFFFF;
32'hFFFF244A: romout <= 16'h2420;
32'hFFFF244C: romout <= 16'h0480;
32'hFFFF244E: romout <= 16'h0000;
32'hFFFF2450: romout <= 16'h0800;
32'hFFFF2452: romout <= 16'h21C0;
32'hFFFF2454: romout <= 16'h062C;
32'hFFFF2456: romout <= 16'h0480;
32'hFFFF2458: romout <= 16'h0000;
32'hFFFF245A: romout <= 16'h1008;
32'hFFFF245C: romout <= 16'h21C0;
32'hFFFF245E: romout <= 16'h0628;
32'hFFFF2460: romout <= 16'h4280;
32'hFFFF2462: romout <= 16'h21C0;
32'hFFFF2464: romout <= 16'h0610;
32'hFFFF2466: romout <= 16'h21C0;
32'hFFFF2468: romout <= 16'h0608;
32'hFFFF246A: romout <= 16'h21C0;
32'hFFFF246C: romout <= 16'h0604;
32'hFFFF246E: romout <= 16'h2E79;
32'hFFFF2470: romout <= 16'hFFFF;
32'hFFFF2472: romout <= 16'h2420;
32'hFFFF2474: romout <= 16'h4DF9;
32'hFFFF2476: romout <= 16'hFFFF;
32'hFFFF2478: romout <= 16'h311E;
32'hFFFF247A: romout <= 16'h6100;
32'hFFFF247C: romout <= 16'h0C18;
32'hFFFF247E: romout <= 16'h103C;
32'hFFFF2480: romout <= 16'h003E;
32'hFFFF2482: romout <= 16'h6100;
32'hFFFF2484: romout <= 16'h0976;
32'hFFFF2486: romout <= 16'h6100;
32'hFFFF2488: romout <= 16'h0BA8;
32'hFFFF248A: romout <= 16'h2848;
32'hFFFF248C: romout <= 16'h41F8;
32'hFFFF248E: romout <= 16'h0630;
32'hFFFF2490: romout <= 16'h6100;
32'hFFFF2492: romout <= 16'h0B5A;
32'hFFFF2494: romout <= 16'h6100;
32'hFFFF2496: romout <= 16'h0B8E;
32'hFFFF2498: romout <= 16'h4A81;
32'hFFFF249A: romout <= 16'h6700;
32'hFFFF249C: romout <= 16'h0152;
32'hFFFF249E: romout <= 16'hB2BC;
32'hFFFF24A0: romout <= 16'h0000;
32'hFFFF24A2: romout <= 16'hFFFF;
32'hFFFF24A4: romout <= 16'h6400;
32'hFFFF24A6: romout <= 16'h094A;
32'hFFFF24A8: romout <= 16'h1101;
32'hFFFF24AA: romout <= 16'hE099;
32'hFFFF24AC: romout <= 16'h1101;
32'hFFFF24AE: romout <= 16'hE199;
32'hFFFF24B0: romout <= 16'h6100;
32'hFFFF24B2: romout <= 16'h09E8;
32'hFFFF24B4: romout <= 16'h2A49;
32'hFFFF24B6: romout <= 16'h6612;
32'hFFFF24B8: romout <= 16'h6100;
32'hFFFF24BA: romout <= 16'h0A08;
32'hFFFF24BC: romout <= 16'h244D;
32'hFFFF24BE: romout <= 16'h2678;
32'hFFFF24C0: romout <= 16'h0624;
32'hFFFF24C2: romout <= 16'h6100;
32'hFFFF24C4: romout <= 16'h0A08;
32'hFFFF24C6: romout <= 16'h21CA;
32'hFFFF24C8: romout <= 16'h0624;
32'hFFFF24CA: romout <= 16'h200C;
32'hFFFF24CC: romout <= 16'h9088;
32'hFFFF24CE: romout <= 16'hB0BC;
32'hFFFF24D0: romout <= 16'h0000;
32'hFFFF24D2: romout <= 16'h0003;
32'hFFFF24D4: romout <= 16'h67A8;
32'hFFFF24D6: romout <= 16'h2678;
32'hFFFF24D8: romout <= 16'h0624;
32'hFFFF24DA: romout <= 16'h2C4B;
32'hFFFF24DC: romout <= 16'hD7C0;
32'hFFFF24DE: romout <= 16'h2038;
32'hFFFF24E0: romout <= 16'h0628;
32'hFFFF24E2: romout <= 16'hB08B;
32'hFFFF24E4: romout <= 16'h6300;
32'hFFFF24E6: romout <= 16'h0900;
32'hFFFF24E8: romout <= 16'h21CB;
32'hFFFF24EA: romout <= 16'h0624;
32'hFFFF24EC: romout <= 16'h224E;
32'hFFFF24EE: romout <= 16'h244D;
32'hFFFF24F0: romout <= 16'h6100;
32'hFFFF24F2: romout <= 16'h09E4;
32'hFFFF24F4: romout <= 16'h2248;
32'hFFFF24F6: romout <= 16'h244D;
32'hFFFF24F8: romout <= 16'h264C;
32'hFFFF24FA: romout <= 16'h6100;
32'hFFFF24FC: romout <= 16'h09D0;
32'hFFFF24FE: romout <= 16'h6000;
32'hFFFF2500: romout <= 16'hFF7E;
32'hFFFF2502: romout <= 16'h4C49;
32'hFFFF2504: romout <= 16'h53D4;
32'hFFFF2506: romout <= 16'h4C4F;
32'hFFFF2508: romout <= 16'h41C4;
32'hFFFF250A: romout <= 16'h4E45;
32'hFFFF250C: romout <= 16'hD752;
32'hFFFF250E: romout <= 16'h55CE;
32'hFFFF2510: romout <= 16'h5341;
32'hFFFF2512: romout <= 16'h56C5;
32'hFFFF2514: romout <= 16'h434C;
32'hFFFF2516: romout <= 16'hD34E;
32'hFFFF2518: romout <= 16'h4558;
32'hFFFF251A: romout <= 16'hD44C;
32'hFFFF251C: romout <= 16'h45D4;
32'hFFFF251E: romout <= 16'h49C6;
32'hFFFF2520: romout <= 16'h474F;
32'hFFFF2522: romout <= 16'h54CF;
32'hFFFF2524: romout <= 16'h474F;
32'hFFFF2526: romout <= 16'h5355;
32'hFFFF2528: romout <= 16'hC252;
32'hFFFF252A: romout <= 16'h4554;
32'hFFFF252C: romout <= 16'h5552;
32'hFFFF252E: romout <= 16'hCE52;
32'hFFFF2530: romout <= 16'h45CD;
32'hFFFF2532: romout <= 16'h464F;
32'hFFFF2534: romout <= 16'hD249;
32'hFFFF2536: romout <= 16'h4E50;
32'hFFFF2538: romout <= 16'h55D4;
32'hFFFF253A: romout <= 16'h5052;
32'hFFFF253C: romout <= 16'h494E;
32'hFFFF253E: romout <= 16'hD450;
32'hFFFF2540: romout <= 16'h4F4B;
32'hFFFF2542: romout <= 16'hC553;
32'hFFFF2544: romout <= 16'h544F;
32'hFFFF2546: romout <= 16'hD042;
32'hFFFF2548: romout <= 16'h59C5;
32'hFFFF254A: romout <= 16'h4341;
32'hFFFF254C: romout <= 16'h4CCC;
32'hFFFF254E: romout <= 16'h4C49;
32'hFFFF2550: romout <= 16'h4EC5;
32'hFFFF2552: romout <= 16'h504F;
32'hFFFF2554: romout <= 16'h494E;
32'hFFFF2556: romout <= 16'hD450;
32'hFFFF2558: romout <= 16'h454E;
32'hFFFF255A: romout <= 16'h434F;
32'hFFFF255C: romout <= 16'h4C4F;
32'hFFFF255E: romout <= 16'hD246;
32'hFFFF2560: romout <= 16'h494C;
32'hFFFF2562: romout <= 16'h4C43;
32'hFFFF2564: romout <= 16'h4F4C;
32'hFFFF2566: romout <= 16'h4FD2;
32'hFFFF2568: romout <= 16'h0050;
32'hFFFF256A: romout <= 16'h4545;
32'hFFFF256C: romout <= 16'hCB52;
32'hFFFF256E: romout <= 16'h4EC4;
32'hFFFF2570: romout <= 16'h4142;
32'hFFFF2572: romout <= 16'hD353;
32'hFFFF2574: romout <= 16'h495A;
32'hFFFF2576: romout <= 16'hC554;
32'hFFFF2578: romout <= 16'h4943;
32'hFFFF257A: romout <= 16'hCB54;
32'hFFFF257C: romout <= 16'h454D;
32'hFFFF257E: romout <= 16'hD053;
32'hFFFF2580: romout <= 16'h47CE;
32'hFFFF2582: romout <= 16'h0054;
32'hFFFF2584: romout <= 16'hCF00;
32'hFFFF2586: romout <= 16'h5354;
32'hFFFF2588: romout <= 16'h45D0;
32'hFFFF258A: romout <= 16'h003E;
32'hFFFF258C: romout <= 16'hBD3C;
32'hFFFF258E: romout <= 16'hBEBE;
32'hFFFF2590: romout <= 16'hBD3C;
32'hFFFF2592: romout <= 16'hBDBC;
32'hFFFF2594: romout <= 16'h00FF;
32'hFFFF2596: romout <= 16'h26B4;
32'hFFFF2598: romout <= 16'h28F6;
32'hFFFF259A: romout <= 16'h264E;
32'hFFFF259C: romout <= 16'h2662;
32'hFFFF259E: romout <= 16'h295A;
32'hFFFF25A0: romout <= 16'h263C;
32'hFFFF25A2: romout <= 16'h2802;
32'hFFFF25A4: romout <= 16'h28E6;
32'hFFFF25A6: romout <= 16'h2852;
32'hFFFF25A8: romout <= 16'h26A0;
32'hFFFF25AA: romout <= 16'h274A;
32'hFFFF25AC: romout <= 16'h2772;
32'hFFFF25AE: romout <= 16'h2850;
32'hFFFF25B0: romout <= 16'h2790;
32'hFFFF25B2: romout <= 16'h2878;
32'hFFFF25B4: romout <= 16'h26E0;
32'hFFFF25B6: romout <= 16'h29DE;
32'hFFFF25B8: romout <= 16'h265A;
32'hFFFF25BA: romout <= 16'h2418;
32'hFFFF25BC: romout <= 16'h2A94;
32'hFFFF25BE: romout <= 16'h2A32;
32'hFFFF25C0: romout <= 16'h29FA;
32'hFFFF25C2: romout <= 16'h2A16;
32'hFFFF25C4: romout <= 16'h2A24;
32'hFFFF25C6: romout <= 16'h28E0;
32'hFFFF25C8: romout <= 16'h2CEE;
32'hFFFF25CA: romout <= 16'h2CFA;
32'hFFFF25CC: romout <= 16'h2D26;
32'hFFFF25CE: romout <= 16'h2D48;
32'hFFFF25D0: romout <= 16'h2D52;
32'hFFFF25D2: romout <= 16'h2D58;
32'hFFFF25D4: romout <= 16'h2D36;
32'hFFFF25D6: romout <= 16'h2BC8;
32'hFFFF25D8: romout <= 16'h27AC;
32'hFFFF25DA: romout <= 16'h2DA4;
32'hFFFF25DC: romout <= 16'h27C4;
32'hFFFF25DE: romout <= 16'h27CA;
32'hFFFF25E0: romout <= 16'h2AC0;
32'hFFFF25E2: romout <= 16'h2AC8;
32'hFFFF25E4: romout <= 16'h2AD0;
32'hFFFF25E6: romout <= 16'h2AE0;
32'hFFFF25E8: romout <= 16'h2AD8;
32'hFFFF25EA: romout <= 16'h2AEA;
32'hFFFF25EC: romout <= 16'h2AFC;
32'hFFFF25EE: romout <= 16'h43F9;
32'hFFFF25F0: romout <= 16'hFFFF;
32'hFFFF25F2: romout <= 16'h2502;
32'hFFFF25F4: romout <= 16'h45F9;
32'hFFFF25F6: romout <= 16'hFFFF;
32'hFFFF25F8: romout <= 16'h2596;
32'hFFFF25FA: romout <= 16'h6100;
32'hFFFF25FC: romout <= 16'h0A28;
32'hFFFF25FE: romout <= 16'h2648;
32'hFFFF2600: romout <= 16'h4202;
32'hFFFF2602: romout <= 16'h1018;
32'hFFFF2604: romout <= 16'h1211;
32'hFFFF2606: romout <= 16'h6604;
32'hFFFF2608: romout <= 16'h204B;
32'hFFFF260A: romout <= 16'h6024;
32'hFFFF260C: romout <= 16'h1600;
32'hFFFF260E: romout <= 16'hC602;
32'hFFFF2610: romout <= 16'hB63C;
32'hFFFF2612: romout <= 16'h002E;
32'hFFFF2614: romout <= 16'h671A;
32'hFFFF2616: romout <= 16'h0201;
32'hFFFF2618: romout <= 16'h007F;
32'hFFFF261A: romout <= 16'hB200;
32'hFFFF261C: romout <= 16'h670C;
32'hFFFF261E: romout <= 16'h548A;
32'hFFFF2620: romout <= 16'h204B;
32'hFFFF2622: romout <= 16'h4202;
32'hFFFF2624: romout <= 16'h4A19;
32'hFFFF2626: romout <= 16'h6AFC;
32'hFFFF2628: romout <= 16'h60D8;
32'hFFFF262A: romout <= 16'h74FF;
32'hFFFF262C: romout <= 16'h4A19;
32'hFFFF262E: romout <= 16'h6AD2;
32'hFFFF2630: romout <= 16'h47F9;
32'hFFFF2632: romout <= 16'hFFFF;
32'hFFFF2634: romout <= 16'h0000;
32'hFFFF2636: romout <= 16'h3452;
32'hFFFF2638: romout <= 16'h4EF3;
32'hFFFF263A: romout <= 16'hA000;
32'hFFFF263C: romout <= 16'h4EB9;
32'hFFFF263E: romout <= 16'hFFFF;
32'hFFFF2640: romout <= 16'h18E8;
32'hFFFF2642: romout <= 16'h4278;
32'hFFFF2644: romout <= 16'h0418;
32'hFFFF2646: romout <= 16'h4278;
32'hFFFF2648: romout <= 16'h041A;
32'hFFFF264A: romout <= 16'h6000;
32'hFFFF264C: romout <= 16'hFE14;
32'hFFFF264E: romout <= 16'h6100;
32'hFFFF2650: romout <= 16'h0748;
32'hFFFF2652: romout <= 16'h21F9;
32'hFFFF2654: romout <= 16'hFFFF;
32'hFFFF2656: romout <= 16'h241C;
32'hFFFF2658: romout <= 16'h0624;
32'hFFFF265A: romout <= 16'h6100;
32'hFFFF265C: romout <= 16'h073C;
32'hFFFF265E: romout <= 16'h6000;
32'hFFFF2660: romout <= 16'hFE00;
32'hFFFF2662: romout <= 16'h6100;
32'hFFFF2664: romout <= 16'h0734;
32'hFFFF2666: romout <= 16'h2079;
32'hFFFF2668: romout <= 16'hFFFF;
32'hFFFF266A: romout <= 16'h241C;
32'hFFFF266C: romout <= 16'h21C8;
32'hFFFF266E: romout <= 16'h0604;
32'hFFFF2670: romout <= 16'h4AB8;
32'hFFFF2672: romout <= 16'h0604;
32'hFFFF2674: romout <= 16'h6700;
32'hFFFF2676: romout <= 16'hFDEA;
32'hFFFF2678: romout <= 16'h4281;
32'hFFFF267A: romout <= 16'h2248;
32'hFFFF267C: romout <= 16'h6100;
32'hFFFF267E: romout <= 16'h082C;
32'hFFFF2680: romout <= 16'h6500;
32'hFFFF2682: romout <= 16'hFDDE;
32'hFFFF2684: romout <= 16'h21C9;
32'hFFFF2686: romout <= 16'h0604;
32'hFFFF2688: romout <= 16'h2049;
32'hFFFF268A: romout <= 16'h5488;
32'hFFFF268C: romout <= 16'h6100;
32'hFFFF268E: romout <= 16'h09EE;
32'hFFFF2690: romout <= 16'h43F9;
32'hFFFF2692: romout <= 16'hFFFF;
32'hFFFF2694: romout <= 16'h2517;
32'hFFFF2696: romout <= 16'h45F9;
32'hFFFF2698: romout <= 16'hFFFF;
32'hFFFF269A: romout <= 16'h25A2;
32'hFFFF269C: romout <= 16'h6000;
32'hFFFF269E: romout <= 16'hFF5C;
32'hFFFF26A0: romout <= 16'h6100;
32'hFFFF26A2: romout <= 16'h0408;
32'hFFFF26A4: romout <= 16'h6100;
32'hFFFF26A6: romout <= 16'h06F2;
32'hFFFF26A8: romout <= 16'h2200;
32'hFFFF26AA: romout <= 16'h6100;
32'hFFFF26AC: romout <= 16'h07EE;
32'hFFFF26AE: romout <= 16'h6600;
32'hFFFF26B0: romout <= 16'h0740;
32'hFFFF26B2: romout <= 16'h60D0;
32'hFFFF26B4: romout <= 16'h6100;
32'hFFFF26B6: romout <= 16'h0936;
32'hFFFF26B8: romout <= 16'h6100;
32'hFFFF26BA: romout <= 16'h06DE;
32'hFFFF26BC: romout <= 16'h6100;
32'hFFFF26BE: romout <= 16'h07DC;
32'hFFFF26C0: romout <= 16'h6500;
32'hFFFF26C2: romout <= 16'hFD9E;
32'hFFFF26C4: romout <= 16'h6100;
32'hFFFF26C6: romout <= 16'h08F0;
32'hFFFF26C8: romout <= 16'h6100;
32'hFFFF26CA: romout <= 16'h09B2;
32'hFFFF26CC: romout <= 16'h670C;
32'hFFFF26CE: romout <= 16'hB03C;
32'hFFFF26D0: romout <= 16'h0013;
32'hFFFF26D2: romout <= 16'h6606;
32'hFFFF26D4: romout <= 16'h6100;
32'hFFFF26D6: romout <= 16'h09A6;
32'hFFFF26D8: romout <= 16'h67FA;
32'hFFFF26DA: romout <= 16'h6100;
32'hFFFF26DC: romout <= 16'h07CE;
32'hFFFF26DE: romout <= 16'h60E0;
32'hFFFF26E0: romout <= 16'h780B;
32'hFFFF26E2: romout <= 16'h6100;
32'hFFFF26E4: romout <= 16'h08EE;
32'hFFFF26E6: romout <= 16'h3A07;
32'hFFFF26E8: romout <= 16'h6100;
32'hFFFF26EA: romout <= 16'h09A4;
32'hFFFF26EC: romout <= 16'h609E;
32'hFFFF26EE: romout <= 16'h6100;
32'hFFFF26F0: romout <= 16'h08E2;
32'hFFFF26F2: romout <= 16'h0D09;
32'hFFFF26F4: romout <= 16'h6100;
32'hFFFF26F6: romout <= 16'h0998;
32'hFFFF26F8: romout <= 16'h6000;
32'hFFFF26FA: romout <= 16'hFF76;
32'hFFFF26FC: romout <= 16'h6100;
32'hFFFF26FE: romout <= 16'h08D4;
32'hFFFF2700: romout <= 16'h2309;
32'hFFFF2702: romout <= 16'h6100;
32'hFFFF2704: romout <= 16'h03A6;
32'hFFFF2706: romout <= 16'h2800;
32'hFFFF2708: romout <= 16'h6016;
32'hFFFF270A: romout <= 16'h6100;
32'hFFFF270C: romout <= 16'h08C6;
32'hFFFF270E: romout <= 16'h240B;
32'hFFFF2710: romout <= 16'h6100;
32'hFFFF2712: romout <= 16'h0398;
32'hFFFF2714: romout <= 16'h6100;
32'hFFFF2716: romout <= 16'hFCF2;
32'hFFFF2718: romout <= 16'h6006;
32'hFFFF271A: romout <= 16'h6100;
32'hFFFF271C: romout <= 16'h081E;
32'hFFFF271E: romout <= 16'h6012;
32'hFFFF2720: romout <= 16'h6100;
32'hFFFF2722: romout <= 16'h08B0;
32'hFFFF2724: romout <= 16'h2C07;
32'hFFFF2726: romout <= 16'h6100;
32'hFFFF2728: romout <= 16'h0656;
32'hFFFF272A: romout <= 16'h60D0;
32'hFFFF272C: romout <= 16'h6100;
32'hFFFF272E: romout <= 16'h0960;
32'hFFFF2730: romout <= 16'h6010;
32'hFFFF2732: romout <= 16'h2F04;
32'hFFFF2734: romout <= 16'h6100;
32'hFFFF2736: romout <= 16'h0374;
32'hFFFF2738: romout <= 16'h281F;
32'hFFFF273A: romout <= 16'h2200;
32'hFFFF273C: romout <= 16'h6100;
32'hFFFF273E: romout <= 16'h083C;
32'hFFFF2740: romout <= 16'h60DE;
32'hFFFF2742: romout <= 16'h6100;
32'hFFFF2744: romout <= 16'h063A;
32'hFFFF2746: romout <= 16'h6000;
32'hFFFF2748: romout <= 16'h065C;
32'hFFFF274A: romout <= 16'h6100;
32'hFFFF274C: romout <= 16'h07AC;
32'hFFFF274E: romout <= 16'h6100;
32'hFFFF2750: romout <= 16'h035A;
32'hFFFF2752: romout <= 16'h2F08;
32'hFFFF2754: romout <= 16'h2200;
32'hFFFF2756: romout <= 16'h6100;
32'hFFFF2758: romout <= 16'h0742;
32'hFFFF275A: romout <= 16'h6600;
32'hFFFF275C: romout <= 16'h0696;
32'hFFFF275E: romout <= 16'h2F38;
32'hFFFF2760: romout <= 16'h0604;
32'hFFFF2762: romout <= 16'h2F38;
32'hFFFF2764: romout <= 16'h0608;
32'hFFFF2766: romout <= 16'h42B8;
32'hFFFF2768: romout <= 16'h0610;
32'hFFFF276A: romout <= 16'h21CF;
32'hFFFF276C: romout <= 16'h0608;
32'hFFFF276E: romout <= 16'h6000;
32'hFFFF2770: romout <= 16'hFF14;
32'hFFFF2772: romout <= 16'h6100;
32'hFFFF2774: romout <= 16'h0624;
32'hFFFF2776: romout <= 16'h2238;
32'hFFFF2778: romout <= 16'h0608;
32'hFFFF277A: romout <= 16'h6700;
32'hFFFF277C: romout <= 16'h0628;
32'hFFFF277E: romout <= 16'h2E41;
32'hFFFF2780: romout <= 16'h21DF;
32'hFFFF2782: romout <= 16'h0608;
32'hFFFF2784: romout <= 16'h21DF;
32'hFFFF2786: romout <= 16'h0604;
32'hFFFF2788: romout <= 16'h205F;
32'hFFFF278A: romout <= 16'h6100;
32'hFFFF278C: romout <= 16'h0752;
32'hFFFF278E: romout <= 16'h60B2;
32'hFFFF2790: romout <= 16'h6100;
32'hFFFF2792: romout <= 16'h0766;
32'hFFFF2794: romout <= 16'h6100;
32'hFFFF2796: romout <= 16'h05CE;
32'hFFFF2798: romout <= 16'h21CE;
32'hFFFF279A: romout <= 16'h0610;
32'hFFFF279C: romout <= 16'h43F9;
32'hFFFF279E: romout <= 16'hFFFF;
32'hFFFF27A0: romout <= 16'h2583;
32'hFFFF27A2: romout <= 16'h45F9;
32'hFFFF27A4: romout <= 16'hFFFF;
32'hFFFF27A6: romout <= 16'h25D8;
32'hFFFF27A8: romout <= 16'h6000;
32'hFFFF27AA: romout <= 16'hFE50;
32'hFFFF27AC: romout <= 16'h6100;
32'hFFFF27AE: romout <= 16'h02FC;
32'hFFFF27B0: romout <= 16'h21C0;
32'hFFFF27B2: romout <= 16'h0618;
32'hFFFF27B4: romout <= 16'h43F9;
32'hFFFF27B6: romout <= 16'hFFFF;
32'hFFFF27B8: romout <= 16'h2586;
32'hFFFF27BA: romout <= 16'h45F9;
32'hFFFF27BC: romout <= 16'hFFFF;
32'hFFFF27BE: romout <= 16'h25DC;
32'hFFFF27C0: romout <= 16'h6000;
32'hFFFF27C2: romout <= 16'hFE38;
32'hFFFF27C4: romout <= 16'h6100;
32'hFFFF27C6: romout <= 16'h02E4;
32'hFFFF27C8: romout <= 16'h6002;
32'hFFFF27CA: romout <= 16'h7001;
32'hFFFF27CC: romout <= 16'h21C0;
32'hFFFF27CE: romout <= 16'h0614;
32'hFFFF27D0: romout <= 16'h21F8;
32'hFFFF27D2: romout <= 16'h0604;
32'hFFFF27D4: romout <= 16'h061C;
32'hFFFF27D6: romout <= 16'h21C8;
32'hFFFF27D8: romout <= 16'h0620;
32'hFFFF27DA: romout <= 16'h2C4F;
32'hFFFF27DC: romout <= 16'h6006;
32'hFFFF27DE: romout <= 16'hDDFC;
32'hFFFF27E0: romout <= 16'h0000;
32'hFFFF27E2: romout <= 16'h0014;
32'hFFFF27E4: romout <= 16'h2016;
32'hFFFF27E6: romout <= 16'h6716;
32'hFFFF27E8: romout <= 16'hB0B8;
32'hFFFF27EA: romout <= 16'h0610;
32'hFFFF27EC: romout <= 16'h66F0;
32'hFFFF27EE: romout <= 16'h244F;
32'hFFFF27F0: romout <= 16'h224E;
32'hFFFF27F2: romout <= 16'h47F8;
32'hFFFF27F4: romout <= 16'h0014;
32'hFFFF27F6: romout <= 16'hD7C9;
32'hFFFF27F8: romout <= 16'h6100;
32'hFFFF27FA: romout <= 16'h06DC;
32'hFFFF27FC: romout <= 16'h2E4B;
32'hFFFF27FE: romout <= 16'h6000;
32'hFFFF2800: romout <= 16'hFF42;
32'hFFFF2802: romout <= 16'h6100;
32'hFFFF2804: romout <= 16'h03F2;
32'hFFFF2806: romout <= 16'h6500;
32'hFFFF2808: romout <= 16'h059C;
32'hFFFF280A: romout <= 16'h2240;
32'hFFFF280C: romout <= 16'h2038;
32'hFFFF280E: romout <= 16'h0610;
32'hFFFF2810: romout <= 16'h6700;
32'hFFFF2812: romout <= 16'h0592;
32'hFFFF2814: romout <= 16'hB3C0;
32'hFFFF2816: romout <= 16'h6706;
32'hFFFF2818: romout <= 16'h6100;
32'hFFFF281A: romout <= 16'h06C4;
32'hFFFF281C: romout <= 16'h60EE;
32'hFFFF281E: romout <= 16'h2011;
32'hFFFF2820: romout <= 16'hD0B8;
32'hFFFF2822: romout <= 16'h0614;
32'hFFFF2824: romout <= 16'h6900;
32'hFFFF2826: romout <= 16'h05CA;
32'hFFFF2828: romout <= 16'h2280;
32'hFFFF282A: romout <= 16'h2238;
32'hFFFF282C: romout <= 16'h0618;
32'hFFFF282E: romout <= 16'h4AB8;
32'hFFFF2830: romout <= 16'h0614;
32'hFFFF2832: romout <= 16'h6A02;
32'hFFFF2834: romout <= 16'hC141;
32'hFFFF2836: romout <= 16'hB280;
32'hFFFF2838: romout <= 16'h6D0E;
32'hFFFF283A: romout <= 16'h21F8;
32'hFFFF283C: romout <= 16'h061C;
32'hFFFF283E: romout <= 16'h0604;
32'hFFFF2840: romout <= 16'h2078;
32'hFFFF2842: romout <= 16'h0620;
32'hFFFF2844: romout <= 16'h6000;
32'hFFFF2846: romout <= 16'hFEFC;
32'hFFFF2848: romout <= 16'h6100;
32'hFFFF284A: romout <= 16'h0694;
32'hFFFF284C: romout <= 16'h6000;
32'hFFFF284E: romout <= 16'hFEF4;
32'hFFFF2850: romout <= 16'h600A;
32'hFFFF2852: romout <= 16'h6100;
32'hFFFF2854: romout <= 16'h0256;
32'hFFFF2856: romout <= 16'h4A80;
32'hFFFF2858: romout <= 16'h6600;
32'hFFFF285A: romout <= 16'hFE32;
32'hFFFF285C: romout <= 16'h2248;
32'hFFFF285E: romout <= 16'h4281;
32'hFFFF2860: romout <= 16'h6100;
32'hFFFF2862: romout <= 16'h0662;
32'hFFFF2864: romout <= 16'h6400;
32'hFFFF2866: romout <= 16'hFE1E;
32'hFFFF2868: romout <= 16'h6000;
32'hFFFF286A: romout <= 16'hFBF6;
32'hFFFF286C: romout <= 16'h2E78;
32'hFFFF286E: romout <= 16'h060C;
32'hFFFF2870: romout <= 16'h21DF;
32'hFFFF2872: romout <= 16'h0604;
32'hFFFF2874: romout <= 16'h588F;
32'hFFFF2876: romout <= 16'h205F;
32'hFFFF2878: romout <= 16'h2F08;
32'hFFFF287A: romout <= 16'h6100;
32'hFFFF287C: romout <= 16'h06BE;
32'hFFFF287E: romout <= 16'h600A;
32'hFFFF2880: romout <= 16'h6100;
32'hFFFF2882: romout <= 16'h0374;
32'hFFFF2884: romout <= 16'h654C;
32'hFFFF2886: romout <= 16'h2440;
32'hFFFF2888: romout <= 16'h601A;
32'hFFFF288A: romout <= 16'h2F08;
32'hFFFF288C: romout <= 16'h6100;
32'hFFFF288E: romout <= 16'h0368;
32'hFFFF2890: romout <= 16'h6500;
32'hFFFF2892: romout <= 16'h0512;
32'hFFFF2894: romout <= 16'h2440;
32'hFFFF2896: romout <= 16'h1410;
32'hFFFF2898: romout <= 16'h4200;
32'hFFFF289A: romout <= 16'h1080;
32'hFFFF289C: romout <= 16'h225F;
32'hFFFF289E: romout <= 16'h6100;
32'hFFFF28A0: romout <= 16'h067E;
32'hFFFF28A2: romout <= 16'h1082;
32'hFFFF28A4: romout <= 16'h2F08;
32'hFFFF28A6: romout <= 16'h2F38;
32'hFFFF28A8: romout <= 16'h0604;
32'hFFFF28AA: romout <= 16'h21FC;
32'hFFFF28AC: romout <= 16'hFFFF;
32'hFFFF28AE: romout <= 16'hFFFF;
32'hFFFF28B0: romout <= 16'h0604;
32'hFFFF28B2: romout <= 16'h21CF;
32'hFFFF28B4: romout <= 16'h060C;
32'hFFFF28B6: romout <= 16'h2F0A;
32'hFFFF28B8: romout <= 16'h103C;
32'hFFFF28BA: romout <= 16'h003A;
32'hFFFF28BC: romout <= 16'h6100;
32'hFFFF28BE: romout <= 16'h053C;
32'hFFFF28C0: romout <= 16'h41F8;
32'hFFFF28C2: romout <= 16'h0630;
32'hFFFF28C4: romout <= 16'h6100;
32'hFFFF28C6: romout <= 16'h01E4;
32'hFFFF28C8: romout <= 16'h245F;
32'hFFFF28CA: romout <= 16'h2480;
32'hFFFF28CC: romout <= 16'h21DF;
32'hFFFF28CE: romout <= 16'h0604;
32'hFFFF28D0: romout <= 16'h205F;
32'hFFFF28D2: romout <= 16'h588F;
32'hFFFF28D4: romout <= 16'h6100;
32'hFFFF28D6: romout <= 16'h06FC;
32'hFFFF28D8: romout <= 16'h2C03;
32'hFFFF28DA: romout <= 16'h609C;
32'hFFFF28DC: romout <= 16'h6000;
32'hFFFF28DE: romout <= 16'hFE64;
32'hFFFF28E0: romout <= 16'h0C10;
32'hFFFF28E2: romout <= 16'h000D;
32'hFFFF28E4: romout <= 16'h670C;
32'hFFFF28E6: romout <= 16'h6100;
32'hFFFF28E8: romout <= 16'h047C;
32'hFFFF28EA: romout <= 16'h6100;
32'hFFFF28EC: romout <= 16'h06E6;
32'hFFFF28EE: romout <= 16'h2C03;
32'hFFFF28F0: romout <= 16'h60F4;
32'hFFFF28F2: romout <= 16'h6000;
32'hFFFF28F4: romout <= 16'hFE4E;
32'hFFFF28F6: romout <= 16'h2079;
32'hFFFF28F8: romout <= 16'hFFFF;
32'hFFFF28FA: romout <= 16'h241C;
32'hFFFF28FC: romout <= 16'h103C;
32'hFFFF28FE: romout <= 16'h000D;
32'hFFFF2900: romout <= 16'h6100;
32'hFFFF2902: romout <= 16'hFB0E;
32'hFFFF2904: romout <= 16'h6100;
32'hFFFF2906: romout <= 16'hFB0E;
32'hFFFF2908: romout <= 16'h67FA;
32'hFFFF290A: romout <= 16'hB03C;
32'hFFFF290C: romout <= 16'h0040;
32'hFFFF290E: romout <= 16'h6722;
32'hFFFF2910: romout <= 16'hB03C;
32'hFFFF2912: romout <= 16'h003A;
32'hFFFF2914: romout <= 16'h66EE;
32'hFFFF2916: romout <= 16'h6100;
32'hFFFF2918: romout <= 16'h0022;
32'hFFFF291A: romout <= 16'h10C1;
32'hFFFF291C: romout <= 16'h6100;
32'hFFFF291E: romout <= 16'h001C;
32'hFFFF2920: romout <= 16'h10C1;
32'hFFFF2922: romout <= 16'h6100;
32'hFFFF2924: romout <= 16'hFAF0;
32'hFFFF2926: romout <= 16'h67FA;
32'hFFFF2928: romout <= 16'h10C0;
32'hFFFF292A: romout <= 16'hB03C;
32'hFFFF292C: romout <= 16'h000D;
32'hFFFF292E: romout <= 16'h66F2;
32'hFFFF2930: romout <= 16'h60D2;
32'hFFFF2932: romout <= 16'h21C8;
32'hFFFF2934: romout <= 16'h0624;
32'hFFFF2936: romout <= 16'h6000;
32'hFFFF2938: romout <= 16'hFB28;
32'hFFFF293A: romout <= 16'h7401;
32'hFFFF293C: romout <= 16'h4281;
32'hFFFF293E: romout <= 16'h6100;
32'hFFFF2940: romout <= 16'hFAD4;
32'hFFFF2942: romout <= 16'h67FA;
32'hFFFF2944: romout <= 16'hB03C;
32'hFFFF2946: romout <= 16'h0041;
32'hFFFF2948: romout <= 16'h6502;
32'hFFFF294A: romout <= 16'h5F00;
32'hFFFF294C: romout <= 16'h0200;
32'hFFFF294E: romout <= 16'h000F;
32'hFFFF2950: romout <= 16'hE909;
32'hFFFF2952: romout <= 16'h8200;
32'hFFFF2954: romout <= 16'h51CA;
32'hFFFF2956: romout <= 16'hFFE8;
32'hFFFF2958: romout <= 16'h4E75;
32'hFFFF295A: romout <= 16'h2079;
32'hFFFF295C: romout <= 16'hFFFF;
32'hFFFF295E: romout <= 16'h241C;
32'hFFFF2960: romout <= 16'h2278;
32'hFFFF2962: romout <= 16'h0624;
32'hFFFF2964: romout <= 16'h103C;
32'hFFFF2966: romout <= 16'h000D;
32'hFFFF2968: romout <= 16'h6100;
32'hFFFF296A: romout <= 16'hFAA6;
32'hFFFF296C: romout <= 16'h103C;
32'hFFFF296E: romout <= 16'h000A;
32'hFFFF2970: romout <= 16'h6100;
32'hFFFF2972: romout <= 16'hFA9E;
32'hFFFF2974: romout <= 16'hB3C8;
32'hFFFF2976: romout <= 16'h6322;
32'hFFFF2978: romout <= 16'h103C;
32'hFFFF297A: romout <= 16'h003A;
32'hFFFF297C: romout <= 16'h6100;
32'hFFFF297E: romout <= 16'hFA92;
32'hFFFF2980: romout <= 16'h1218;
32'hFFFF2982: romout <= 16'h6100;
32'hFFFF2984: romout <= 16'h003A;
32'hFFFF2986: romout <= 16'h1218;
32'hFFFF2988: romout <= 16'h6100;
32'hFFFF298A: romout <= 16'h0034;
32'hFFFF298C: romout <= 16'h1018;
32'hFFFF298E: romout <= 16'hB03C;
32'hFFFF2990: romout <= 16'h000D;
32'hFFFF2992: romout <= 16'h67D0;
32'hFFFF2994: romout <= 16'h6100;
32'hFFFF2996: romout <= 16'hFA7A;
32'hFFFF2998: romout <= 16'h60F2;
32'hFFFF299A: romout <= 16'h103C;
32'hFFFF299C: romout <= 16'h0040;
32'hFFFF299E: romout <= 16'h6100;
32'hFFFF29A0: romout <= 16'hFA70;
32'hFFFF29A2: romout <= 16'h103C;
32'hFFFF29A4: romout <= 16'h000D;
32'hFFFF29A6: romout <= 16'h6100;
32'hFFFF29A8: romout <= 16'hFA68;
32'hFFFF29AA: romout <= 16'h103C;
32'hFFFF29AC: romout <= 16'h000A;
32'hFFFF29AE: romout <= 16'h6100;
32'hFFFF29B0: romout <= 16'hFA60;
32'hFFFF29B2: romout <= 16'h103C;
32'hFFFF29B4: romout <= 16'h001A;
32'hFFFF29B6: romout <= 16'h6100;
32'hFFFF29B8: romout <= 16'hFA58;
32'hFFFF29BA: romout <= 16'h6000;
32'hFFFF29BC: romout <= 16'hFAA4;
32'hFFFF29BE: romout <= 16'h7401;
32'hFFFF29C0: romout <= 16'hE919;
32'hFFFF29C2: romout <= 16'h1001;
32'hFFFF29C4: romout <= 16'h0200;
32'hFFFF29C6: romout <= 16'h000F;
32'hFFFF29C8: romout <= 16'h0600;
32'hFFFF29CA: romout <= 16'h0030;
32'hFFFF29CC: romout <= 16'hB03C;
32'hFFFF29CE: romout <= 16'h0039;
32'hFFFF29D0: romout <= 16'h6302;
32'hFFFF29D2: romout <= 16'h5E00;
32'hFFFF29D4: romout <= 16'h6100;
32'hFFFF29D6: romout <= 16'hFA3A;
32'hFFFF29D8: romout <= 16'h51CA;
32'hFFFF29DA: romout <= 16'hFFE6;
32'hFFFF29DC: romout <= 16'h4E75;
32'hFFFF29DE: romout <= 16'h6100;
32'hFFFF29E0: romout <= 16'h00CA;
32'hFFFF29E2: romout <= 16'h6100;
32'hFFFF29E4: romout <= 16'h05EE;
32'hFFFF29E6: romout <= 16'h2C0F;
32'hFFFF29E8: romout <= 16'h2F00;
32'hFFFF29EA: romout <= 16'h6100;
32'hFFFF29EC: romout <= 16'h00BE;
32'hFFFF29EE: romout <= 16'h225F;
32'hFFFF29F0: romout <= 16'h1280;
32'hFFFF29F2: romout <= 16'h6000;
32'hFFFF29F4: romout <= 16'hFD4E;
32'hFFFF29F6: romout <= 16'h6000;
32'hFFFF29F8: romout <= 16'h03AC;
32'hFFFF29FA: romout <= 16'h6100;
32'hFFFF29FC: romout <= 16'h00AE;
32'hFFFF29FE: romout <= 16'h6100;
32'hFFFF2A00: romout <= 16'h05D2;
32'hFFFF2A02: romout <= 16'h2CF3;
32'hFFFF2A04: romout <= 16'h2F00;
32'hFFFF2A06: romout <= 16'h6100;
32'hFFFF2A08: romout <= 16'h00A2;
32'hFFFF2A0A: romout <= 16'h221F;
32'hFFFF2A0C: romout <= 16'h2400;
32'hFFFF2A0E: romout <= 16'h6100;
32'hFFFF2A10: romout <= 16'hEAEE;
32'hFFFF2A12: romout <= 16'h6000;
32'hFFFF2A14: romout <= 16'hFD2E;
32'hFFFF2A16: romout <= 16'h6100;
32'hFFFF2A18: romout <= 16'h0092;
32'hFFFF2A1A: romout <= 16'h23C0;
32'hFFFF2A1C: romout <= 16'hFFDA;
32'hFFFF2A1E: romout <= 16'hE000;
32'hFFFF2A20: romout <= 16'h6000;
32'hFFFF2A22: romout <= 16'hFD20;
32'hFFFF2A24: romout <= 16'h6100;
32'hFFFF2A26: romout <= 16'h0084;
32'hFFFF2A28: romout <= 16'h23C0;
32'hFFFF2A2A: romout <= 16'hFFDA;
32'hFFFF2A2C: romout <= 16'hE004;
32'hFFFF2A2E: romout <= 16'h6000;
32'hFFFF2A30: romout <= 16'hFD12;
32'hFFFF2A32: romout <= 16'h6100;
32'hFFFF2A34: romout <= 16'h0076;
32'hFFFF2A36: romout <= 16'h6100;
32'hFFFF2A38: romout <= 16'h059A;
32'hFFFF2A3A: romout <= 16'h2C49;
32'hFFFF2A3C: romout <= 16'h2F00;
32'hFFFF2A3E: romout <= 16'h6100;
32'hFFFF2A40: romout <= 16'h006A;
32'hFFFF2A42: romout <= 16'h6100;
32'hFFFF2A44: romout <= 16'h058E;
32'hFFFF2A46: romout <= 16'h2C41;
32'hFFFF2A48: romout <= 16'h2F00;
32'hFFFF2A4A: romout <= 16'h6100;
32'hFFFF2A4C: romout <= 16'h005E;
32'hFFFF2A4E: romout <= 16'h6100;
32'hFFFF2A50: romout <= 16'h0582;
32'hFFFF2A52: romout <= 16'h2C3B;
32'hFFFF2A54: romout <= 16'h2F00;
32'hFFFF2A56: romout <= 16'h6100;
32'hFFFF2A58: romout <= 16'h0052;
32'hFFFF2A5A: romout <= 16'h33C0;
32'hFFFF2A5C: romout <= 16'hFFDA;
32'hFFFF2A5E: romout <= 16'hE00E;
32'hFFFF2A60: romout <= 16'h201F;
32'hFFFF2A62: romout <= 16'h33C0;
32'hFFFF2A64: romout <= 16'hFFDA;
32'hFFFF2A66: romout <= 16'hE00C;
32'hFFFF2A68: romout <= 16'h201F;
32'hFFFF2A6A: romout <= 16'h33C0;
32'hFFFF2A6C: romout <= 16'hFFDA;
32'hFFFF2A6E: romout <= 16'hE00A;
32'hFFFF2A70: romout <= 16'h201F;
32'hFFFF2A72: romout <= 16'h33C0;
32'hFFFF2A74: romout <= 16'hFFDA;
32'hFFFF2A76: romout <= 16'hE008;
32'hFFFF2A78: romout <= 16'h33FC;
32'hFFFF2A7A: romout <= 16'h0002;
32'hFFFF2A7C: romout <= 16'hFFDA;
32'hFFFF2A7E: romout <= 16'hE01E;
32'hFFFF2A80: romout <= 16'h6000;
32'hFFFF2A82: romout <= 16'hFCC0;
32'hFFFF2A84: romout <= 16'h6000;
32'hFFFF2A86: romout <= 16'h031E;
32'hFFFF2A88: romout <= 16'h588F;
32'hFFFF2A8A: romout <= 16'h6000;
32'hFFFF2A8C: romout <= 16'h0318;
32'hFFFF2A8E: romout <= 16'h508F;
32'hFFFF2A90: romout <= 16'h6000;
32'hFFFF2A92: romout <= 16'h0312;
32'hFFFF2A94: romout <= 16'h6100;
32'hFFFF2A96: romout <= 16'h0014;
32'hFFFF2A98: romout <= 16'h4A80;
32'hFFFF2A9A: romout <= 16'h6700;
32'hFFFF2A9C: romout <= 16'h0354;
32'hFFFF2A9E: romout <= 16'h2F08;
32'hFFFF2AA0: romout <= 16'h2240;
32'hFFFF2AA2: romout <= 16'h4E91;
32'hFFFF2AA4: romout <= 16'h205F;
32'hFFFF2AA6: romout <= 16'h6000;
32'hFFFF2AA8: romout <= 16'hFC9A;
32'hFFFF2AAA: romout <= 16'h6100;
32'hFFFF2AAC: romout <= 16'h0066;
32'hFFFF2AAE: romout <= 16'h2F00;
32'hFFFF2AB0: romout <= 16'h43F9;
32'hFFFF2AB2: romout <= 16'hFFFF;
32'hFFFF2AB4: romout <= 16'h258B;
32'hFFFF2AB6: romout <= 16'h45F9;
32'hFFFF2AB8: romout <= 16'hFFFF;
32'hFFFF2ABA: romout <= 16'h25E0;
32'hFFFF2ABC: romout <= 16'h6000;
32'hFFFF2ABE: romout <= 16'hFB3C;
32'hFFFF2AC0: romout <= 16'h6100;
32'hFFFF2AC2: romout <= 16'h003E;
32'hFFFF2AC4: romout <= 16'h6D2E;
32'hFFFF2AC6: romout <= 16'h6030;
32'hFFFF2AC8: romout <= 16'h6100;
32'hFFFF2ACA: romout <= 16'h0036;
32'hFFFF2ACC: romout <= 16'h6726;
32'hFFFF2ACE: romout <= 16'h6028;
32'hFFFF2AD0: romout <= 16'h6100;
32'hFFFF2AD2: romout <= 16'h002E;
32'hFFFF2AD4: romout <= 16'h6F1E;
32'hFFFF2AD6: romout <= 16'h6020;
32'hFFFF2AD8: romout <= 16'h6100;
32'hFFFF2ADA: romout <= 16'h0026;
32'hFFFF2ADC: romout <= 16'h6E16;
32'hFFFF2ADE: romout <= 16'h6018;
32'hFFFF2AE0: romout <= 16'h6100;
32'hFFFF2AE2: romout <= 16'h001E;
32'hFFFF2AE4: romout <= 16'h660E;
32'hFFFF2AE6: romout <= 16'h6010;
32'hFFFF2AE8: romout <= 16'h4E75;
32'hFFFF2AEA: romout <= 16'h6100;
32'hFFFF2AEC: romout <= 16'h0014;
32'hFFFF2AEE: romout <= 16'h6C04;
32'hFFFF2AF0: romout <= 16'h6006;
32'hFFFF2AF2: romout <= 16'h4E75;
32'hFFFF2AF4: romout <= 16'h4280;
32'hFFFF2AF6: romout <= 16'h4E75;
32'hFFFF2AF8: romout <= 16'h7001;
32'hFFFF2AFA: romout <= 16'h4E75;
32'hFFFF2AFC: romout <= 16'h201F;
32'hFFFF2AFE: romout <= 16'h4E75;
32'hFFFF2B00: romout <= 16'h201F;
32'hFFFF2B02: romout <= 16'h221F;
32'hFFFF2B04: romout <= 16'h2F00;
32'hFFFF2B06: romout <= 16'h2F01;
32'hFFFF2B08: romout <= 16'h6100;
32'hFFFF2B0A: romout <= 16'h0008;
32'hFFFF2B0C: romout <= 16'h221F;
32'hFFFF2B0E: romout <= 16'hB280;
32'hFFFF2B10: romout <= 16'h4E75;
32'hFFFF2B12: romout <= 16'h6100;
32'hFFFF2B14: romout <= 16'h04BE;
32'hFFFF2B16: romout <= 16'h2D05;
32'hFFFF2B18: romout <= 16'h4280;
32'hFFFF2B1A: romout <= 16'h603C;
32'hFFFF2B1C: romout <= 16'h6100;
32'hFFFF2B1E: romout <= 16'h04B4;
32'hFFFF2B20: romout <= 16'h2111;
32'hFFFF2B22: romout <= 16'h4280;
32'hFFFF2B24: romout <= 16'h2F00;
32'hFFFF2B26: romout <= 16'h6100;
32'hFFFF2B28: romout <= 16'h0062;
32'hFFFF2B2A: romout <= 16'h4680;
32'hFFFF2B2C: romout <= 16'h4EF9;
32'hFFFF2B2E: romout <= 16'hFFFF;
32'hFFFF2B30: romout <= 16'h2B48;
32'hFFFF2B32: romout <= 16'h6100;
32'hFFFF2B34: romout <= 16'h049E;
32'hFFFF2B36: romout <= 16'h2B01;
32'hFFFF2B38: romout <= 16'h6100;
32'hFFFF2B3A: romout <= 16'h0050;
32'hFFFF2B3C: romout <= 16'h6100;
32'hFFFF2B3E: romout <= 16'h0494;
32'hFFFF2B40: romout <= 16'h2B11;
32'hFFFF2B42: romout <= 16'h2F00;
32'hFFFF2B44: romout <= 16'h6100;
32'hFFFF2B46: romout <= 16'h0044;
32'hFFFF2B48: romout <= 16'h221F;
32'hFFFF2B4A: romout <= 16'hD081;
32'hFFFF2B4C: romout <= 16'h6900;
32'hFFFF2B4E: romout <= 16'h02A2;
32'hFFFF2B50: romout <= 16'h60EA;
32'hFFFF2B52: romout <= 16'h6100;
32'hFFFF2B54: romout <= 16'h047E;
32'hFFFF2B56: romout <= 16'h2D0F;
32'hFFFF2B58: romout <= 16'h2F00;
32'hFFFF2B5A: romout <= 16'h6100;
32'hFFFF2B5C: romout <= 16'h002E;
32'hFFFF2B5E: romout <= 16'h4480;
32'hFFFF2B60: romout <= 16'h4EF9;
32'hFFFF2B62: romout <= 16'hFFFF;
32'hFFFF2B64: romout <= 16'h2B48;
32'hFFFF2B66: romout <= 16'h6100;
32'hFFFF2B68: romout <= 16'h046A;
32'hFFFF2B6A: romout <= 16'h260D;
32'hFFFF2B6C: romout <= 16'h2F00;
32'hFFFF2B6E: romout <= 16'h6100;
32'hFFFF2B70: romout <= 16'h001A;
32'hFFFF2B72: romout <= 16'h221F;
32'hFFFF2B74: romout <= 16'hC081;
32'hFFFF2B76: romout <= 16'h60C4;
32'hFFFF2B78: romout <= 16'h6100;
32'hFFFF2B7A: romout <= 16'h0458;
32'hFFFF2B7C: romout <= 16'h7C73;
32'hFFFF2B7E: romout <= 16'h2F00;
32'hFFFF2B80: romout <= 16'h6100;
32'hFFFF2B82: romout <= 16'h0008;
32'hFFFF2B84: romout <= 16'h221F;
32'hFFFF2B86: romout <= 16'h8081;
32'hFFFF2B88: romout <= 16'h60B2;
32'hFFFF2B8A: romout <= 16'h6100;
32'hFFFF2B8C: romout <= 16'h002C;
32'hFFFF2B8E: romout <= 16'h6100;
32'hFFFF2B90: romout <= 16'h0442;
32'hFFFF2B92: romout <= 16'h2A0F;
32'hFFFF2B94: romout <= 16'h2F00;
32'hFFFF2B96: romout <= 16'h6100;
32'hFFFF2B98: romout <= 16'h0020;
32'hFFFF2B9A: romout <= 16'h221F;
32'hFFFF2B9C: romout <= 16'h6100;
32'hFFFF2B9E: romout <= 16'h00D2;
32'hFFFF2BA0: romout <= 16'h60EC;
32'hFFFF2BA2: romout <= 16'h6100;
32'hFFFF2BA4: romout <= 16'h042E;
32'hFFFF2BA6: romout <= 16'h2F49;
32'hFFFF2BA8: romout <= 16'h2F00;
32'hFFFF2BAA: romout <= 16'h6100;
32'hFFFF2BAC: romout <= 16'h000C;
32'hFFFF2BAE: romout <= 16'h221F;
32'hFFFF2BB0: romout <= 16'hC141;
32'hFFFF2BB2: romout <= 16'h6100;
32'hFFFF2BB4: romout <= 16'h00FE;
32'hFFFF2BB6: romout <= 16'h60D6;
32'hFFFF2BB8: romout <= 16'h43F9;
32'hFFFF2BBA: romout <= 16'hFFFF;
32'hFFFF2BBC: romout <= 16'h2569;
32'hFFFF2BBE: romout <= 16'h45F9;
32'hFFFF2BC0: romout <= 16'hFFFF;
32'hFFFF2BC2: romout <= 16'h25C8;
32'hFFFF2BC4: romout <= 16'h6000;
32'hFFFF2BC6: romout <= 16'hFA34;
32'hFFFF2BC8: romout <= 16'h6100;
32'hFFFF2BCA: romout <= 16'h002C;
32'hFFFF2BCC: romout <= 16'h6508;
32'hFFFF2BCE: romout <= 16'h2240;
32'hFFFF2BD0: romout <= 16'h4280;
32'hFFFF2BD2: romout <= 16'h2011;
32'hFFFF2BD4: romout <= 16'h4E75;
32'hFFFF2BD6: romout <= 16'h6100;
32'hFFFF2BD8: romout <= 16'h0414;
32'hFFFF2BDA: romout <= 16'h2001;
32'hFFFF2BDC: romout <= 16'h4A82;
32'hFFFF2BDE: romout <= 16'h66F4;
32'hFFFF2BE0: romout <= 16'h6100;
32'hFFFF2BE2: romout <= 16'h03F0;
32'hFFFF2BE4: romout <= 16'h280D;
32'hFFFF2BE6: romout <= 16'h6100;
32'hFFFF2BE8: romout <= 16'hFEC2;
32'hFFFF2BEA: romout <= 16'h6100;
32'hFFFF2BEC: romout <= 16'h03E6;
32'hFFFF2BEE: romout <= 16'h2903;
32'hFFFF2BF0: romout <= 16'h4E75;
32'hFFFF2BF2: romout <= 16'h6000;
32'hFFFF2BF4: romout <= 16'h01B0;
32'hFFFF2BF6: romout <= 16'h6100;
32'hFFFF2BF8: romout <= 16'h042C;
32'hFFFF2BFA: romout <= 16'h4280;
32'hFFFF2BFC: romout <= 16'h1010;
32'hFFFF2BFE: romout <= 16'h0400;
32'hFFFF2C00: romout <= 16'h0040;
32'hFFFF2C02: romout <= 16'h6554;
32'hFFFF2C04: romout <= 16'h6628;
32'hFFFF2C06: romout <= 16'h5288;
32'hFFFF2C08: romout <= 16'h6100;
32'hFFFF2C0A: romout <= 16'hFFD6;
32'hFFFF2C0C: romout <= 16'hD080;
32'hFFFF2C0E: romout <= 16'h6500;
32'hFFFF2C10: romout <= 16'h01E0;
32'hFFFF2C12: romout <= 16'hD080;
32'hFFFF2C14: romout <= 16'h6500;
32'hFFFF2C16: romout <= 16'h01DA;
32'hFFFF2C18: romout <= 16'h2F00;
32'hFFFF2C1A: romout <= 16'h6100;
32'hFFFF2C1C: romout <= 16'h012C;
32'hFFFF2C1E: romout <= 16'h221F;
32'hFFFF2C20: romout <= 16'hB081;
32'hFFFF2C22: romout <= 16'h6300;
32'hFFFF2C24: romout <= 16'h01C2;
32'hFFFF2C26: romout <= 16'h2038;
32'hFFFF2C28: romout <= 16'h0628;
32'hFFFF2C2A: romout <= 16'h9081;
32'hFFFF2C2C: romout <= 16'h4E75;
32'hFFFF2C2E: romout <= 16'hB03C;
32'hFFFF2C30: romout <= 16'h001B;
32'hFFFF2C32: romout <= 16'h0A3C;
32'hFFFF2C34: romout <= 16'h0001;
32'hFFFF2C36: romout <= 16'h6520;
32'hFFFF2C38: romout <= 16'h5288;
32'hFFFF2C3A: romout <= 16'h4281;
32'hFFFF2C3C: romout <= 16'h1210;
32'hFFFF2C3E: romout <= 16'h6100;
32'hFFFF2C40: romout <= 16'h001A;
32'hFFFF2C42: romout <= 16'h0C01;
32'hFFFF2C44: romout <= 16'h00FF;
32'hFFFF2C46: romout <= 16'h6706;
32'hFFFF2C48: romout <= 16'h5288;
32'hFFFF2C4A: romout <= 16'hEB81;
32'hFFFF2C4C: romout <= 16'hD081;
32'hFFFF2C4E: romout <= 16'hD080;
32'hFFFF2C50: romout <= 16'hD080;
32'hFFFF2C52: romout <= 16'h2238;
32'hFFFF2C54: romout <= 16'h0628;
32'hFFFF2C56: romout <= 16'hD081;
32'hFFFF2C58: romout <= 16'h4E75;
32'hFFFF2C5A: romout <= 16'h0C01;
32'hFFFF2C5C: romout <= 16'h0041;
32'hFFFF2C5E: romout <= 16'h650C;
32'hFFFF2C60: romout <= 16'h0C01;
32'hFFFF2C62: romout <= 16'h005A;
32'hFFFF2C64: romout <= 16'h6206;
32'hFFFF2C66: romout <= 16'h0401;
32'hFFFF2C68: romout <= 16'h0041;
32'hFFFF2C6A: romout <= 16'h4E75;
32'hFFFF2C6C: romout <= 16'h72FF;
32'hFFFF2C6E: romout <= 16'h4E75;
32'hFFFF2C70: romout <= 16'h2801;
32'hFFFF2C72: romout <= 16'hB184;
32'hFFFF2C74: romout <= 16'h4A80;
32'hFFFF2C76: romout <= 16'h6A02;
32'hFFFF2C78: romout <= 16'h4480;
32'hFFFF2C7A: romout <= 16'h4A81;
32'hFFFF2C7C: romout <= 16'h6A02;
32'hFFFF2C7E: romout <= 16'h4481;
32'hFFFF2C80: romout <= 16'hB2BC;
32'hFFFF2C82: romout <= 16'h0000;
32'hFFFF2C84: romout <= 16'hFFFF;
32'hFFFF2C86: romout <= 16'h630C;
32'hFFFF2C88: romout <= 16'hC141;
32'hFFFF2C8A: romout <= 16'hB2BC;
32'hFFFF2C8C: romout <= 16'h0000;
32'hFFFF2C8E: romout <= 16'hFFFF;
32'hFFFF2C90: romout <= 16'h6200;
32'hFFFF2C92: romout <= 16'h015E;
32'hFFFF2C94: romout <= 16'h2400;
32'hFFFF2C96: romout <= 16'hC4C1;
32'hFFFF2C98: romout <= 16'h4840;
32'hFFFF2C9A: romout <= 16'hC0C1;
32'hFFFF2C9C: romout <= 16'h4840;
32'hFFFF2C9E: romout <= 16'h4A80;
32'hFFFF2CA0: romout <= 16'h6600;
32'hFFFF2CA2: romout <= 16'h014E;
32'hFFFF2CA4: romout <= 16'hD082;
32'hFFFF2CA6: romout <= 16'h6B00;
32'hFFFF2CA8: romout <= 16'h0148;
32'hFFFF2CAA: romout <= 16'h4A84;
32'hFFFF2CAC: romout <= 16'h6A02;
32'hFFFF2CAE: romout <= 16'h4480;
32'hFFFF2CB0: romout <= 16'h4E75;
32'hFFFF2CB2: romout <= 16'h4A81;
32'hFFFF2CB4: romout <= 16'h6700;
32'hFFFF2CB6: romout <= 16'h013A;
32'hFFFF2CB8: romout <= 16'h2401;
32'hFFFF2CBA: romout <= 16'h2801;
32'hFFFF2CBC: romout <= 16'hB184;
32'hFFFF2CBE: romout <= 16'h4A80;
32'hFFFF2CC0: romout <= 16'h6A02;
32'hFFFF2CC2: romout <= 16'h4480;
32'hFFFF2CC4: romout <= 16'h4A81;
32'hFFFF2CC6: romout <= 16'h6A02;
32'hFFFF2CC8: romout <= 16'h4481;
32'hFFFF2CCA: romout <= 16'h761F;
32'hFFFF2CCC: romout <= 16'h2200;
32'hFFFF2CCE: romout <= 16'h4280;
32'hFFFF2CD0: romout <= 16'hD281;
32'hFFFF2CD2: romout <= 16'hD180;
32'hFFFF2CD4: romout <= 16'h6708;
32'hFFFF2CD6: romout <= 16'hB082;
32'hFFFF2CD8: romout <= 16'h6B04;
32'hFFFF2CDA: romout <= 16'h5281;
32'hFFFF2CDC: romout <= 16'h9082;
32'hFFFF2CDE: romout <= 16'h51CB;
32'hFFFF2CE0: romout <= 16'hFFF0;
32'hFFFF2CE2: romout <= 16'hC141;
32'hFFFF2CE4: romout <= 16'h4A84;
32'hFFFF2CE6: romout <= 16'h6A04;
32'hFFFF2CE8: romout <= 16'h4480;
32'hFFFF2CEA: romout <= 16'h4481;
32'hFFFF2CEC: romout <= 16'h4E75;
32'hFFFF2CEE: romout <= 16'h6100;
32'hFFFF2CF0: romout <= 16'hFEF0;
32'hFFFF2CF2: romout <= 16'h2240;
32'hFFFF2CF4: romout <= 16'h4280;
32'hFFFF2CF6: romout <= 16'h1011;
32'hFFFF2CF8: romout <= 16'h4E75;
32'hFFFF2CFA: romout <= 16'h6100;
32'hFFFF2CFC: romout <= 16'hFEE4;
32'hFFFF2CFE: romout <= 16'h4A80;
32'hFFFF2D00: romout <= 16'h6700;
32'hFFFF2D02: romout <= 16'h00EE;
32'hFFFF2D04: romout <= 16'h6B00;
32'hFFFF2D06: romout <= 16'h00EA;
32'hFFFF2D08: romout <= 16'h2200;
32'hFFFF2D0A: romout <= 16'h3039;
32'hFFFF2D0C: romout <= 16'hFFDC;
32'hFFFF2D0E: romout <= 16'h0C02;
32'hFFFF2D10: romout <= 16'h4840;
32'hFFFF2D12: romout <= 16'h3039;
32'hFFFF2D14: romout <= 16'hFFDC;
32'hFFFF2D16: romout <= 16'h0C00;
32'hFFFF2D18: romout <= 16'h0880;
32'hFFFF2D1A: romout <= 16'h001F;
32'hFFFF2D1C: romout <= 16'h6100;
32'hFFFF2D1E: romout <= 16'hFF94;
32'hFFFF2D20: romout <= 16'h2001;
32'hFFFF2D22: romout <= 16'h5280;
32'hFFFF2D24: romout <= 16'h4E75;
32'hFFFF2D26: romout <= 16'h6100;
32'hFFFF2D28: romout <= 16'hFEB8;
32'hFFFF2D2A: romout <= 16'h4A80;
32'hFFFF2D2C: romout <= 16'h6A06;
32'hFFFF2D2E: romout <= 16'h4480;
32'hFFFF2D30: romout <= 16'h6B00;
32'hFFFF2D32: romout <= 16'h00BE;
32'hFFFF2D34: romout <= 16'h4E75;
32'hFFFF2D36: romout <= 16'h6100;
32'hFFFF2D38: romout <= 16'hFEA8;
32'hFFFF2D3A: romout <= 16'h4A80;
32'hFFFF2D3C: romout <= 16'h6704;
32'hFFFF2D3E: romout <= 16'h6B04;
32'hFFFF2D40: romout <= 16'h7001;
32'hFFFF2D42: romout <= 16'h4E75;
32'hFFFF2D44: romout <= 16'h70FF;
32'hFFFF2D46: romout <= 16'h4E75;
32'hFFFF2D48: romout <= 16'h2038;
32'hFFFF2D4A: romout <= 16'h0628;
32'hFFFF2D4C: romout <= 16'h90B8;
32'hFFFF2D4E: romout <= 16'h0624;
32'hFFFF2D50: romout <= 16'h4E75;
32'hFFFF2D52: romout <= 16'h2038;
32'hFFFF2D54: romout <= 16'h0400;
32'hFFFF2D56: romout <= 16'h4E75;
32'hFFFF2D58: romout <= 16'h6100;
32'hFFFF2D5A: romout <= 16'hF154;
32'hFFFF2D5C: romout <= 16'h0280;
32'hFFFF2D5E: romout <= 16'h0000;
32'hFFFF2D60: romout <= 16'hFFFF;
32'hFFFF2D62: romout <= 16'h4E75;
32'hFFFF2D64: romout <= 16'h6100;
32'hFFFF2D66: romout <= 16'hFE90;
32'hFFFF2D68: romout <= 16'h653A;
32'hFFFF2D6A: romout <= 16'h2F00;
32'hFFFF2D6C: romout <= 16'h6100;
32'hFFFF2D6E: romout <= 16'h0264;
32'hFFFF2D70: romout <= 16'h3D0B;
32'hFFFF2D72: romout <= 16'h6100;
32'hFFFF2D74: romout <= 16'hFD36;
32'hFFFF2D76: romout <= 16'h2C5F;
32'hFFFF2D78: romout <= 16'h2C80;
32'hFFFF2D7A: romout <= 16'h4E75;
32'hFFFF2D7C: romout <= 16'h6026;
32'hFFFF2D7E: romout <= 16'h6100;
32'hFFFF2D80: romout <= 16'h0252;
32'hFFFF2D82: romout <= 16'h3A07;
32'hFFFF2D84: romout <= 16'h588F;
32'hFFFF2D86: romout <= 16'h6000;
32'hFFFF2D88: romout <= 16'hF904;
32'hFFFF2D8A: romout <= 16'h6100;
32'hFFFF2D8C: romout <= 16'h0246;
32'hFFFF2D8E: romout <= 16'h0D07;
32'hFFFF2D90: romout <= 16'h588F;
32'hFFFF2D92: romout <= 16'h6000;
32'hFFFF2D94: romout <= 16'hF8DC;
32'hFFFF2D96: romout <= 16'h4E75;
32'hFFFF2D98: romout <= 16'h6100;
32'hFFFF2D9A: romout <= 16'h028A;
32'hFFFF2D9C: romout <= 16'h0C10;
32'hFFFF2D9E: romout <= 16'h000D;
32'hFFFF2DA0: romout <= 16'h6602;
32'hFFFF2DA2: romout <= 16'h4E75;
32'hFFFF2DA4: romout <= 16'h2F08;
32'hFFFF2DA6: romout <= 16'h4DF9;
32'hFFFF2DA8: romout <= 16'hFFFF;
32'hFFFF2DAA: romout <= 16'h312C;
32'hFFFF2DAC: romout <= 16'h6100;
32'hFFFF2DAE: romout <= 16'h02E6;
32'hFFFF2DB0: romout <= 16'h205F;
32'hFFFF2DB2: romout <= 16'h2038;
32'hFFFF2DB4: romout <= 16'h0604;
32'hFFFF2DB6: romout <= 16'h6700;
32'hFFFF2DB8: romout <= 16'hF6A8;
32'hFFFF2DBA: romout <= 16'hB0BC;
32'hFFFF2DBC: romout <= 16'hFFFF;
32'hFFFF2DBE: romout <= 16'hFFFF;
32'hFFFF2DC0: romout <= 16'h6700;
32'hFFFF2DC2: romout <= 16'hFAAA;
32'hFFFF2DC4: romout <= 16'h1F10;
32'hFFFF2DC6: romout <= 16'h4210;
32'hFFFF2DC8: romout <= 16'h2278;
32'hFFFF2DCA: romout <= 16'h0604;
32'hFFFF2DCC: romout <= 16'h6100;
32'hFFFF2DCE: romout <= 16'h01E8;
32'hFFFF2DD0: romout <= 16'h109F;
32'hFFFF2DD2: romout <= 16'h103C;
32'hFFFF2DD4: romout <= 16'h003F;
32'hFFFF2DD6: romout <= 16'h6100;
32'hFFFF2DD8: romout <= 16'hF630;
32'hFFFF2DDA: romout <= 16'h4280;
32'hFFFF2DDC: romout <= 16'h5389;
32'hFFFF2DDE: romout <= 16'h6100;
32'hFFFF2DE0: romout <= 16'h013E;
32'hFFFF2DE2: romout <= 16'h6000;
32'hFFFF2DE4: romout <= 16'hF67C;
32'hFFFF2DE6: romout <= 16'h2F08;
32'hFFFF2DE8: romout <= 16'h4DF9;
32'hFFFF2DEA: romout <= 16'hFFFF;
32'hFFFF2DEC: romout <= 16'h3134;
32'hFFFF2DEE: romout <= 16'h60BC;
32'hFFFF2DF0: romout <= 16'h2F08;
32'hFFFF2DF2: romout <= 16'h4DF9;
32'hFFFF2DF4: romout <= 16'hFFFF;
32'hFFFF2DF6: romout <= 16'h3125;
32'hFFFF2DF8: romout <= 16'h60B2;
32'hFFFF2DFA: romout <= 16'h6100;
32'hFFFF2DFC: romout <= 16'hF60C;
32'hFFFF2DFE: romout <= 16'h103C;
32'hFFFF2E00: romout <= 16'h0020;
32'hFFFF2E02: romout <= 16'h6100;
32'hFFFF2E04: romout <= 16'hF604;
32'hFFFF2E06: romout <= 16'h41F8;
32'hFFFF2E08: romout <= 16'h0630;
32'hFFFF2E0A: romout <= 16'h6100;
32'hFFFF2E0C: romout <= 16'h0270;
32'hFFFF2E0E: romout <= 16'h67FA;
32'hFFFF2E10: romout <= 16'hB03C;
32'hFFFF2E12: romout <= 16'h0008;
32'hFFFF2E14: romout <= 16'h6726;
32'hFFFF2E16: romout <= 16'hB03C;
32'hFFFF2E18: romout <= 16'h0018;
32'hFFFF2E1A: romout <= 16'h6744;
32'hFFFF2E1C: romout <= 16'hB03C;
32'hFFFF2E1E: romout <= 16'h000D;
32'hFFFF2E20: romout <= 16'h6706;
32'hFFFF2E22: romout <= 16'hB03C;
32'hFFFF2E24: romout <= 16'h0020;
32'hFFFF2E26: romout <= 16'h65E2;
32'hFFFF2E28: romout <= 16'h10C0;
32'hFFFF2E2A: romout <= 16'h6100;
32'hFFFF2E2C: romout <= 16'hF5DC;
32'hFFFF2E2E: romout <= 16'hB03C;
32'hFFFF2E30: romout <= 16'h000D;
32'hFFFF2E32: romout <= 16'h675C;
32'hFFFF2E34: romout <= 16'hB1FC;
32'hFFFF2E36: romout <= 16'h0000;
32'hFFFF2E38: romout <= 16'h067F;
32'hFFFF2E3A: romout <= 16'h65CE;
32'hFFFF2E3C: romout <= 16'h103C;
32'hFFFF2E3E: romout <= 16'h0008;
32'hFFFF2E40: romout <= 16'h6100;
32'hFFFF2E42: romout <= 16'hF5C6;
32'hFFFF2E44: romout <= 16'h103C;
32'hFFFF2E46: romout <= 16'h0020;
32'hFFFF2E48: romout <= 16'h6100;
32'hFFFF2E4A: romout <= 16'hF5BE;
32'hFFFF2E4C: romout <= 16'hB1FC;
32'hFFFF2E4E: romout <= 16'h0000;
32'hFFFF2E50: romout <= 16'h0630;
32'hFFFF2E52: romout <= 16'h63B6;
32'hFFFF2E54: romout <= 16'h103C;
32'hFFFF2E56: romout <= 16'h0008;
32'hFFFF2E58: romout <= 16'h6100;
32'hFFFF2E5A: romout <= 16'hF5AE;
32'hFFFF2E5C: romout <= 16'h5388;
32'hFFFF2E5E: romout <= 16'h60AA;
32'hFFFF2E60: romout <= 16'h2208;
32'hFFFF2E62: romout <= 16'h0481;
32'hFFFF2E64: romout <= 16'h0000;
32'hFFFF2E66: romout <= 16'h0630;
32'hFFFF2E68: romout <= 16'h671E;
32'hFFFF2E6A: romout <= 16'h5381;
32'hFFFF2E6C: romout <= 16'h103C;
32'hFFFF2E6E: romout <= 16'h0008;
32'hFFFF2E70: romout <= 16'h6100;
32'hFFFF2E72: romout <= 16'hF596;
32'hFFFF2E74: romout <= 16'h103C;
32'hFFFF2E76: romout <= 16'h0020;
32'hFFFF2E78: romout <= 16'h6100;
32'hFFFF2E7A: romout <= 16'hF58E;
32'hFFFF2E7C: romout <= 16'h103C;
32'hFFFF2E7E: romout <= 16'h0008;
32'hFFFF2E80: romout <= 16'h6100;
32'hFFFF2E82: romout <= 16'hF586;
32'hFFFF2E84: romout <= 16'h51C9;
32'hFFFF2E86: romout <= 16'hFFE6;
32'hFFFF2E88: romout <= 16'h41F8;
32'hFFFF2E8A: romout <= 16'h0630;
32'hFFFF2E8C: romout <= 16'h6000;
32'hFFFF2E8E: romout <= 16'hFF7C;
32'hFFFF2E90: romout <= 16'h103C;
32'hFFFF2E92: romout <= 16'h000A;
32'hFFFF2E94: romout <= 16'h6100;
32'hFFFF2E96: romout <= 16'hF572;
32'hFFFF2E98: romout <= 16'h4E75;
32'hFFFF2E9A: romout <= 16'hB2BC;
32'hFFFF2E9C: romout <= 16'h0000;
32'hFFFF2E9E: romout <= 16'hFFFF;
32'hFFFF2EA0: romout <= 16'h6400;
32'hFFFF2EA2: romout <= 16'hFF4E;
32'hFFFF2EA4: romout <= 16'h2279;
32'hFFFF2EA6: romout <= 16'hFFFF;
32'hFFFF2EA8: romout <= 16'h241C;
32'hFFFF2EAA: romout <= 16'h2478;
32'hFFFF2EAC: romout <= 16'h0624;
32'hFFFF2EAE: romout <= 16'h538A;
32'hFFFF2EB0: romout <= 16'hB5C9;
32'hFFFF2EB2: romout <= 16'h650C;
32'hFFFF2EB4: romout <= 16'h1411;
32'hFFFF2EB6: romout <= 16'hE14A;
32'hFFFF2EB8: romout <= 16'h1429;
32'hFFFF2EBA: romout <= 16'h0001;
32'hFFFF2EBC: romout <= 16'hB441;
32'hFFFF2EBE: romout <= 16'h6502;
32'hFFFF2EC0: romout <= 16'h4E75;
32'hFFFF2EC2: romout <= 16'h5489;
32'hFFFF2EC4: romout <= 16'h0C19;
32'hFFFF2EC6: romout <= 16'h000D;
32'hFFFF2EC8: romout <= 16'h66FA;
32'hFFFF2ECA: romout <= 16'h60DE;
32'hFFFF2ECC: romout <= 16'hB7C9;
32'hFFFF2ECE: romout <= 16'h6704;
32'hFFFF2ED0: romout <= 16'h14D9;
32'hFFFF2ED2: romout <= 16'h60F8;
32'hFFFF2ED4: romout <= 16'h4E75;
32'hFFFF2ED6: romout <= 16'hB5C9;
32'hFFFF2ED8: romout <= 16'h67FA;
32'hFFFF2EDA: romout <= 16'h1721;
32'hFFFF2EDC: romout <= 16'h60F8;
32'hFFFF2EDE: romout <= 16'h2C5F;
32'hFFFF2EE0: romout <= 16'h21DF;
32'hFFFF2EE2: romout <= 16'h0610;
32'hFFFF2EE4: romout <= 16'h6710;
32'hFFFF2EE6: romout <= 16'h21DF;
32'hFFFF2EE8: romout <= 16'h0614;
32'hFFFF2EEA: romout <= 16'h21DF;
32'hFFFF2EEC: romout <= 16'h0618;
32'hFFFF2EEE: romout <= 16'h21DF;
32'hFFFF2EF0: romout <= 16'h061C;
32'hFFFF2EF2: romout <= 16'h21DF;
32'hFFFF2EF4: romout <= 16'h0620;
32'hFFFF2EF6: romout <= 16'h4ED6;
32'hFFFF2EF8: romout <= 16'h2238;
32'hFFFF2EFA: romout <= 16'h062C;
32'hFFFF2EFC: romout <= 16'h928F;
32'hFFFF2EFE: romout <= 16'h6400;
32'hFFFF2F00: romout <= 16'hFEE6;
32'hFFFF2F02: romout <= 16'h2C5F;
32'hFFFF2F04: romout <= 16'h2238;
32'hFFFF2F06: romout <= 16'h0610;
32'hFFFF2F08: romout <= 16'h6710;
32'hFFFF2F0A: romout <= 16'h2F38;
32'hFFFF2F0C: romout <= 16'h0620;
32'hFFFF2F0E: romout <= 16'h2F38;
32'hFFFF2F10: romout <= 16'h061C;
32'hFFFF2F12: romout <= 16'h2F38;
32'hFFFF2F14: romout <= 16'h0618;
32'hFFFF2F16: romout <= 16'h2F38;
32'hFFFF2F18: romout <= 16'h0614;
32'hFFFF2F1A: romout <= 16'h2F01;
32'hFFFF2F1C: romout <= 16'h4ED6;
32'hFFFF2F1E: romout <= 16'h1200;
32'hFFFF2F20: romout <= 16'h1019;
32'hFFFF2F22: romout <= 16'hB200;
32'hFFFF2F24: romout <= 16'h6712;
32'hFFFF2F26: romout <= 16'h6100;
32'hFFFF2F28: romout <= 16'hF4E0;
32'hFFFF2F2A: romout <= 16'hB03C;
32'hFFFF2F2C: romout <= 16'h000D;
32'hFFFF2F2E: romout <= 16'h66F0;
32'hFFFF2F30: romout <= 16'h103C;
32'hFFFF2F32: romout <= 16'h000A;
32'hFFFF2F34: romout <= 16'h6100;
32'hFFFF2F36: romout <= 16'hF4D2;
32'hFFFF2F38: romout <= 16'h4E75;
32'hFFFF2F3A: romout <= 16'h6100;
32'hFFFF2F3C: romout <= 16'h0096;
32'hFFFF2F3E: romout <= 16'h221B;
32'hFFFF2F40: romout <= 16'h103C;
32'hFFFF2F42: romout <= 16'h0022;
32'hFFFF2F44: romout <= 16'h2248;
32'hFFFF2F46: romout <= 16'h6100;
32'hFFFF2F48: romout <= 16'hFFD6;
32'hFFFF2F4A: romout <= 16'h2049;
32'hFFFF2F4C: romout <= 16'h225F;
32'hFFFF2F4E: romout <= 16'hB03C;
32'hFFFF2F50: romout <= 16'h000A;
32'hFFFF2F52: romout <= 16'h6700;
32'hFFFF2F54: romout <= 16'hF71C;
32'hFFFF2F56: romout <= 16'h5489;
32'hFFFF2F58: romout <= 16'h4ED1;
32'hFFFF2F5A: romout <= 16'h6100;
32'hFFFF2F5C: romout <= 16'h0076;
32'hFFFF2F5E: romout <= 16'h2707;
32'hFFFF2F60: romout <= 16'h103C;
32'hFFFF2F62: romout <= 16'h0027;
32'hFFFF2F64: romout <= 16'h60DE;
32'hFFFF2F66: romout <= 16'h6100;
32'hFFFF2F68: romout <= 16'h006A;
32'hFFFF2F6A: romout <= 16'h5F0D;
32'hFFFF2F6C: romout <= 16'h103C;
32'hFFFF2F6E: romout <= 16'h000D;
32'hFFFF2F70: romout <= 16'h6100;
32'hFFFF2F72: romout <= 16'hF496;
32'hFFFF2F74: romout <= 16'h225F;
32'hFFFF2F76: romout <= 16'h60DE;
32'hFFFF2F78: romout <= 16'h4E75;
32'hFFFF2F7A: romout <= 16'h48E7;
32'hFFFF2F7C: romout <= 16'hC844;
32'hFFFF2F7E: romout <= 16'h4BF8;
32'hFFFF2F80: romout <= 16'h0700;
32'hFFFF2F82: romout <= 16'h2001;
32'hFFFF2F84: romout <= 16'h4EB9;
32'hFFFF2F86: romout <= 16'hFFFF;
32'hFFFF2F88: romout <= 16'h313E;
32'hFFFF2F8A: romout <= 16'h4BF8;
32'hFFFF2F8C: romout <= 16'h0700;
32'hFFFF2F8E: romout <= 16'h101D;
32'hFFFF2F90: romout <= 16'h6704;
32'hFFFF2F92: romout <= 16'h51CC;
32'hFFFF2F94: romout <= 16'hFFFA;
32'hFFFF2F96: romout <= 16'h4A44;
32'hFFFF2F98: romout <= 16'h6B0C;
32'hFFFF2F9A: romout <= 16'h103C;
32'hFFFF2F9C: romout <= 16'h0020;
32'hFFFF2F9E: romout <= 16'h6100;
32'hFFFF2FA0: romout <= 16'hF468;
32'hFFFF2FA2: romout <= 16'h51CC;
32'hFFFF2FA4: romout <= 16'hFFF2;
32'hFFFF2FA6: romout <= 16'h43F8;
32'hFFFF2FA8: romout <= 16'h0700;
32'hFFFF2FAA: romout <= 16'h4EB9;
32'hFFFF2FAC: romout <= 16'hFFFF;
32'hFFFF2FAE: romout <= 16'h1858;
32'hFFFF2FB0: romout <= 16'h4CDF;
32'hFFFF2FB2: romout <= 16'h2213;
32'hFFFF2FB4: romout <= 16'h4E75;
32'hFFFF2FB6: romout <= 16'h4281;
32'hFFFF2FB8: romout <= 16'h1219;
32'hFFFF2FBA: romout <= 16'hE189;
32'hFFFF2FBC: romout <= 16'h1219;
32'hFFFF2FBE: romout <= 16'h7805;
32'hFFFF2FC0: romout <= 16'h6100;
32'hFFFF2FC2: romout <= 16'hFFB8;
32'hFFFF2FC4: romout <= 16'h103C;
32'hFFFF2FC6: romout <= 16'h0020;
32'hFFFF2FC8: romout <= 16'h6100;
32'hFFFF2FCA: romout <= 16'hF43E;
32'hFFFF2FCC: romout <= 16'h4280;
32'hFFFF2FCE: romout <= 16'h6000;
32'hFFFF2FD0: romout <= 16'hFF4E;
32'hFFFF2FD2: romout <= 16'h6100;
32'hFFFF2FD4: romout <= 16'h0050;
32'hFFFF2FD6: romout <= 16'h225F;
32'hFFFF2FD8: romout <= 16'h1219;
32'hFFFF2FDA: romout <= 16'hB210;
32'hFFFF2FDC: romout <= 16'h6708;
32'hFFFF2FDE: romout <= 16'h4281;
32'hFFFF2FE0: romout <= 16'h1211;
32'hFFFF2FE2: romout <= 16'hD3C1;
32'hFFFF2FE4: romout <= 16'h4ED1;
32'hFFFF2FE6: romout <= 16'h5288;
32'hFFFF2FE8: romout <= 16'h5289;
32'hFFFF2FEA: romout <= 16'h4ED1;
32'hFFFF2FEC: romout <= 16'h4281;
32'hFFFF2FEE: romout <= 16'h4282;
32'hFFFF2FF0: romout <= 16'h6100;
32'hFFFF2FF2: romout <= 16'h0032;
32'hFFFF2FF4: romout <= 16'h0C10;
32'hFFFF2FF6: romout <= 16'h0030;
32'hFFFF2FF8: romout <= 16'h6528;
32'hFFFF2FFA: romout <= 16'h0C10;
32'hFFFF2FFC: romout <= 16'h0039;
32'hFFFF2FFE: romout <= 16'h6222;
32'hFFFF3000: romout <= 16'hB2BC;
32'hFFFF3002: romout <= 16'h0CCC;
32'hFFFF3004: romout <= 16'hCCCC;
32'hFFFF3006: romout <= 16'h6400;
32'hFFFF3008: romout <= 16'hFDE8;
32'hFFFF300A: romout <= 16'h2001;
32'hFFFF300C: romout <= 16'hD281;
32'hFFFF300E: romout <= 16'hD281;
32'hFFFF3010: romout <= 16'hD280;
32'hFFFF3012: romout <= 16'hD281;
32'hFFFF3014: romout <= 16'h1018;
32'hFFFF3016: romout <= 16'h0280;
32'hFFFF3018: romout <= 16'h0000;
32'hFFFF301A: romout <= 16'h000F;
32'hFFFF301C: romout <= 16'hD280;
32'hFFFF301E: romout <= 16'h5282;
32'hFFFF3020: romout <= 16'h60D2;
32'hFFFF3022: romout <= 16'h4E75;
32'hFFFF3024: romout <= 16'h0C10;
32'hFFFF3026: romout <= 16'h0020;
32'hFFFF3028: romout <= 16'h6604;
32'hFFFF302A: romout <= 16'h5288;
32'hFFFF302C: romout <= 16'h60F6;
32'hFFFF302E: romout <= 16'h4E75;
32'hFFFF3030: romout <= 16'h41F8;
32'hFFFF3032: romout <= 16'h0630;
32'hFFFF3034: romout <= 16'h4201;
32'hFFFF3036: romout <= 16'h1018;
32'hFFFF3038: romout <= 16'hB03C;
32'hFFFF303A: romout <= 16'h000D;
32'hFFFF303C: romout <= 16'h671A;
32'hFFFF303E: romout <= 16'hB03C;
32'hFFFF3040: romout <= 16'h0022;
32'hFFFF3042: romout <= 16'h6716;
32'hFFFF3044: romout <= 16'hB03C;
32'hFFFF3046: romout <= 16'h0027;
32'hFFFF3048: romout <= 16'h6710;
32'hFFFF304A: romout <= 16'h4A01;
32'hFFFF304C: romout <= 16'h66E8;
32'hFFFF304E: romout <= 16'h6100;
32'hFFFF3050: romout <= 16'h001A;
32'hFFFF3052: romout <= 16'h1100;
32'hFFFF3054: romout <= 16'h5288;
32'hFFFF3056: romout <= 16'h60DE;
32'hFFFF3058: romout <= 16'h4E75;
32'hFFFF305A: romout <= 16'h4A01;
32'hFFFF305C: romout <= 16'h6604;
32'hFFFF305E: romout <= 16'h1200;
32'hFFFF3060: romout <= 16'h60D4;
32'hFFFF3062: romout <= 16'hB200;
32'hFFFF3064: romout <= 16'h66D0;
32'hFFFF3066: romout <= 16'h4201;
32'hFFFF3068: romout <= 16'h60CC;
32'hFFFF306A: romout <= 16'hB03C;
32'hFFFF306C: romout <= 16'h0061;
32'hFFFF306E: romout <= 16'h650A;
32'hFFFF3070: romout <= 16'hB03C;
32'hFFFF3072: romout <= 16'h007A;
32'hFFFF3074: romout <= 16'h6204;
32'hFFFF3076: romout <= 16'h0400;
32'hFFFF3078: romout <= 16'h0020;
32'hFFFF307A: romout <= 16'h4E75;
32'hFFFF307C: romout <= 16'h6100;
32'hFFFF307E: romout <= 16'hF38E;
32'hFFFF3080: romout <= 16'h670A;
32'hFFFF3082: romout <= 16'hB03C;
32'hFFFF3084: romout <= 16'h0003;
32'hFFFF3086: romout <= 16'h6604;
32'hFFFF3088: romout <= 16'h6000;
32'hFFFF308A: romout <= 16'hF3D6;
32'hFFFF308C: romout <= 16'h4E75;
32'hFFFF308E: romout <= 16'h4DF9;
32'hFFFF3090: romout <= 16'hFFFF;
32'hFFFF3092: romout <= 16'h313A;
32'hFFFF3094: romout <= 16'h101E;
32'hFFFF3096: romout <= 16'h6706;
32'hFFFF3098: romout <= 16'h6100;
32'hFFFF309A: romout <= 16'hF36E;
32'hFFFF309C: romout <= 16'h60F6;
32'hFFFF309E: romout <= 16'h4E75;
32'hFFFF30A0: romout <= 16'h48E7;
32'hFFFF30A2: romout <= 16'hC000;
32'hFFFF30A4: romout <= 16'h2200;
32'hFFFF30A6: romout <= 16'h4EB9;
32'hFFFF30A8: romout <= 16'hFFFF;
32'hFFFF30AA: romout <= 16'h1732;
32'hFFFF30AC: romout <= 16'h4CDF;
32'hFFFF30AE: romout <= 16'h0003;
32'hFFFF30B0: romout <= 16'h4E75;
32'hFFFF30B2: romout <= 16'h3039;
32'hFFFF30B4: romout <= 16'hFFDC;
32'hFFFF30B6: romout <= 16'h0000;
32'hFFFF30B8: romout <= 16'h6A0C;
32'hFFFF30BA: romout <= 16'h4279;
32'hFFFF30BC: romout <= 16'hFFDC;
32'hFFFF30BE: romout <= 16'h0002;
32'hFFFF30C0: romout <= 16'h0240;
32'hFFFF30C2: romout <= 16'h00FF;
32'hFFFF30C4: romout <= 16'h4E75;
32'hFFFF30C6: romout <= 16'h7000;
32'hFFFF30C8: romout <= 16'h4E75;
32'hFFFF30CA: romout <= 16'h0839;
32'hFFFF30CC: romout <= 16'h0005;
32'hFFFF30CE: romout <= 16'hFFDC;
32'hFFFF30D0: romout <= 16'h0A01;
32'hFFFF30D2: romout <= 16'h67F6;
32'hFFFF30D4: romout <= 16'h13C0;
32'hFFFF30D6: romout <= 16'hFFDC;
32'hFFFF30D8: romout <= 16'h0A00;
32'hFFFF30DA: romout <= 16'h4E75;
32'hFFFF30DC: romout <= 16'h0839;
32'hFFFF30DE: romout <= 16'h0000;
32'hFFFF30E0: romout <= 16'hFFDC;
32'hFFFF30E2: romout <= 16'h0A01;
32'hFFFF30E4: romout <= 16'h670A;
32'hFFFF30E6: romout <= 16'h1039;
32'hFFFF30E8: romout <= 16'hFFDC;
32'hFFFF30EA: romout <= 16'h0A00;
32'hFFFF30EC: romout <= 16'h0200;
32'hFFFF30EE: romout <= 16'h007F;
32'hFFFF30F0: romout <= 16'h4E75;
32'hFFFF30F2: romout <= 16'h4EF9;
32'hFFFF30F4: romout <= 16'hFFFF;
32'hFFFF30F6: romout <= 16'h1A7A;
32'hFFFF30F8: romout <= 16'h0D0A;
32'hFFFF30FA: romout <= 16'h476F;
32'hFFFF30FC: romout <= 16'h7264;
32'hFFFF30FE: romout <= 16'h6F27;
32'hFFFF3100: romout <= 16'h7320;
32'hFFFF3102: romout <= 16'h4D43;
32'hFFFF3104: romout <= 16'h3638;
32'hFFFF3106: romout <= 16'h3030;
32'hFFFF3108: romout <= 16'h3020;
32'hFFFF310A: romout <= 16'h5469;
32'hFFFF310C: romout <= 16'h6E79;
32'hFFFF310E: romout <= 16'h2042;
32'hFFFF3110: romout <= 16'h4153;
32'hFFFF3112: romout <= 16'h4943;
32'hFFFF3114: romout <= 16'h2C20;
32'hFFFF3116: romout <= 16'h7631;
32'hFFFF3118: romout <= 16'h2E33;
32'hFFFF311A: romout <= 16'h0D0A;
32'hFFFF311C: romout <= 16'h0A00;
32'hFFFF311E: romout <= 16'h0D0A;
32'hFFFF3120: romout <= 16'h4F4B;
32'hFFFF3122: romout <= 16'h0D0A;
32'hFFFF3124: romout <= 16'h0048;
32'hFFFF3126: romout <= 16'h6F77;
32'hFFFF3128: romout <= 16'h3F0D;
32'hFFFF312A: romout <= 16'h0A00;
32'hFFFF312C: romout <= 16'h5768;
32'hFFFF312E: romout <= 16'h6174;
32'hFFFF3130: romout <= 16'h3F0D;
32'hFFFF3132: romout <= 16'h0A00;
32'hFFFF3134: romout <= 16'h536F;
32'hFFFF3136: romout <= 16'h7272;
32'hFFFF3138: romout <= 16'h792E;
32'hFFFF313A: romout <= 16'h0D0A;
32'hFFFF313C: romout <= 16'h00FF;
32'hFFFF313E: romout <= 16'h48E7;
32'hFFFF3140: romout <= 16'h7F00;
32'hFFFF3142: romout <= 16'h2E00;
32'hFFFF3144: romout <= 16'h6A08;
32'hFFFF3146: romout <= 16'h4487;
32'hFFFF3148: romout <= 16'h6B4E;
32'hFFFF314A: romout <= 16'h1AFC;
32'hFFFF314C: romout <= 16'h002D;
32'hFFFF314E: romout <= 16'h4244;
32'hFFFF3150: romout <= 16'h7C0A;
32'hFFFF3152: romout <= 16'h7401;
32'hFFFF3154: romout <= 16'h2206;
32'hFFFF3156: romout <= 16'h5381;
32'hFFFF3158: romout <= 16'h671A;
32'hFFFF315A: romout <= 16'h3602;
32'hFFFF315C: romout <= 16'hC6FC;
32'hFFFF315E: romout <= 16'h000A;
32'hFFFF3160: romout <= 16'h4842;
32'hFFFF3162: romout <= 16'hC4FC;
32'hFFFF3164: romout <= 16'h000A;
32'hFFFF3166: romout <= 16'h4843;
32'hFFFF3168: romout <= 16'hD443;
32'hFFFF316A: romout <= 16'h4842;
32'hFFFF316C: romout <= 16'h4843;
32'hFFFF316E: romout <= 16'h3403;
32'hFFFF3170: romout <= 16'h5381;
32'hFFFF3172: romout <= 16'h66E6;
32'hFFFF3174: romout <= 16'h4280;
32'hFFFF3176: romout <= 16'hBE82;
32'hFFFF3178: romout <= 16'h6D06;
32'hFFFF317A: romout <= 16'h5280;
32'hFFFF317C: romout <= 16'h9E82;
32'hFFFF317E: romout <= 16'h60F6;
32'hFFFF3180: romout <= 16'h4A00;
32'hFFFF3182: romout <= 16'h6604;
32'hFFFF3184: romout <= 16'h4A44;
32'hFFFF3186: romout <= 16'h6708;
32'hFFFF3188: romout <= 16'h0600;
32'hFFFF318A: romout <= 16'h0030;
32'hFFFF318C: romout <= 16'h1AC0;
32'hFFFF318E: romout <= 16'h1800;
32'hFFFF3190: romout <= 16'h5386;
32'hFFFF3192: romout <= 16'h66BE;
32'hFFFF3194: romout <= 16'h4A44;
32'hFFFF3196: romout <= 16'h6604;
32'hFFFF3198: romout <= 16'h1AFC;
32'hFFFF319A: romout <= 16'h0030;
32'hFFFF319C: romout <= 16'h1ABC;
32'hFFFF319E: romout <= 16'h0000;
32'hFFFF31A0: romout <= 16'h4CDF;
32'hFFFF31A2: romout <= 16'h00FE;
32'hFFFF31A4: romout <= 16'h4E75;
default: romout <= 16'h0000;
endcase
always @(posedge clk)
    romo <= romout;
endmodule
