`include "mips789_defs.v"

module mips_core (
        clk,rst,zz_ins_i,iack_o,qa,qb,wb_din_o,rdaddra_o,rdaddrb_o,wb_addr_o,wb_we_o,
       zz_pc_o,dmem_ctl_ur_o,alu_ur_o,dmem_data_ur_o,dout,size,branch,hold,imds,dmds,asi_pass2, pc_next
    );

    input clk;
    wire clk;
    input rst;
    wire rst;
    input [31:0] zz_ins_i;
    wire [31:0] zz_ins_i;
	 wire [31:0] zz_ins_o; 
    input [31:0] dout;
    wire [31:0] dout;
	 input [31:0] qa;
	 wire [31:0] qa;
	 input [31:0] qb;
	 wire [31:0] qb;
    output [31:0] zz_pc_o;
    wire [31:0] zz_pc_o;
    output iack_o;
    wire iack_o;
    wire [31:0] cop_addr_o;
    output [4:0] dmem_ctl_ur_o;
    output [31:0] alu_ur_o;
    output [31:0] dmem_data_ur_o;
    wire [4:0] dmem_ctl_ur_o;
    wire [31:0] alu_ur_o;
    wire [31:0] dmem_data_ur_o;
	 output [31:0] wb_din_o;
	 wire [31:0] wb_din_o;
	 output [4:0] rdaddra_o;
	 wire [4:0] rdaddra_o;
	 output [4:0] rdaddrb_o;
	 wire [4:0] rdaddrb_o;
	 output [4:0] wb_addr_o;
	 wire [4:0] wb_addr_o;
	 output wb_we_o;
	 wire wb_we_o;
	 output [1:0] size;
	 wire [1:0] size;
	 output branch;
	 wire branch;
	 input hold;
	 wire hold;
	 input imds;
	 wire imds;
	 input dmds;
	 wire dmds;
	 output [4:0] asi_pass2;
	 output [31:0] pc_next;
	 
	 wire [31:0] pc_next;
    wire load;
	 wire load_o;
	 wire [4:0]rt_o;
    wire NET1375;
    wire NET1572;
    wire NET1606;
    wire NET1640;
    wire NET21531;
    wire NET457;
    wire NET767;
    wire [2:0] BUS109;
    wire [2:0] BUS1158;
    wire [2:0] BUS117;
    wire [2:0] BUS1196;
    wire [31:0] BUS15471;
    wire [4:0] BUS1724;
    wire [4:0] BUS1726;
    wire [4:0] BUS18211;
    wire [2:0] BUS197;
    wire [2:0] BUS2140;
    wire [2:0] BUS2156;
    wire [31:0] BUS22401;
    wire [31:0] BUS24839;
    wire [31:0] BUS27031;
    wire [2:0] BUS271;
    wire [31:0] BUS28013;
    wire [1:0] BUS371;
    wire [31:0] BUS422;
    wire [1:0] BUS5832;
    wire [1:0] BUS5840;
    wire [2:0] BUS5993;
    wire [4:0] BUS6275;
    wire [31:0] BUS7101;
    wire [31:0] BUS7117;
    wire [31:0] BUS7160;
    wire [31:0] BUS7219;
    wire [31:0] BUS7231;
    wire [4:0] BUS748;
    wire [4:0] BUS756;
    wire [4:0] BUS775;
    wire [31:0] BUS7772;
    wire [31:0] BUS7780;
    wire [31:0] BUS9884;
	 wire [4:0] asi_o;
	 wire [4:0] asi_pass1;
	 wire [4:0] asi_pass2;
	 wire [4:0] rdaddra1;
	 wire [4:0] rdaddrb1;
	 
	

    assign NET21531 = NET1572 | iack_o;

    rf_stage iRF_stage
             (   .hold(hold),
                 .clk(clk),
                 .cmp_ctl_i(BUS109),
                 .ext_ctl_i(BUS117),
                 .ext_o(BUS7219),
                 .fw_alu_i(cop_addr_o),
                 .fw_cmp_rs(BUS2140),
                 .fw_cmp_rt(BUS2156),
                 .fw_mem_i(wb_din_o),
                 .iack_o(iack_o),
                 .id2ra_ctl_clr_o(NET1606),
                 .id2ra_ctl_cls_o(NET1572),
                 .id_cmd(BUS197),
                 .ins_i(zz_ins_o),
                 .pc_gen_ctl(BUS271),
					  .branch(branch),
                 .pc_i(zz_pc_o),
                 .pc_next(pc_next),
                 .ra2ex_ctl_clr_o(NET1640),
                 .rd_index_o(BUS775),
                 .rd_sel_i(BUS371),
                 .rs_n_o(BUS748),
                 .rs_o(BUS24839),
                 .rst_i(rst),
                 .rt_n_o(BUS756),
                 .rt_o(BUS7160),
                 .wb_din_i(wb_din_o),
                 .zz_spc_i(BUS28013),
					  .rdaddra1(rdaddra1),
					  .rdaddrb1(rdaddrb1),
					  .qa(qa),
					  .qb(qb)
             );



    exec_stage iexec_stage
               (.hold(hold),
                   .alu_func(BUS6275),
                   .alu_ur_o(alu_ur_o),
                   .clk(clk),
                   .dmem_data_ur_o(dmem_data_ur_o),
                   .dmem_fw_ctl(BUS5993),
                   .ext_i(BUS7231),
                   .fw_alu(cop_addr_o),
                   .fw_dmem(wb_din_o),
                   .muxa_ctl_i(BUS5832),
                   .muxa_fw_ctl(BUS1158),
                   .muxb_ctl_i(BUS5840),
                   .muxb_fw_ctl(BUS1196),
                   .pc_i(zz_pc_o),
                   .rs_i(BUS7101),
                   .rst(rst),
                   .rt_i(BUS7117),
                   .spc_cls_i(NET21531),
                   .zz_spc_o(BUS28013)
               );



    r32_reg alu_pass0
            (.hold(hold),
                .clk(clk),
                .r32_i(alu_ur_o),
                .r32_o(cop_addr_o)
            );



    r32_reg alu_pass1
            (.hold(hold),
                .clk(clk),
                .r32_i(cop_addr_o),
                .r32_o(BUS422)
            );
	
	r32_inst_reg instruction
            (	 .hold(hold),
					 .branch(branch),
					 .imds(imds),
                .clk(clk),
                .r32_i(zz_ins_i),
                .r32_o(zz_ins_o)
            );



//    or32 cop_data_or
//         (
//             .a(cop_dout),
//             .b(BUS7772),
//             .c(BUS7780)
//         );



//    r32_reg cop_data_reg
//            (
//                .clk(clk),
//                .r32_i(BUS9884),
//                .r32_o(cop_data_o)
//            );



/*    r32_reg cop_dout_reg
            (.hold(hold),
                .clk(clk),
                .r32_i(dout),
                .r32_o(BUS7780)
            );
	*/
	
	r32_data_reg cop_dout_reg
            (	 .hold(hold),
					 .dmds(dmds),
                .clk(clk),
                .r32_i(dout),
                .r32_o(BUS7780)
            );



    decode_pipe decoder_pipe
                (.hold(hold),
						  .rt1(rt_o),
						  .load(load_o),
						  .load_o(load),
                    .alu_func_o(BUS6275),
						  .size(size),
                    .alu_we_o(NET767),
                    .clk(clk),
                    .cmp_ctl_o(BUS109),
                    .dmem_ctl_ur_o(dmem_ctl_ur_o),
                    .ext_ctl_o(BUS117),
                    .fsm_dly(BUS197),
                    .id2ra_ctl_clr(NET1606),
                    .id2ra_ctl_cls(NET1572),
                    .ins_i(zz_ins_o),
                    .muxa_ctl_o(BUS5832),
                    .muxb_ctl_o(BUS5840),
                    .pc_gen_ctl_o(BUS271),
                    .ra2ex_ctl_clr(NET1640),
                    .rd_sel_o(BUS371),
                    .wb_mux_ctl_o(NET457),
                    .wb_we_o(wb_we_o),
						  .asi(asi_o)
                );



    r32_reg ext_reg
            (.hold(hold),
                .clk(clk),
                .r32_i(BUS7219),
                .r32_o(BUS7231)
            );



    forward iforward
            (.hold(hold),
                .alu_rs_fw(BUS1158),
                .alu_rt_fw(BUS1196),
                .alu_we(NET767),
                .clk(clk),
                .cmp_rs_fw(BUS2140),
                .cmp_rt_fw(BUS2156),
                .dmem_fw(BUS5993),
                .fw_alu_rn(BUS1724),
                .fw_mem_rn(wb_addr_o),
                .mem_We(wb_we_o),
                .rns_i(BUS748),
                .rnt_i(BUS756)
            );



    r32_reg pc
            (.hold(hold),
                .clk(clk),
                .r32_i(pc_next),
                .r32_o(zz_pc_o)
            );



    r5_reg rnd_pass0
           (.hold(hold),
               .clk(clk),
               .r5_i(BUS775),
               .r5_o(BUS1726)
           );



    r5_reg rnd_pass1
           (.hold(hold),
               .clk(clk),
               .r5_i(BUS1726),
               .r5_o(BUS1724)
           );



    r5_reg rnd_pass2
           (.hold(hold),
               .clk(clk),
               .r5_i(BUS1724),
               .r5_o(wb_addr_o)
           );



    r32_reg rs_reg
            (.hold(hold),
                .clk(clk),
                .r32_i(BUS24839),
                .r32_o(BUS7101)
            );



    r32_reg rt_reg
            (.hold(hold),
                .clk(clk),
                .r32_i(BUS7160),
                .r32_o(BUS7117)
            );



    wb_mux wb_mux
           (
               .alu_i(BUS422),
               .dmem_i(BUS7780),
               .sel(NET457),
               .wb_o(wb_din_o)
           );
			  
	 hazard_unit ihazard_unit
			(.hold(hold),
					.clk(clk),
					.rt(rdaddrb_o),
					.load(load),
					.load_o(load_o),
					.rt_o(rt_o)
			);  
			
			r4_asi_reg reg_asi_pass1
            (	 .hold(hold),
                .clk(clk),
                .r4_i(asi_o),
                .r4_o(asi_pass1)
            );
				
			r4_asi_reg reg_asi_pass2
            (	 .hold(hold),
                .clk(clk),
                .r4_i(asi_pass1),
                .r4_o(asi_pass2)
            );

			r4_rdaddr_reg reg_rdaddra
            (	 .hold(hold),
                .clk(clk),
                .clr(NET1606),
                .cls(NET1572),
                .r4_i(rdaddra1),
                .r4_o(rdaddra_o)
            );
				
				r4_rdaddr_reg reg_rdaddrb
            (	 .hold(hold),
                .clk(clk),
                .clr(NET1606),
                .cls(NET1572),
                .r4_i(rdaddrb1),
                .r4_o(rdaddrb_o)
            );
			
			
endmodule
