-------------------------------------------------------------------------------
--
-- SD/MMC Bootloader
--
-- $Id: card-c.vhd 77 2009-04-01 19:53:14Z arniml $
--
-------------------------------------------------------------------------------

configuration card_behav_c0 of card is

  for behav
  end for;

end card_behav_c0;
