-- DSU UART
  constant CFG_AHB_UART	: integer := CONFIG_DSU_UART;

