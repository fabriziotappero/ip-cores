library ieee;
use ieee.std_logic_1164.all;

package asci_types is
  type lcd_char is (
    NUL, SOH, STX, ETX, EOT, ENQ, ACK, BEL, 
    BS,  HT,  LF,  VT,  FF,  CR,  SO,  SI,
    DLE, DC1, DC2, DC3, DC4, NAK, SYN, ETB, 
    CAN,  EM, SUB, ESC, FSP, GSP, RSP, USP,
    ' ', '!', '"', '#', '$', '%', '&', ''',
    '(', ')', '*', '+', ',', '-', '.', '/', 
    '0', '1', '2', '3', '4', '5', '6', '7', 
    '8', '9', ':', ';', '<', '=', '>', '?', 
    '@', 'A', 'B', 'C', 'D', 'E', 'F', 'G',
    'H', 'I', 'J', 'K', 'L', 'M', 'N', 'O', 
    'P', 'Q', 'R', 'S', 'T', 'U', 'V', 'W', 
    'X', 'Y', 'Z', '[', '\', ']', '^', '_', 
    '`', 'a', 'b', 'c', 'd', 'e', 'f', 'g', 
    'h', 'i', 'j', 'k', 'l', 'm', 'n', 'o', 
    'p', 'q', 'r', 's', 't', 'u', 'v', 'w', 
    'x', 'y', 'z', '{', '|', '}', '~', DEL );
  type lcd_matrix is array(natural range 1 TO 80) of lcd_char;
  TYPE char_std_matrix IS array(lcd_char RANGE NUL TO DEL) OF std_logic_vector(7 DOWNTO 0);
  constant char2std : char_std_matrix :=
    ("00000000", "00000001", "00000010", "00000011",
     "00000100", "00000101", "00000110", "00000111",
     "00001000", "00001001", "00001010", "00001011",
     "00001100", "00001101", "10010001", "00001111",
     "00010000", "00010001", "00010010", "00010011",
     "10110110", "01011111", "00010110", "00010111",
     "11011110", "11100000", "11010000", "11100001",
     "00011100", "00011101", "00011110", "00011111",
     "00100000", "00100001", "00100010", "00100011",
     "10100010", "00100101", "00100110", "00100111",
     "00101000", "00101001", "00101010", "00101011",
     "00101100", "00101101", "00101110", "00101111",
     "00110000", "00110001", "00110010", "00110011",
     "00110100", "00110101", "00110110", "00110111",
     "00111000", "00111001", "00111010", "00111011",
     "00111100", "00111101", "00111110", "00111111",
     "10100000", "01000001", "01000010", "01000011",
     "01000100", "01000101", "01000110", "01000111",
     "01001000", "01001001", "01001010", "01001011",
     "01001100", "01001101", "01001110", "01001111",
     "01010000", "01010001", "01010010", "01010011",
     "01010100", "01010101", "01010110", "01010111",
     "01011000", "01011001", "01011010", "11111010",
     "11111011", "11111100", "00011101", "11000100",
     "00100111", "01100001", "01100010", "01100011",
     "01100100", "01100101", "01100110", "01100111",
     "01101000", "01101001", "01101010", "01101011",
     "01101100", "01101101", "01101110", "01101111",
     "01110000", "01110001", "01110010", "01110011",
     "01110100", "01110101", "01110110", "01110111",
     "01111000", "01111001", "01111010", "11111101",
     "11111110", "11111111", "11001110", "10110000");
END asci_types;
  
  
