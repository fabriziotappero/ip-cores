-- USB Host Controller
  constant CFG_GRUSBHC          : integer := CONFIG_GRUSBHC_ENABLE;
  constant CFG_GRUSBHC_NPORTS   : integer := CONFIG_GRUSBHC_NPORTS;
  constant CFG_GRUSBHC_EHC      : integer := CONFIG_GRUSBHC_EHC;
  constant CFG_GRUSBHC_UHC      : integer := CONFIG_GRUSBHC_UHC;
  constant CFG_GRUSBHC_NCC      : integer := CONFIG_GRUSBHC_NCC;
  constant CFG_GRUSBHC_NPCC     : integer := CONFIG_GRUSBHC_NPCC;
  constant CFG_GRUSBHC_PRR      : integer := CONFIG_GRUSBHC_PRR;
  constant CFG_GRUSBHC_PR1      : integer := CONFIG_GRUSBHC_PORTROUTE1;
  constant CFG_GRUSBHC_PR2      : integer := CONFIG_GRUSBHC_PORTROUTE2;
  constant CFG_GRUSBHC_ENDIAN   : integer := CONFIG_GRUSBHC_ENDIAN;
  constant CFG_GRUSBHC_BEREGS   : integer := CONFIG_GRUSBHC_BEREGS;
  constant CFG_GRUSBHC_BEDESC   : integer := CONFIG_GRUSBHC_BEDESC;
  constant CFG_GRUSBHC_BLO      : integer := CONFIG_GRUSBHC_BLO;
  constant CFG_GRUSBHC_BWRD     : integer := CONFIG_GRUSBHC_BWRD;
  constant CFG_GRUSBHC_UTM      : integer := CONFIG_GRUSBHC_UTMTYPE;
  constant CFG_GRUSBHC_VBUSCONF : integer := CONFIG_GRUSBHC_VBUSCONF;

