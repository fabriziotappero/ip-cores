000000 => x"cafe",
000001 => x"0017",
000002 => x"aa75",
000003 => x"424c",
000004 => x"494e",
000005 => x"4b5f",
000006 => x"4445",
000007 => x"4d4f",
000008 => x"bc05",
000009 => x"bc00",
000010 => x"bc00",
000011 => x"bc00",
000012 => x"bc00",
000013 => x"2800",
000014 => x"ed0f",
000015 => x"c2b2",
000016 => x"be09",
000017 => x"ed0f",
000018 => x"3c00",
000019 => x"0001",
000020 => x"c08f",
000021 => x"2001",
000022 => x"3c00",
000023 => x"ed0f",
000024 => x"bdf7",
000025 => x"c77f",
000026 => x"0769",
000027 => x"85ff",
000028 => x"06d9",
000029 => x"85fc",
000030 => x"3470",
others => x"0000"