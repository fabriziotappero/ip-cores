// --------------------------------------------------------------------
//
// --------------------------------------------------------------------


`timescale 1ps/1ps


module tb_top();

  // --------------------------------------------------------------------
  // system wires
  wire CLK_20;
  wire CLK_50;
  wire CLK_100;
  wire CLK_125;
  wire CLK_156_25;

  wire tb_clk = CLK_50;

  wire tb_rst;


  // --------------------------------------------------------------------
  // clock & reset
  parameter CLK_PERIOD = 2000;

  tb_clk #( .CLK_PERIOD(5000) ) i_CLK_20    ( CLK_20 );
  tb_clk #( .CLK_PERIOD(2000) ) i_CLK_50    ( CLK_50 );
  tb_clk #( .CLK_PERIOD(1000) ) i_CLK_100   ( CLK_100 );
  tb_clk #( .CLK_PERIOD(640) ) i_CLK_156_25 ( CLK_156_25 );
  tb_clk #( .CLK_PERIOD(800) ) i_CLK_125    ( CLK_125 );

  tb_reset #( .ASSERT_TIME(CLK_PERIOD*10) ) i_tb_rst( tb_rst );

  initial
    begin
      $display("\n^^^---------------------------------");
      i_tb_rst.assert_delayed_reset(CLK_PERIOD/3);
    end
    

  // --------------------------------------------------------------------
  //



  // --------------------------------------------------------------------
  // sim models
  //  |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   | 
  // \|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/-\|/
  //  '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   ' 



  // --------------------------------------------------------------------
  //
  tb_log log();
  

  //  '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   '   ' 
  // /|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\-/|\
  //  |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   |   | 
  // sim models 
  // --------------------------------------------------------------------


  // --------------------------------------------------------------------
  //  debug wires



  // --------------------------------------------------------------------
  // test
  the_test test( tb_clk, tb_rst );

  initial
    begin

      test.run_the_test();

      $display("^^^---------------------------------");
      $display("^^^ %16.t | Testbench done.", $time);
      $display("^^^---------------------------------");

      log.log_fail_count();
      $display("^^^---------------------------------");

`ifdef MAKEFILE_TEST_RUN
      $finish();
`else
      $stop();
`endif

    end

endmodule



