-- ------------------------------------------------------------------------
-- Copyright (C) 2005 Arif Endro Nugroho
-- All rights reserved.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY ARIF ENDRO NUGROHO "AS IS" AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL ARIF ENDRO NUGROHO BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
-- ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
-- POSSIBILITY OF SUCH DAMAGE.
-- 
-- End Of License.
-- ------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity reference is
   port (
      clear    : in  bit;
      start    : in  bit;
      y0       : in  bit;
      y1       : in  bit;
      y2       : in  bit;
      y3       : in  bit;
      senddata : out bit_vector (3 downto 0);
      match    : out bit_vector (3 downto 0)
      );
end reference;

architecture verify of reference is

type senddata_rom is array (000 to 2499) of bit_vector (3 downto 0);
constant senddata_tbl : senddata_rom :=
(

 B"0010", B"0001", B"1101", B"1011", 
 B"1000", B"1011", B"1101", B"1100", 
 B"0010", B"0011", B"1100", B"1010", 
 B"1001", B"1111", B"0110", B"0010", 
 B"1100", B"1000", B"0001", B"1010", 
 B"0110", B"1011", B"0101", B"0001", 
 B"1100", B"1001", B"1100", B"1000", 
 B"0110", B"1101", B"0000", B"0100", 
 B"0000", B"0110", B"1101", B"1011", 
 B"0000", B"1001", B"1001", B"1000", 
 B"0110", B"1100", B"0110", B"1101", 
 B"1101", B"1011", B"0101", B"1101", 
 B"1111", B"0110", B"1000", B"0010", 
 B"1111", B"0110", B"0000", B"1110", 
 B"0001", B"0101", B"0111", B"1111", 
 B"0100", B"1010", B"1011", B"0111", 
 B"0011", B"1101", B"1000", B"1000", 
 B"0001", B"1000", B"1110", B"0110", 
 B"1111", B"1101", B"0000", B"0000", 
 B"1111", B"1010", B"1001", B"0011", 
 B"1110", B"0010", B"0010", B"0011", 
 B"1000", B"1101", B"1101", B"0000", 
 B"0000", B"1001", B"1010", B"1010", 
 B"0000", B"0111", B"0001", B"1111", 
 B"1010", B"0110", B"0100", B"0000", 
 B"1011", B"1100", B"0000", B"0011", 
 B"1111", B"0001", B"0000", B"0000", 
 B"1011", B"0100", B"1101", B"0011", 
 B"0001", B"1000", B"0101", B"0000", 
 B"0100", B"1111", B"0100", B"0010", 
 B"0101", B"0000", B"0001", B"0100", 
 B"1000", B"0000", B"1101", B"1100", 
 B"1110", B"1100", B"1001", B"0010", 
 B"0101", B"0001", B"0101", B"1001", 
 B"0011", B"1010", B"0111", B"1101", 
 B"0010", B"1111", B"1010", B"0011", 
 B"0011", B"0010", B"0111", B"0010", 
 B"0000", B"0001", B"0110", B"1100", 
 B"0001", B"0110", B"1110", B"0110", 
 B"1101", B"0001", B"1101", B"0001", 
 B"0011", B"1000", B"1001", B"1010", 
 B"0110", B"1101", B"0110", B"1010", 
 B"0011", B"0010", B"1110", B"1101", 
 B"1011", B"0010", B"1110", B"1000", 
 B"0010", B"1111", B"0010", B"0110", 
 B"1110", B"1100", B"0000", B"0000", 
 B"0000", B"0110", B"1110", B"0101", 
 B"1010", B"1000", B"0100", B"0001", 
 B"0101", B"0110", B"1101", B"1011", 
 B"1000", B"1111", B"1111", B"1101", 
 B"0001", B"1011", B"1000", B"0011", 
 B"0010", B"0100", B"0010", B"0010", 
 B"0010", B"0101", B"0111", B"1101", 
 B"1000", B"1101", B"1001", B"1001", 
 B"0101", B"0011", B"0100", B"0000", 
 B"1100", B"1100", B"1000", B"1001", 
 B"0000", B"1110", B"0110", B"1101", 
 B"0010", B"0000", B"1111", B"1010", 
 B"1010", B"0100", B"1101", B"0010", 
 B"1001", B"1001", B"1011", B"1000", 
 B"0000", B"1001", B"1110", B"0000", 
 B"0110", B"1000", B"0101", B"0010", 
 B"1100", B"0100", B"1000", B"0110", 
 B"0100", B"1111", B"0011", B"0101", 
 B"0000", B"1100", B"0110", B"1110", 
 B"1111", B"1000", B"1000", B"0110", 
 B"1000", B"1000", B"1100", B"1000", 
 B"1100", B"0011", B"0110", B"1001", 
 B"0101", B"0011", B"0111", B"0100", 
 B"0010", B"1011", B"1001", B"0111", 
 B"1110", B"0001", B"1001", B"0110", 
 B"1001", B"0111", B"1111", B"0010", 
 B"1010", B"0011", B"0101", B"1010", 
 B"0000", B"0000", B"0001", B"0110", 
 B"1111", B"0010", B"0100", B"1100", 
 B"0100", B"0001", B"0000", B"1010", 
 B"1001", B"1011", B"0101", B"1101", 
 B"1100", B"1010", B"0010", B"1101", 
 B"1111", B"1000", B"0111", B"0101", 
 B"0010", B"1101", B"0111", B"1110", 
 B"1011", B"0110", B"0101", B"1010", 
 B"1001", B"0001", B"0001", B"1000", 
 B"0100", B"1010", B"1111", B"1100", 
 B"1000", B"0101", B"1010", B"0011", 
 B"0010", B"1010", B"1010", B"0110", 
 B"0101", B"0000", B"0011", B"0011", 
 B"0110", B"0011", B"1100", B"1111", 
 B"0001", B"1101", B"1011", B"1111", 
 B"1100", B"1000", B"0010", B"1100", 
 B"0010", B"1100", B"0001", B"1101", 
 B"0111", B"0001", B"1110", B"1010", 
 B"0010", B"1111", B"0101", B"1011", 
 B"1110", B"0001", B"0001", B"1000", 
 B"1000", B"1000", B"1011", B"0101", 
 B"1000", B"1011", B"0011", B"0001", 
 B"1110", B"1111", B"0111", B"0010", 
 B"0101", B"0110", B"0000", B"1110", 
 B"0000", B"0110", B"1011", B"0101", 
 B"0001", B"0001", B"1111", B"1100", 
 B"1110", B"0000", B"0101", B"1011", 
 B"1011", B"0000", B"0110", B"0111", 
 B"0111", B"1110", B"0011", B"0000", 
 B"1100", B"0110", B"0000", B"1000", 
 B"0010", B"0100", B"1101", B"0000", 
 B"0000", B"0001", B"0100", B"1101", 
 B"0011", B"1001", B"0110", B"1001", 
 B"0000", B"0000", B"0001", B"1011", 
 B"1000", B"1001", B"0000", B"1000", 
 B"1101", B"0111", B"0110", B"0100", 
 B"1011", B"0010", B"0000", B"0100", 
 B"1010", B"1101", B"1011", B"1100", 
 B"0111", B"1111", B"0110", B"0011", 
 B"0001", B"0100", B"0001", B"1010", 
 B"1011", B"0110", B"1111", B"1010", 
 B"1110", B"0010", B"1000", B"0100", 
 B"0010", B"1010", B"1010", B"1010", 
 B"0001", B"1010", B"0000", B"1010", 
 B"0101", B"1011", B"0000", B"0100", 
 B"1000", B"1111", B"0100", B"1010", 
 B"1111", B"1000", B"1110", B"0111", 
 B"1110", B"1011", B"0000", B"1100", 
 B"0011", B"0000", B"1011", B"1100", 
 B"0010", B"1000", B"1011", B"0110", 
 B"1000", B"1111", B"1000", B"0110", 
 B"1100", B"1001", B"1101", B"1001", 
 B"0010", B"0100", B"0101", B"0101", 
 B"1010", B"0000", B"1000", B"1010", 
 B"1100", B"0110", B"0110", B"1100", 
 B"0011", B"0010", B"0000", B"0100", 
 B"0010", B"1010", B"1010", B"0101", 
 B"0110", B"1000", B"0001", B"0100", 
 B"1111", B"0011", B"0111", B"1001", 
 B"0111", B"0110", B"1100", B"1010", 
 B"1001", B"0011", B"0000", B"0010", 
 B"0110", B"0000", B"1100", B"1101", 
 B"0100", B"0010", B"1110", B"0011", 
 B"0001", B"1011", B"0000", B"1010", 
 B"0011", B"0011", B"0111", B"0100", 
 B"0001", B"1100", B"1000", B"1101", 
 B"0100", B"1101", B"0010", B"1011", 
 B"1010", B"1011", B"0011", B"1000", 
 B"1000", B"0010", B"1010", B"0010", 
 B"0110", B"1100", B"1110", B"0010", 
 B"0110", B"0001", B"0111", B"1101", 
 B"1101", B"1111", B"0010", B"0001", 
 B"0011", B"0110", B"0100", B"0101", 
 B"1001", B"0011", B"0000", B"0101", 
 B"1111", B"0010", B"1110", B"1010", 
 B"1111", B"0011", B"1101", B"0011", 
 B"0000", B"0101", B"0011", B"0100", 
 B"0101", B"0111", B"1100", B"0101", 
 B"0010", B"1101", B"0010", B"1100", 
 B"1110", B"1110", B"0011", B"0101", 
 B"1001", B"0111", B"0001", B"0011", 
 B"1000", B"0010", B"0001", B"1000", 
 B"1010", B"0110", B"0101", B"0010", 
 B"0101", B"0010", B"1011", B"1111", 
 B"1110", B"0100", B"0110", B"1001", 
 B"0110", B"0111", B"0111", B"1000", 
 B"0001", B"0111", B"1101", B"1110", 
 B"1011", B"1111", B"0010", B"0100", 
 B"1110", B"0111", B"0000", B"1011", 
 B"0001", B"0010", B"0000", B"1011", 
 B"0000", B"0101", B"0001", B"1111", 
 B"0000", B"1101", B"1101", B"0010", 
 B"1011", B"1110", B"1110", B"0001", 
 B"0010", B"1011", B"0011", B"1101", 
 B"0101", B"1011", B"1100", B"1100", 
 B"1001", B"0101", B"0000", B"0111", 
 B"1111", B"1000", B"0010", B"0100", 
 B"1100", B"1001", B"0111", B"1001", 
 B"0101", B"0000", B"1110", B"1000", 
 B"1011", B"0111", B"0101", B"1001", 
 B"0101", B"0000", B"1100", B"0111", 
 B"1001", B"1110", B"1001", B"1011", 
 B"1010", B"0011", B"1101", B"1101", 
 B"0101", B"0101", B"1110", B"1011", 
 B"1011", B"1101", B"0111", B"0101", 
 B"1010", B"1101", B"1101", B"1000", 
 B"1101", B"0001", B"1110", B"0101", 
 B"0100", B"0001", B"0010", B"1011", 
 B"1001", B"1001", B"1110", B"1101", 
 B"0101", B"0110", B"0001", B"1101", 
 B"0011", B"0111", B"0110", B"0001", 
 B"0011", B"1111", B"0101", B"1101", 
 B"1111", B"0000", B"1000", B"1001", 
 B"1111", B"1100", B"0110", B"0001", 
 B"1100", B"1010", B"1111", B"0011", 
 B"1000", B"0100", B"1101", B"0100", 
 B"0100", B"0111", B"1011", B"1110", 
 B"0101", B"0101", B"1011", B"1001", 
 B"0001", B"0110", B"0110", B"1111", 
 B"1110", B"1100", B"1100", B"1011", 
 B"1000", B"1010", B"1100", B"1001", 
 B"0101", B"0010", B"0010", B"0011", 
 B"1001", B"0010", B"0010", B"0111", 
 B"1111", B"0100", B"0001", B"0000", 
 B"1001", B"1100", B"0010", B"1010", 
 B"0100", B"0110", B"0010", B"0001", 
 B"1111", B"0100", B"0001", B"0101", 
 B"0001", B"0010", B"0111", B"0010", 
 B"1110", B"0100", B"0001", B"1100", 
 B"0111", B"1100", B"1010", B"0011", 
 B"1010", B"1110", B"0100", B"0101", 
 B"0001", B"0000", B"0100", B"1000", 
 B"1001", B"0010", B"0100", B"0000", 
 B"0011", B"1111", B"1010", B"0010", 
 B"0110", B"0111", B"1110", B"0101", 
 B"1111", B"0110", B"0010", B"0011", 
 B"1101", B"0001", B"1000", B"1101", 
 B"0001", B"1111", B"1110", B"1111", 
 B"1011", B"1100", B"0001", B"0001", 
 B"1111", B"0000", B"1000", B"0000", 
 B"1111", B"1110", B"0011", B"0110", 
 B"1000", B"0101", B"0100", B"1000", 
 B"0001", B"0001", B"1001", B"0100", 
 B"1000", B"1101", B"1100", B"0000", 
 B"1101", B"1111", B"1011", B"1011", 
 B"1110", B"1100", B"0010", B"0111", 
 B"0000", B"0000", B"1101", B"1101", 
 B"0010", B"0000", B"1000", B"0100", 
 B"1001", B"1001", B"1111", B"1001", 
 B"0001", B"1110", B"1110", B"1111", 
 B"0111", B"1010", B"0000", B"1100", 
 B"0111", B"1110", B"1010", B"0100", 
 B"0100", B"0010", B"1101", B"0000", 
 B"1100", B"0011", B"1100", B"0011", 
 B"0010", B"1001", B"0010", B"1011", 
 B"0110", B"1010", B"1011", B"1110", 
 B"0001", B"0110", B"1001", B"0000", 
 B"1111", B"0100", B"0100", B"0011", 
 B"1101", B"0110", B"1101", B"0101", 
 B"0001", B"1100", B"1101", B"0100", 
 B"0001", B"1110", B"0011", B"1101", 
 B"1101", B"0000", B"1110", B"0010", 
 B"1001", B"0110", B"1000", B"0000", 
 B"1000", B"1010", B"1011", B"1000", 
 B"0110", B"0010", B"1010", B"1111", 
 B"1000", B"0011", B"1010", B"0000", 
 B"0010", B"1011", B"1110", B"1000", 
 B"0011", B"0100", B"0101", B"1001", 
 B"0100", B"0111", B"1110", B"0111", 
 B"0011", B"0111", B"0100", B"1100", 
 B"1010", B"0110", B"1011", B"1111", 
 B"1110", B"1011", B"0111", B"1110", 
 B"0011", B"0011", B"0011", B"0001", 
 B"0110", B"1110", B"1000", B"0000", 
 B"1100", B"0001", B"0100", B"0001", 
 B"0010", B"1001", B"0011", B"0100", 
 B"0011", B"0011", B"0111", B"1001", 
 B"1111", B"1101", B"0000", B"0000", 
 B"1010", B"0000", B"0110", B"0110", 
 B"0001", B"1100", B"1111", B"1100", 
 B"0000", B"1001", B"1101", B"0001", 
 B"1001", B"0101", B"0101", B"0101", 
 B"1000", B"0101", B"0001", B"1100", 
 B"1111", B"1111", B"1000", B"1110", 
 B"1000", B"0101", B"0011", B"1111", 
 B"0110", B"1001", B"1010", B"0011", 
 B"1101", B"1011", B"0010", B"1100", 
 B"0000", B"0101", B"0000", B"0011", 
 B"1110", B"1001", B"0111", B"0110", 
 B"0110", B"0011", B"1010", B"0000", 
 B"1000", B"0111", B"0111", B"1101", 
 B"1001", B"0001", B"1011", B"1100", 
 B"1101", B"0110", B"1101", B"0010", 
 B"1010", B"0001", B"0001", B"0111", 
 B"0001", B"1011", B"1100", B"1101", 
 B"0010", B"0001", B"0110", B"1101", 
 B"1111", B"0001", B"0011", B"0001", 
 B"1010", B"0100", B"0001", B"1111", 
 B"0011", B"1010", B"1011", B"1000", 
 B"1101", B"0011", B"0010", B"0001", 
 B"1110", B"0101", B"1111", B"0101", 
 B"1000", B"1001", B"0101", B"1011", 
 B"0111", B"1111", B"0001", B"0100", 
 B"1111", B"1000", B"1000", B"0111", 
 B"0101", B"0011", B"0001", B"0000", 
 B"0101", B"1101", B"1110", B"0001", 
 B"0110", B"1011", B"0110", B"0000", 
 B"1100", B"0001", B"1100", B"1101", 
 B"1111", B"0111", B"0001", B"0100", 
 B"0100", B"1100", B"1100", B"1101", 
 B"1010", B"1011", B"1010", B"1011", 
 B"1101", B"0100", B"0100", B"0011", 
 B"1111", B"1010", B"0110", B"1001", 
 B"1111", B"0110", B"0110", B"0000", 
 B"1010", B"0111", B"0111", B"0011", 
 B"0101", B"1001", B"0000", B"0111", 
 B"0110", B"1100", B"0001", B"1100", 
 B"1010", B"0101", B"0000", B"0010", 
 B"1111", B"0011", B"1001", B"1000", 
 B"0101", B"0110", B"1001", B"1110", 
 B"0111", B"1011", B"1000", B"0001", 
 B"1001", B"1110", B"1011", B"0101", 
 B"0001", B"1111", B"1111", B"0010", 
 B"1101", B"0010", B"0010", B"0001", 
 B"0100", B"0100", B"1101", B"1001", 
 B"1001", B"1100", B"1000", B"1001", 
 B"0010", B"0111", B"1010", B"0011", 
 B"0010", B"1011", B"0011", B"0110", 
 B"1010", B"0111", B"0010", B"0111", 
 B"0011", B"0011", B"0100", B"1110", 
 B"1110", B"1100", B"0001", B"0011", 
 B"0000", B"1010", B"1110", B"0010", 
 B"1001", B"1000", B"1100", B"1000", 
 B"0010", B"0001", B"0110", B"0100", 
 B"1011", B"1000", B"1111", B"1001", 
 B"0001", B"1101", B"0001", B"0000", 
 B"0101", B"0111", B"1001", B"1011", 
 B"1000", B"0111", B"1001", B"1000", 
 B"0011", B"1100", B"1000", B"1111", 
 B"1010", B"0111", B"0001", B"0101", 
 B"1001", B"1111", B"1101", B"1010", 
 B"0100", B"0010", B"0101", B"1010", 
 B"1011", B"0100", B"1000", B"0110", 
 B"1001", B"1100", B"1000", B"1100", 
 B"0011", B"1001", B"0011", B"1101", 
 B"1100", B"0000", B"1010", B"1000", 
 B"1001", B"0111", B"1001", B"1100", 
 B"0000", B"0101", B"0101", B"0010", 
 B"1011", B"0101", B"1100", B"0101", 
 B"1001", B"1010", B"1000", B"1100", 
 B"1000", B"1101", B"1101", B"0001", 
 B"0110", B"0110", B"1011", B"1010", 
 B"0010", B"1100", B"0111", B"0010", 
 B"0110", B"0001", B"0010", B"1111", 
 B"0110", B"0101", B"1111", B"0011", 
 B"1110", B"0000", B"1010", B"0110", 
 B"1101", B"0011", B"1010", B"0111", 
 B"0000", B"0110", B"0010", B"0001", 
 B"0100", B"1011", B"0011", B"0111", 
 B"0100", B"1010", B"0111", B"1110", 
 B"1100", B"1110", B"1101", B"0011", 
 B"0111", B"0010", B"0000", B"1111", 
 B"0010", B"1100", B"0110", B"0110", 
 B"0000", B"0000", B"1010", B"1101", 
 B"0100", B"0111", B"0001", B"1010", 
 B"0000", B"0011", B"1011", B"1010", 
 B"1100", B"1000", B"0101", B"1110", 
 B"1101", B"1001", B"1110", B"1111", 
 B"1110", B"0111", B"1101", B"1010", 
 B"1001", B"1010", B"1111", B"0111", 
 B"0110", B"1000", B"1010", B"0101", 
 B"1110", B"1010", B"0000", B"0111", 
 B"0110", B"1111", B"1000", B"1001", 
 B"0110", B"0101", B"0010", B"1011", 
 B"1111", B"0000", B"1100", B"0101", 
 B"0101", B"1101", B"0111", B"0111", 
 B"0101", B"0011", B"0101", B"0011", 
 B"0011", B"1000", B"1101", B"1011", 
 B"1000", B"0111", B"1010", B"1100", 
 B"1110", B"0100", B"0011", B"1110", 
 B"1001", B"1011", B"0100", B"1010", 
 B"1010", B"0101", B"1011", B"0101", 
 B"1011", B"0100", B"0110", B"0110", 
 B"1000", B"0010", B"1111", B"0010", 
 B"1111", B"1011", B"1000", B"0000", 
 B"0100", B"0110", B"0001", B"0010", 
 B"0001", B"0110", B"0100", B"1111", 
 B"0110", B"0001", B"0010", B"1001", 
 B"0011", B"0011", B"0100", B"0111", 
 B"0100", B"1111", B"0100", B"0101", 
 B"0100", B"1000", B"0011", B"1000", 
 B"0011", B"0110", B"1001", B"0101", 
 B"1001", B"1100", B"1011", B"0010", 
 B"0000", B"0010", B"0010", B"1110", 
 B"0100", B"0010", B"0100", B"0110", 
 B"1001", B"1101", B"1010", B"1111", 
 B"1101", B"0110", B"0100", B"0111", 
 B"0111", B"1000", B"0111", B"1000", 
 B"0010", B"0110", B"1000", B"1001", 
 B"0011", B"1100", B"0010", B"0010", 
 B"1111", B"0011", B"0000", B"1111", 
 B"1100", B"0001", B"1000", B"0001", 
 B"1000", B"0110", B"1010", B"1111", 
 B"0100", B"0111", B"0010", B"0111", 
 B"1001", B"0100", B"0001", B"1000", 
 B"0100", B"1110", B"0010", B"1110", 
 B"0110", B"1000", B"0110", B"0111", 
 B"0110", B"0001", B"0110", B"0001", 
 B"1101", B"1000", B"1111", B"1001", 
 B"0011", B"0011", B"1011", B"1111", 
 B"1100", B"1001", B"1101", B"1111", 
 B"0010", B"1101", B"0010", B"1010", 
 B"0100", B"1000", B"0000", B"0000", 
 B"1100", B"1011", B"0100", B"0011", 
 B"0100", B"1001", B"1001", B"0011", 
 B"1001", B"0110", B"1111", B"1011", 
 B"0001", B"1011", B"0000", B"0110", 
 B"0101", B"0111", B"0101", B"1101", 
 B"0011", B"0110", B"1100", B"1001", 
 B"1110", B"1111", B"1101", B"0110", 
 B"1010", B"0101", B"1000", B"1010", 
 B"0000", B"1011", B"1100", B"1000", 
 B"1111", B"0101", B"0111", B"1011", 
 B"0101", B"1101", B"1110", B"0101", 
 B"1000", B"0011", B"1101", B"1110", 
 B"0110", B"1100", B"1110", B"0000", 
 B"1011", B"1011", B"0000", B"0001", 
 B"0011", B"1101", B"0011", B"1111", 
 B"1000", B"1101", B"1001", B"1110", 
 B"1100", B"0100", B"0111", B"0010", 
 B"0010", B"1001", B"0111", B"1101", 
 B"0101", B"0100", B"0010", B"1000", 
 B"0000", B"1001", B"1011", B"0110", 
 B"1110", B"0100", B"0011", B"1100", 
 B"0001", B"0111", B"0000", B"1001", 
 B"1101", B"0000", B"1111", B"0011", 
 B"1000", B"1011", B"0001", B"0101", 
 B"0001", B"1110", B"1100", B"0101", 
 B"1110", B"0110", B"0011", B"0100", 
 B"0101", B"1111", B"0110", B"0101", 
 B"0011", B"1011", B"0100", B"1110", 
 B"0110", B"1100", B"1010", B"0111", 
 B"1111", B"1100", B"0011", B"1011", 
 B"1101", B"1101", B"1011", B"1011", 
 B"1100", B"0101", B"0001", B"1000", 
 B"1101", B"1100", B"1100", B"0001", 
 B"1101", B"1110", B"0101", B"0110", 
 B"0010", B"1000", B"1100", B"1101", 
 B"0101", B"1001", B"0110", B"1000", 
 B"1011", B"0100", B"0001", B"0100", 
 B"1111", B"1110", B"1000", B"1000", 
 B"0000", B"0001", B"1100", B"1100", 
 B"0101", B"1001", B"1001", B"1101", 
 B"0000", B"0010", B"1001", B"0001", 
 B"1001", B"0111", B"1111", B"1101", 
 B"0001", B"0010", B"0011", B"0010", 
 B"0001", B"0110", B"1111", B"0010", 
 B"0001", B"1000", B"1011", B"1010", 
 B"0100", B"1001", B"0100", B"1110", 
 B"1010", B"1000", B"1100", B"0010", 
 B"1100", B"0101", B"1100", B"1111", 
 B"0100", B"1011", B"0000", B"0101", 
 B"0111", B"0001", B"0110", B"0101", 
 B"0110", B"1011", B"1111", B"1101", 
 B"0111", B"1010", B"0110", B"0011", 
 B"0000", B"0001", B"0101", B"1001", 
 B"1001", B"1001", B"0001", B"1100", 
 B"1010", B"0110", B"0011", B"1111", 
 B"0010", B"1001", B"1110", B"1111", 
 B"0000", B"1011", B"0110", B"1001", 
 B"1101", B"0011", B"0010", B"1100", 
 B"1101", B"1000", B"0001", B"0011", 
 B"0101", B"0110", B"1001", B"0111", 
 B"1010", B"0010", B"1000", B"0100", 
 B"1111", B"0010", B"0000", B"0011", 
 B"1010", B"1010", B"1101", B"0111", 
 B"1011", B"0011", B"0100", B"1111", 
 B"1110", B"0111", B"0111", B"0010", 
 B"0011", B"0111", B"1100", B"0010", 
 B"0101", B"1010", B"0110", B"1111", 
 B"1101", B"0101", B"1100", B"1011", 
 B"1011", B"1011", B"1110", B"0100", 
 B"0111", B"0010", B"1100", B"1101", 
 B"1000", B"0000", B"0110", B"1011", 
 B"0011", B"0001", B"1111", B"0010", 
 B"1101", B"0001", B"0101", B"0111", 
 B"1000", B"1010", B"0000", B"1110", 
 B"1111", B"1111", B"1111", B"1011", 
 B"1110", B"1011", B"1111", B"0001", 
 B"1001", B"0101", B"0011", B"0001", 
 B"0110", B"1001", B"0010", B"0111", 
 B"1111", B"1101", B"1110", B"0110", 
 B"1010", B"1110", B"1100", B"1100", 
 B"1110", B"1111", B"0001", B"1010", 
 B"0111", B"0111", B"1011", B"1000", 
 B"1011", B"0000", B"0011", B"0100", 
 B"1001", B"0110", B"0010", B"1000", 
 B"0001", B"1101", B"1101", B"1010", 
 B"0001", B"1100", B"0000", B"1101", 
 B"0010", B"1111", B"1001", B"1000", 
 B"0100", B"1111", B"0111", B"1011", 
 B"0110", B"0000", B"0001", B"0010", 
 B"1101", B"0110", B"0110", B"0101", 
 B"1111", B"0011", B"1110", B"0101", 
 B"1010", B"1100", B"0101", B"1100", 
 B"0110", B"0010", B"0001", B"0000", 
 B"1101", B"1001", B"0001", B"0100", 
 B"1110", B"1000", B"0110", B"1100", 
 B"1000", B"1100", B"0111", B"1001", 
 B"1001", B"0110", B"1010", B"0001", 
 B"0110", B"0001", B"0101", B"1000", 
 B"0101", B"0101", B"0111", B"0000", 
 B"0111", B"1101", B"0010", B"0001", 
 B"0100", B"0011", B"1110", B"0100", 
 B"1110", B"1000", B"0110", B"1001", 
 B"1101", B"0100", B"0111", B"1000", 
 B"1011", B"0010", B"0111", B"0010", 
 B"1000", B"0110", B"0000", B"1000", 
 B"0101", B"1101", B"0010", B"1100", 
 B"1010", B"0000", B"1111", B"1001", 
 B"0000", B"1001", B"0101", B"0111", 
 B"1000", B"1100", B"0010", B"0001", 
 B"0010", B"1011", B"1000", B"0010", 
 B"0000", B"0100", B"0010", B"0001", 
 B"0100", B"1011", B"0001", B"1100", 
 B"1100", B"0110", B"1001", B"0100", 
 B"0101", B"1110", B"1010", B"0001", 
 B"0110", B"0100", B"1110", B"0111", 
 B"1111", B"1110", B"0001", B"1100", 
 B"0101", B"0000", B"1100", B"0011", 
 B"1001", B"0101", B"0101", B"1100", 
 B"0000", B"0100", B"1011", B"1011", 
 B"0001", B"1011", B"1001", B"1111", 
 B"0100", B"1001", B"0011", B"0000", 
 B"1010", B"1000", B"0110", B"1000", 
 B"0000", B"1101", B"0100", B"1100", 
 B"1110", B"0001", B"0111", B"0001", 
 B"0101", B"0001", B"0101", B"1000", 
 B"1111", B"1000", B"0111", B"1100", 
 B"0111", B"1010", B"0011", B"0010", 
 B"1101", B"0011", B"1011", B"0100", 
 B"1111", B"1101", B"1100", B"1000", 
 B"0100", B"1001", B"0011", B"1110", 
 B"0101", B"0101", B"1100", B"1111", 
 B"1100", B"1100", B"0001", B"1110", 
 B"1000", B"0101", B"1111", B"0101", 
 B"1011", B"1101", B"1001", B"1011", 
 B"1111", B"0001", B"0101", B"0001", 
 B"1000", B"1100", B"0110", B"1010", 
 B"1000", B"0011", B"1111", B"0011", 
 B"1100", B"1101", B"1101", B"1011", 
 B"0000", B"0011", B"1000", B"0001", 
 B"0011", B"1010", B"1000", B"0000", 
 B"0000", B"0111", B"1101", B"1100", 
 B"1110", B"1111", B"0010", B"0100", 
 B"1101", B"1000", B"1010", B"1011", 
 B"1001", B"0010", B"1111", B"1011", 
 B"0111", B"1010", B"1001", B"1110", 
 B"1110", B"0110", B"1101", B"1001", 
 B"0101", B"0101", B"1101", B"1001", 
 B"0101", B"0011", B"1001", B"0101", 
 B"0110", B"1111", B"1101", B"0100", 
 B"1111", B"1011", B"1001", B"1001", 
 B"0111", B"1010", B"0101", B"0010", 
 B"1000", B"1011", B"0100", B"0111", 
 B"0011", B"1101", B"1110", B"0001", 
 B"0101", B"0011", B"1000", B"1101", 
 B"0001", B"0000", B"0111", B"1010", 
 B"1000", B"0010", B"0000", B"0011", 
 B"0100", B"0100", B"0000", B"0111", 
 B"1000", B"0101", B"1001", B"1111", 
 B"1110", B"0010", B"0010", B"0000", 
 B"1100", B"0010", B"0111", B"0000", 
 B"1011", B"1110", B"1101", B"1110", 
 B"0000", B"0010", B"1001", B"0011", 
 B"1111", B"1100", B"0000", B"0101", 
 B"1101", B"0001", B"1110", B"0001", 
 B"1101", B"0000", B"0010", B"0110", 
 B"0000", B"0010", B"0011", B"0100", 
 B"1000", B"1011", B"0001", B"1101", 
 B"1110", B"1000", B"0001", B"0011", 
 B"0100", B"1001", B"0101", B"1001", 
 B"0010", B"1010", B"0001", B"0000", 
 B"1010", B"1110", B"0111", B"1101", 
 B"1111", B"1111", B"0100", B"1111", 
 B"1101", B"1110", B"0101", B"0111", 
 B"0011", B"1101", B"1100", B"1011", 
 B"1110", B"1110", B"0001", B"0101", 
 B"1110", B"1000", B"0111", B"0010", 
 B"0110", B"0111", B"1011", B"0100", 
 B"1110", B"0010", B"0001", B"1110", 
 B"0110", B"1010", B"0101", B"1000", 
 B"0110", B"1010", B"0101", B"1100", 
 B"0001", B"1001", B"1110", B"1000", 
 B"1000", B"1110", B"0101", B"0000", 
 B"1000", B"1101", B"1101", B"0101", 
 B"0001", B"1100", B"1101", B"1110", 
 B"0100", B"1101", B"0100", B"1011", 
 B"0010", B"1110", B"1100", B"0110", 
 B"1101", B"0001", B"0111", B"0001", 
 B"0100", B"0110", B"0100", B"0110", 
 B"1110", B"1011", B"1010", B"0100", 
 B"1011", B"0110", B"1010", B"0010", 
 B"1100", B"1110", B"0011", B"0010", 
 B"1100", B"0110", B"0011", B"1110", 
 B"1010", B"0111", B"0111", B"0010", 
 B"1101", B"1000", B"1111", B"1010", 
 B"1101", B"1001", B"1101", B"0110", 
 B"1010", B"0011", B"0010", B"1001", 
 B"0000", B"0101", B"0100", B"1010", 
 B"1110", B"1001", B"0110", B"1011", 
 B"1000", B"1101", B"1010", B"0010", 
 B"1111", B"1000", B"1011", B"0110", 
 B"1000", B"1010", B"0010", B"1100", 
 B"0000", B"1001", B"0110", B"1111", 
 B"1000", B"0100", B"1111", B"1101", 
 B"1011", B"0000", B"1010", B"0001", 
 B"0011", B"1011", B"1011", B"0010", 
 B"0110", B"1010", B"1000", B"1110", 
 B"0101", B"1010", B"1100", B"1010", 
 B"1110", B"1101", B"0001", B"0101", 
 B"0001", B"0110", B"1101", B"0111", 
 B"1100", B"1111", B"1111", B"0011", 
 B"0111", B"0000", B"0110", B"0100", 
 B"1001", B"1001", B"0100", B"0010", 
 B"1011", B"0010", B"1101", B"0000", 
 B"1110", B"0110", B"1111", B"1101", 
 B"0011", B"0111", B"1100", B"1110", 
 B"1011", B"1101", B"0001", B"1101", 
 B"0011", B"0010", B"1011", B"0011", 
 B"0001", B"1100", B"0001", B"1011", 
 B"0111", B"0101", B"1010", B"1010", 
 B"0001", B"0011", B"1110", B"0000", 
 B"1100", B"0111", B"0001", B"1000", 
 B"0010", B"0000", B"1111", B"0010", 
 B"1110", B"0111", B"1101", B"0011", 
 B"1101", B"1001", B"0001", B"0111", 
 B"1011", B"0101", B"0111", B"0010", 
 B"0100", B"0011", B"1011", B"1110", 
 B"1110", B"1111", B"1101", B"1110", 
 B"1001", B"1011", B"0100", B"0011", 
 B"1001", B"0011", B"1111", B"0100", 
 B"1000", B"1110", B"1001", B"1111", 
 B"1110", B"1100", B"1011", B"0111", 
 B"1001", B"0000", B"0100", B"1010", 
 B"0101", B"0010", B"1001", B"0110", 
 B"0111", B"1111", B"0111", B"0110", 
 B"1000", B"1101", B"0011", B"0111", 
 B"1101", B"1011", B"0000", B"0000", 
 B"1101", B"0100", B"1110", B"0110", 
 B"1010", B"0100", B"1111", B"1010", 
 B"1101", B"1101", B"0110", B"1100"

);

signal data_in          : bit_vector (3 downto 0);
signal reference_data   : bit_vector (3 downto 0);
signal senddata_counter : integer range 0 to 2499 := 2497;

begin

data_in        <= (y0 & y1 & y2 & y3);
senddata       <= senddata_tbl(senddata_counter);
reference_data <= senddata_tbl(senddata_counter);

process (start, clear)
begin
if (clear = '1') then
  senddata_counter <= 2497;
elsif (start = '0' and start'event) then
  if (senddata_counter < 2499) then
     senddata_counter <= senddata_counter + 1;
  else
     senddata_counter <= 0;
  end if;
end if;
end process;

match <= not(data_in xor reference_data);

end verify;
