--------------------------------------------------------------------------------
----                                                                        ----
---- This file is part of the yaVGA project                                 ----
---- http://www.opencores.org/?do=project&who=yavga                         ----
----                                                                        ----
---- Description                                                            ----
---- Implementation of yaVGA IP core                                        ----
----                                                                        ----
---- To Do:                                                                 ----
----                                                                        ----
----                                                                        ----
---- Author(s):                                                             ----
---- Sandro Amato, sdroamt@netscape.net                                     ----
----                                                                        ----
--------------------------------------------------------------------------------
----                                                                        ----
---- Copyright (c) 2009, Sandro Amato                                       ----
---- All rights reserved.                                                   ----
----                                                                        ----
---- Redistribution  and  use in  source  and binary forms, with or without ----
---- modification,  are  permitted  provided that  the following conditions ----
---- are met:                                                               ----
----                                                                        ----
----     * Redistributions  of  source  code  must  retain the above        ----
----       copyright   notice,  this  list  of  conditions  and  the        ----
----       following disclaimer.                                            ----
----     * Redistributions  in  binary form must reproduce the above        ----
----       copyright   notice,  this  list  of  conditions  and  the        ----
----       following  disclaimer in  the documentation and/or  other        ----
----       materials provided with the distribution.                        ----
----     * Neither  the  name  of  SANDRO AMATO nor the names of its        ----
----       contributors may be used to  endorse or  promote products        ----
----       derived from this software without specific prior written        ----
----       permission.                                                      ----
----                                                                        ----
---- THIS SOFTWARE IS PROVIDED  BY THE COPYRIGHT  HOLDERS AND  CONTRIBUTORS ----
---- "AS IS"  AND  ANY EXPRESS OR  IMPLIED  WARRANTIES, INCLUDING,  BUT NOT ----
---- LIMITED  TO, THE  IMPLIED  WARRANTIES  OF MERCHANTABILITY  AND FITNESS ----
---- FOR  A PARTICULAR  PURPOSE  ARE  DISCLAIMED. IN  NO  EVENT  SHALL  THE ----
---- COPYRIGHT  OWNER  OR CONTRIBUTORS  BE LIABLE FOR ANY DIRECT, INDIRECT, ----
---- INCIDENTAL,  SPECIAL,  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, ----
---- BUT  NOT LIMITED  TO,  PROCUREMENT OF  SUBSTITUTE  GOODS  OR SERVICES; ----
---- LOSS  OF  USE,  DATA,  OR PROFITS;  OR  BUSINESS INTERRUPTION) HOWEVER ----
---- CAUSED  AND  ON  ANY THEORY  OF LIABILITY, WHETHER IN CONTRACT, STRICT ----
---- LIABILITY,  OR  TORT  (INCLUDING  NEGLIGENCE  OR OTHERWISE) ARISING IN ----
---- ANY  WAY OUT  OF THE  USE  OF  THIS  SOFTWARE,  EVEN IF ADVISED OF THE ----
---- POSSIBILITY OF SUCH DAMAGE.                                            ----
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

use work.yavga_pkg.all;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity waveform_RAM is
  port (
    i_DIA    : in  std_logic_vector(c_WAVFRM_DATA_BUS_W - 1 downto 0);  -- 16-bit Data Input
    -- i_DIPA   : in std_logic;                       -- 2-bit parity Input
    -- i_ENA    : in std_logic;                       -- RAM Enable Input
    i_WEA    : in  std_logic;           -- Write Enable Input
    -- i_SSRA   : in std_logic;                       -- Synchronous Set/Reset Input
    i_clockA : in  std_logic;           -- Clock
    i_ADDRA  : in  std_logic_vector(c_WAVFRM_ADDR_BUS_W - 1 downto 0);  -- 10-bit Address Input
    --o_DOA     : out std_logic_vector(c_WAVFRM_DATA_BUS_W - 1 downto 0);  -- 16-bit Data Output
    -- o_DOPA   : out std_logic                       -- 2-bit parity Output
    --
    i_DIB    : in  std_logic_vector(c_WAVFRM_DATA_BUS_W - 1 downto 0);  -- 16-bit Data Input
    -- i_DIPB   : in std_logic;                       -- 2-bit parity Input
    -- i_ENB    : in std_logic;                       -- RAM Enable Input
    i_WEB    : in  std_logic;           -- Write Enable Input
    -- i_SSRB   : in std_logic;                       -- Synchronous Set/Reset Input
    i_clockB : in  std_logic;           -- Clock
    i_ADDRB  : in  std_logic_vector(c_WAVFRM_ADDR_BUS_W - 1 downto 0);  -- 10-bit Address Input
    o_DOB    : out std_logic_vector(c_WAVFRM_DATA_BUS_W - 1 downto 0)  -- 16-bit Data Output
    -- o_DOPB   : out std_logic                       -- 2-bit parity Output
    );
end waveform_RAM;

architecture Behavioral of waveform_RAM is

  constant c_ram_size : natural := 2**(c_WAVFRM_ADDR_BUS_W);

  type t_ram is array (c_ram_size-1 downto 0) of
    std_logic_vector (c_WAVFRM_DATA_BUS_W - 1 downto 0);

  shared variable v_ram : t_ram := (
    0      => X"1000" or X"00BF",
    1      => X"1000" or X"00BE",
    2      => X"1000" or X"00BD",
    3      => X"1000" or X"00BD",
    4      => X"1000" or X"00BC",
    5      => X"1000" or X"00BB",
    6      => X"1000" or X"00BB",
    7      => X"1000" or X"00BA",
    8      => X"1000" or X"00B9",
    9      => X"1000" or X"00B9",
    10     => X"1000" or X"00B8",
    11     => X"1000" or X"00B7",
    12     => X"1000" or X"00B7",
    13     => X"1000" or X"00B6",
    14     => X"1000" or X"00B5",
    15     => X"1000" or X"00B5",
    16     => X"1000" or X"00B4",
    17     => X"1000" or X"00B3",
    18     => X"1000" or X"00B3",
    19     => X"1000" or X"00B2",
    20     => X"1000" or X"00B1",
    21     => X"1000" or X"00B1",
    22     => X"1000" or X"00B0",
    23     => X"1000" or X"00B0",
    24     => X"1000" or X"00AF",
    25     => X"1000" or X"00AE",
    26     => X"1000" or X"00AE",
    27     => X"1000" or X"00AD",
    28     => X"1000" or X"00AD",
    29     => X"1000" or X"00AC",
    30     => X"1000" or X"00AB",
    31     => X"1000" or X"00AB",
    32     => X"1000" or X"00AA",
    33     => X"1000" or X"00AA",
    34     => X"1000" or X"00A9",
    35     => X"1000" or X"00A9",
    36     => X"1000" or X"00A8",
    37     => X"1000" or X"00A8",
    38     => X"1000" or X"00A7",
    39     => X"1000" or X"00A7",
    40     => X"1000" or X"00A6",
    41     => X"1000" or X"00A6",
    42     => X"1000" or X"00A5",
    43     => X"1000" or X"00A5",
    44     => X"1000" or X"00A4",
    45     => X"1000" or X"00A4",
    46     => X"1000" or X"00A3",
    47     => X"1000" or X"00A3",
    48     => X"1000" or X"00A2",
    49     => X"1000" or X"00A2",
    50     => X"1000" or X"00A2",
    51     => X"1000" or X"00A1",
    52     => X"1000" or X"00A1",
    53     => X"1000" or X"00A1",
    54     => X"1000" or X"00A0",
    55     => X"1000" or X"00A0",
    56     => X"1000" or X"00A0",
    57     => X"1000" or X"009F",
    58     => X"1000" or X"009F",
    59     => X"1000" or X"009F",
    60     => X"1000" or X"009E",
    61     => X"1000" or X"009E",
    62     => X"1000" or X"009E",
    63     => X"1000" or X"009E",
    64     => X"1000" or X"009E",
    65     => X"1000" or X"009D",
    66     => X"1000" or X"009D",
    67     => X"1000" or X"009D",
    68     => X"1000" or X"009D",
    69     => X"1000" or X"009D",
    70     => X"1000" or X"009D",
    71     => X"1000" or X"009D",
    72     => X"1000" or X"009D",
    73     => X"1000" or X"009D",
    74     => X"1000" or X"009D",
    75     => X"1000" or X"009D",
    76     => X"1000" or X"009D",
    77     => X"1000" or X"009D",
    78     => X"1000" or X"009D",
    79     => X"1000" or X"009D",
    80     => X"1000" or X"009D",
    81     => X"1000" or X"009D",
    82     => X"1000" or X"009D",
    83     => X"1000" or X"009D",
    84     => X"1000" or X"009D",
    85     => X"1000" or X"009D",
    86     => X"1000" or X"009E",
    87     => X"1000" or X"009E",
    88     => X"1000" or X"009E",
    89     => X"1000" or X"009E",
    90     => X"1000" or X"009E",
    91     => X"1000" or X"009F",
    92     => X"1000" or X"009F",
    93     => X"1000" or X"009F",
    94     => X"1000" or X"00A0",
    95     => X"1000" or X"00A0",
    96     => X"1000" or X"00A0",
    97     => X"1000" or X"00A1",
    98     => X"1000" or X"00A1",
    99     => X"1000" or X"00A2",
    100    => X"1000" or X"00A2",
    101    => X"1000" or X"00A3",
    102    => X"1000" or X"00A3",
    103    => X"1000" or X"00A4",
    104    => X"1000" or X"00A4",
    105    => X"1000" or X"00A5",
    106    => X"1000" or X"00A5",
    107    => X"1000" or X"00A6",
    108    => X"1000" or X"00A7",
    109    => X"1000" or X"00A7",
    110    => X"1000" or X"00A8",
    111    => X"1000" or X"00A8",
    112    => X"1000" or X"00A9",
    113    => X"1000" or X"00AA",
    114    => X"1000" or X"00AB",
    115    => X"1000" or X"00AB",
    116    => X"1000" or X"00AC",
    117    => X"1000" or X"00AD",
    118    => X"1000" or X"00AE",
    119    => X"1000" or X"00AF",
    120    => X"1000" or X"00AF",
    121    => X"1000" or X"00B0",
    122    => X"1000" or X"00B1",
    123    => X"1000" or X"00B2",
    124    => X"1000" or X"00B3",
    125    => X"1000" or X"00B4",
    126    => X"1000" or X"00B5",
    127    => X"1000" or X"00B6",
    128    => X"1000" or X"00B7",
    129    => X"1000" or X"00B8",
    130    => X"1000" or X"00B9",
    131    => X"1000" or X"00BA",
    132    => X"1000" or X"00BB",
    133    => X"1000" or X"00BC",
    134    => X"1000" or X"00BD",
    135    => X"1000" or X"00BE",
    136    => X"1000" or X"00C0",
    137    => X"1000" or X"00C1",
    138    => X"1000" or X"00C2",
    139    => X"1000" or X"00C3",
    140    => X"1000" or X"00C4",
    141    => X"1000" or X"00C6",
    142    => X"1000" or X"00C7",
    143    => X"1000" or X"00C8",
    144    => X"1000" or X"00C9",
    145    => X"1000" or X"00CB",
    146    => X"1000" or X"00CC",
    147    => X"1000" or X"00CD",
    148    => X"1000" or X"00CF",
    149    => X"1000" or X"00D0",
    150    => X"1000" or X"00D1",
    151    => X"1000" or X"00D3",
    152    => X"1000" or X"00D4",
    153    => X"1000" or X"00D6",
    154    => X"1000" or X"00D7",
    155    => X"1000" or X"00D8",
    156    => X"1000" or X"00DA",
    157    => X"1000" or X"00DB",
    158    => X"1000" or X"00DD",
    159    => X"1000" or X"00DE",
    160    => X"1000" or X"00E0",
    161    => X"1000" or X"00E1",
    162    => X"1000" or X"00E3",
    163    => X"1000" or X"00E5",
    164    => X"1000" or X"00E6",
    165    => X"1000" or X"00E8",
    166    => X"1000" or X"00E9",
    167    => X"1000" or X"00EB",
    168    => X"1000" or X"00EC",
    169    => X"1000" or X"00EE",
    170    => X"1000" or X"00F0",
    171    => X"1000" or X"00F1",
    172    => X"1000" or X"00F3",
    173    => X"1000" or X"00F5",
    174    => X"1000" or X"00F6",
    175    => X"1000" or X"00F8",
    176    => X"1000" or X"00FA",
    177    => X"1000" or X"00FB",
    178    => X"1000" or X"00FD",
    179    => X"1000" or X"00FF",
    180    => X"1000" or X"0100",
    181    => X"1000" or X"0102",
    182    => X"1000" or X"0104",
    183    => X"1000" or X"0105",
    184    => X"1000" or X"0107",
    185    => X"1000" or X"0109",
    186    => X"1000" or X"010B",
    187    => X"1000" or X"010C",
    188    => X"1000" or X"010E",
    189    => X"1000" or X"0110",
    190    => X"1000" or X"0111",
    191    => X"1000" or X"0113",
    192    => X"1000" or X"0115",
    193    => X"1000" or X"0117",
    194    => X"1000" or X"0118",
    195    => X"1000" or X"011A",
    196    => X"1000" or X"011C",
    197    => X"1000" or X"011E",
    198    => X"1000" or X"011F",
    199    => X"1000" or X"0121",
    200    => X"1000" or X"0123",
    201    => X"1000" or X"0125",
    202    => X"1000" or X"0126",
    203    => X"1000" or X"0128",
    204    => X"1000" or X"012A",
    205    => X"1000" or X"012C",
    206    => X"1000" or X"012D",
    207    => X"1000" or X"012F",
    208    => X"1000" or X"0131",
    209    => X"1000" or X"0132",
    210    => X"1000" or X"0134",
    211    => X"1000" or X"0136",
    212    => X"1000" or X"0138",
    213    => X"1000" or X"0139",
    214    => X"1000" or X"013B",
    215    => X"1000" or X"013D",
    216    => X"1000" or X"013E",
    217    => X"1000" or X"0140",
    218    => X"1000" or X"0142",
    219    => X"1000" or X"0143",
    220    => X"1000" or X"0145",
    221    => X"1000" or X"0147",
    222    => X"1000" or X"0148",
    223    => X"1000" or X"014A",
    224    => X"1000" or X"014B",
    225    => X"1000" or X"014D",
    226    => X"1000" or X"014F",
    227    => X"1000" or X"0150",
    228    => X"1000" or X"0152",
    229    => X"1000" or X"0153",
    230    => X"1000" or X"0155",
    231    => X"1000" or X"0156",
    232    => X"1000" or X"0158",
    233    => X"1000" or X"0159",
    234    => X"1000" or X"015B",
    235    => X"1000" or X"015C",
    236    => X"1000" or X"015E",
    237    => X"1000" or X"015F",
    238    => X"1000" or X"0161",
    239    => X"1000" or X"0162",
    240    => X"1000" or X"0163",
    241    => X"1000" or X"0165",
    242    => X"1000" or X"0166",
    243    => X"1000" or X"0167",
    244    => X"1000" or X"0169",
    245    => X"1000" or X"016A",
    246    => X"1000" or X"016B",
    247    => X"1000" or X"016D",
    248    => X"1000" or X"016E",
    249    => X"1000" or X"016F",
    250    => X"1000" or X"0170",
    251    => X"1000" or X"0171",
    252    => X"1000" or X"0173",
    253    => X"1000" or X"0174",
    254    => X"1000" or X"0175",
    255    => X"1000" or X"0176",
    256    => X"1000" or X"0177",
    257    => X"1000" or X"0178",
    258    => X"1000" or X"0179",
    259    => X"1000" or X"017A",
    260    => X"1000" or X"017B",
    261    => X"1000" or X"017C",
    262    => X"1000" or X"017D",
    263    => X"1000" or X"017E",
    264    => X"1000" or X"017F",
    265    => X"1000" or X"0180",
    266    => X"1000" or X"0181",
    267    => X"1000" or X"0182",
    268    => X"1000" or X"0183",
    269    => X"1000" or X"0183",
    270    => X"1000" or X"0184",
    271    => X"1000" or X"0185",
    272    => X"1000" or X"0186",
    273    => X"1000" or X"0186",
    274    => X"1000" or X"0187",
    275    => X"1000" or X"0188",
    276    => X"1000" or X"0188",
    277    => X"1000" or X"0189",
    278    => X"1000" or X"018A",
    279    => X"1000" or X"018A",
    280    => X"1000" or X"018B",
    281    => X"1000" or X"018B",
    282    => X"1000" or X"018C",
    283    => X"1000" or X"018C",
    284    => X"1000" or X"018D",
    285    => X"1000" or X"018D",
    286    => X"1000" or X"018D",
    287    => X"1000" or X"018E",
    288    => X"1000" or X"018E",
    289    => X"1000" or X"018E",
    290    => X"1000" or X"018F",
    291    => X"1000" or X"018F",
    292    => X"1000" or X"018F",
    293    => X"1000" or X"018F",
    294    => X"1000" or X"0190",
    295    => X"1000" or X"0190",
    296    => X"1000" or X"0190",
    297    => X"1000" or X"0190",
    298    => X"1000" or X"0190",
    299    => X"1000" or X"0190",
    300    => X"1000" or X"0190",
    301    => X"1000" or X"0190",
    302    => X"1000" or X"0190",
    303    => X"1000" or X"0190",
    304    => X"1000" or X"0190",
    305    => X"1000" or X"0190",
    306    => X"1000" or X"0190",
    307    => X"1000" or X"018F",
    308    => X"1000" or X"018F",
    309    => X"1000" or X"018F",
    310    => X"1000" or X"018F",
    311    => X"1000" or X"018E",
    312    => X"1000" or X"018E",
    313    => X"1000" or X"018E",
    314    => X"1000" or X"018D",
    315    => X"1000" or X"018D",
    316    => X"1000" or X"018D",
    317    => X"1000" or X"018C",
    318    => X"1000" or X"018C",
    319    => X"1000" or X"018B",
    320    => X"1000" or X"018B",
    321    => X"1000" or X"018A",
    322    => X"1000" or X"018A",
    323    => X"1000" or X"0189",
    324    => X"1000" or X"0188",
    325    => X"1000" or X"0188",
    326    => X"1000" or X"0187",
    327    => X"1000" or X"0186",
    328    => X"1000" or X"0186",
    329    => X"1000" or X"0185",
    330    => X"1000" or X"0184",
    331    => X"1000" or X"0183",
    332    => X"1000" or X"0183",
    333    => X"1000" or X"0182",
    334    => X"1000" or X"0181",
    335    => X"1000" or X"0180",
    336    => X"1000" or X"017F",
    337    => X"1000" or X"017E",
    338    => X"1000" or X"017D",
    339    => X"1000" or X"017C",
    340    => X"1000" or X"017B",
    341    => X"1000" or X"017A",
    342    => X"1000" or X"0179",
    343    => X"1000" or X"0178",
    344    => X"1000" or X"0177",
    345    => X"1000" or X"0176",
    346    => X"1000" or X"0175",
    347    => X"1000" or X"0174",
    348    => X"1000" or X"0173",
    349    => X"1000" or X"0171",
    350    => X"1000" or X"0170",
    351    => X"1000" or X"016F",
    352    => X"1000" or X"016E",
    353    => X"1000" or X"016D",
    354    => X"1000" or X"016B",
    355    => X"1000" or X"016A",
    356    => X"1000" or X"0169",
    357    => X"1000" or X"0167",
    358    => X"1000" or X"0166",
    359    => X"1000" or X"0165",
    360    => X"1000" or X"0163",
    361    => X"1000" or X"0162",
    362    => X"1000" or X"0161",
    363    => X"1000" or X"015F",
    364    => X"1000" or X"015E",
    365    => X"1000" or X"015C",
    366    => X"1000" or X"015B",
    367    => X"1000" or X"0159",
    368    => X"1000" or X"0158",
    369    => X"1000" or X"0156",
    370    => X"1000" or X"0155",
    371    => X"1000" or X"0153",
    372    => X"1000" or X"0152",
    373    => X"1000" or X"0150",
    374    => X"1000" or X"014F",
    375    => X"1000" or X"014D",
    376    => X"1000" or X"014B",
    377    => X"1000" or X"014A",
    378    => X"1000" or X"0148",
    379    => X"1000" or X"0147",
    380    => X"1000" or X"0145",
    381    => X"1000" or X"0143",
    382    => X"1000" or X"0142",
    383    => X"1000" or X"0140",
    384    => X"1000" or X"013E",
    385    => X"1000" or X"013D",
    386    => X"1000" or X"013B",
    387    => X"1000" or X"0139",
    388    => X"1000" or X"0138",
    389    => X"1000" or X"0136",
    390    => X"1000" or X"0134",
    391    => X"1000" or X"0132",
    392    => X"1000" or X"0131",
    393    => X"1000" or X"012F",
    394    => X"1000" or X"012D",
    395    => X"1000" or X"012C",
    396    => X"1000" or X"012A",
    397    => X"1000" or X"0128",
    398    => X"1000" or X"0126",
    399    => X"1000" or X"0125",
    400    => X"1000" or X"0123",
    401    => X"1000" or X"0121",
    402    => X"1000" or X"011F",
    403    => X"1000" or X"011E",
    404    => X"1000" or X"011C",
    405    => X"1000" or X"011A",
    406    => X"1000" or X"0118",
    407    => X"1000" or X"0117",
    408    => X"1000" or X"0115",
    409    => X"1000" or X"0113",
    410    => X"1000" or X"0111",
    411    => X"1000" or X"0110",
    412    => X"1000" or X"010E",
    413    => X"1000" or X"010C",
    414    => X"1000" or X"010B",
    415    => X"1000" or X"0109",
    416    => X"1000" or X"0107",
    417    => X"1000" or X"0105",
    418    => X"1000" or X"0104",
    419    => X"1000" or X"0102",
    420    => X"1000" or X"0100",
    421    => X"1000" or X"00FF",
    422    => X"1000" or X"00FD",
    423    => X"1000" or X"00FB",
    424    => X"1000" or X"00FA",
    425    => X"1000" or X"00F8",
    426    => X"1000" or X"00F6",
    427    => X"1000" or X"00F5",
    428    => X"1000" or X"00F3",
    429    => X"1000" or X"00F1",
    430    => X"1000" or X"00F0",
    431    => X"1000" or X"00EE",
    432    => X"1000" or X"00EC",
    433    => X"1000" or X"00EB",
    434    => X"1000" or X"00E9",
    435    => X"1000" or X"00E8",
    436    => X"1000" or X"00E6",
    437    => X"1000" or X"00E5",
    438    => X"1000" or X"00E3",
    439    => X"1000" or X"00E1",
    440    => X"1000" or X"00E0",
    441    => X"1000" or X"00DE",
    442    => X"1000" or X"00DD",
    443    => X"1000" or X"00DB",
    444    => X"1000" or X"00DA",
    445    => X"1000" or X"00D8",
    446    => X"1000" or X"00D7",
    447    => X"1000" or X"00D6",
    448    => X"1000" or X"00D4",
    449    => X"1000" or X"00D3",
    450    => X"1000" or X"00D1",
    451    => X"1000" or X"00D0",
    452    => X"1000" or X"00CF",
    453    => X"1000" or X"00CD",
    454    => X"1000" or X"00CC",
    455    => X"1000" or X"00CB",
    456    => X"1000" or X"00C9",
    457    => X"1000" or X"00C8",
    458    => X"1000" or X"00C7",
    459    => X"1000" or X"00C6",
    460    => X"1000" or X"00C4",
    461    => X"1000" or X"00C3",
    462    => X"1000" or X"00C2",
    463    => X"1000" or X"00C1",
    464    => X"1000" or X"00C0",
    465    => X"1000" or X"00BE",
    466    => X"1000" or X"00BD",
    467    => X"1000" or X"00BC",
    468    => X"1000" or X"00BB",
    469    => X"1000" or X"00BA",
    470    => X"1000" or X"00B9",
    471    => X"1000" or X"00B8",
    472    => X"1000" or X"00B7",
    473    => X"1000" or X"00B6",
    474    => X"1000" or X"00B5",
    475    => X"1000" or X"00B4",
    476    => X"1000" or X"00B3",
    477    => X"1000" or X"00B2",
    478    => X"1000" or X"00B1",
    479    => X"1000" or X"00B0",
    480    => X"1000" or X"00AF",
    481    => X"1000" or X"00AF",
    482    => X"1000" or X"00AE",
    483    => X"1000" or X"00AD",
    484    => X"1000" or X"00AC",
    485    => X"1000" or X"00AB",
    486    => X"1000" or X"00AB",
    487    => X"1000" or X"00AA",
    488    => X"1000" or X"00A9",
    489    => X"1000" or X"00A8",
    490    => X"1000" or X"00A8",
    491    => X"1000" or X"00A7",
    492    => X"1000" or X"00A7",
    493    => X"1000" or X"00A6",
    494    => X"1000" or X"00A5",
    495    => X"1000" or X"00A5",
    496    => X"1000" or X"00A4",
    497    => X"1000" or X"00A4",
    498    => X"1000" or X"00A3",
    499    => X"1000" or X"00A3",
    500    => X"1000" or X"00A2",
    501    => X"1000" or X"00A2",
    502    => X"1000" or X"00A1",
    503    => X"1000" or X"00A1",
    504    => X"1000" or X"00A0",
    505    => X"1000" or X"00A0",
    506    => X"1000" or X"00A0",
    507    => X"1000" or X"009F",
    508    => X"1000" or X"009F",
    509    => X"1000" or X"009F",
    510    => X"1000" or X"009E",
    511    => X"1000" or X"009E",
    512    => X"1000" or X"009E",
    513    => X"1000" or X"009E",
    514    => X"1000" or X"009E",
    515    => X"1000" or X"009D",
    516    => X"1000" or X"009D",
    517    => X"1000" or X"009D",
    518    => X"1000" or X"009D",
    519    => X"1000" or X"009D",
    520    => X"1000" or X"009D",
    521    => X"1000" or X"009D",
    522    => X"1000" or X"009D",
    523    => X"1000" or X"009D",
    524    => X"1000" or X"009D",
    525    => X"1000" or X"009D",
    526    => X"1000" or X"009D",
    527    => X"1000" or X"009D",
    528    => X"1000" or X"009D",
    529    => X"1000" or X"009D",
    530    => X"1000" or X"009D",
    531    => X"1000" or X"009D",
    532    => X"1000" or X"009D",
    533    => X"1000" or X"009D",
    534    => X"1000" or X"009D",
    535    => X"1000" or X"009D",
    536    => X"1000" or X"009E",
    537    => X"1000" or X"009E",
    538    => X"1000" or X"009E",
    539    => X"1000" or X"009E",
    540    => X"1000" or X"009E",
    541    => X"1000" or X"009F",
    542    => X"1000" or X"009F",
    543    => X"1000" or X"009F",
    544    => X"1000" or X"00A0",
    545    => X"1000" or X"00A0",
    546    => X"1000" or X"00A0",
    547    => X"1000" or X"00A1",
    548    => X"1000" or X"00A1",
    549    => X"1000" or X"00A1",
    550    => X"1000" or X"00A2",
    551    => X"1000" or X"00A2",
    552    => X"1000" or X"00A2",
    553    => X"1000" or X"00A3",
    554    => X"1000" or X"00A3",
    555    => X"1000" or X"00A4",
    556    => X"1000" or X"00A4",
    557    => X"1000" or X"00A5",
    558    => X"1000" or X"00A5",
    559    => X"1000" or X"00A6",
    560    => X"1000" or X"00A6",
    561    => X"1000" or X"00A7",
    562    => X"1000" or X"00A7",
    563    => X"1000" or X"00A8",
    564    => X"1000" or X"00A8",
    565    => X"1000" or X"00A9",
    566    => X"1000" or X"00A9",
    567    => X"1000" or X"00AA",
    568    => X"1000" or X"00AA",
    569    => X"1000" or X"00AB",
    570    => X"1000" or X"00AB",
    571    => X"1000" or X"00AC",
    572    => X"1000" or X"00AD",
    573    => X"1000" or X"00AD",
    574    => X"1000" or X"00AE",
    575    => X"1000" or X"00AE",
    576    => X"1000" or X"00AF",
    577    => X"1000" or X"00B0",
    578    => X"1000" or X"00B0",
    579    => X"1000" or X"00B1",
    580    => X"1000" or X"00B1",
    581    => X"1000" or X"00B2",
    582    => X"1000" or X"00B3",
    583    => X"1000" or X"00B3",
    584    => X"1000" or X"00B4",
    585    => X"1000" or X"00B5",
    586    => X"1000" or X"00B5",
    587    => X"1000" or X"00B6",
    588    => X"1000" or X"00B7",
    589    => X"1000" or X"00B7",
    590    => X"1000" or X"00B8",
    591    => X"1000" or X"00B9",
    592    => X"1000" or X"00B9",
    593    => X"1000" or X"00BA",
    594    => X"1000" or X"00BB",
    595    => X"1000" or X"00BB",
    596    => X"1000" or X"00BC",
    597    => X"1000" or X"00BD",
    598    => X"1000" or X"00BD",
    599    => X"1000" or X"00BE",
    600    => X"1000" or X"00BF",
    601    => X"1000" or X"00BF",
    602    => X"1000" or X"00C0",
    603    => X"1000" or X"00C1",
    604    => X"1000" or X"00C1",
    605    => X"1000" or X"00C2",
    606    => X"1000" or X"00C3",
    607    => X"1000" or X"00C3",
    608    => X"1000" or X"00C4",
    609    => X"1000" or X"00C5",
    610    => X"1000" or X"00C5",
    611    => X"1000" or X"00C6",
    612    => X"1000" or X"00C7",
    613    => X"1000" or X"00C7",
    614    => X"1000" or X"00C8",
    615    => X"1000" or X"00C9",
    616    => X"1000" or X"00C9",
    617    => X"1000" or X"00CA",
    618    => X"1000" or X"00CA",
    619    => X"1000" or X"00CB",
    620    => X"1000" or X"00CC",
    621    => X"1000" or X"00CC",
    622    => X"1000" or X"00CD",
    623    => X"1000" or X"00CD",
    624    => X"1000" or X"00CE",
    625    => X"1000" or X"00CF",
    626    => X"1000" or X"00CF",
    627    => X"1000" or X"00D0",
    628    => X"1000" or X"00D0",
    629    => X"1000" or X"00D1",
    630    => X"1000" or X"00D1",
    631    => X"1000" or X"00D2",
    632    => X"1000" or X"00D3",
    633    => X"1000" or X"00D3",
    634    => X"1000" or X"00D4",
    635    => X"1000" or X"00D4",
    636    => X"1000" or X"00D5",
    637    => X"1000" or X"00D5",
    638    => X"1000" or X"00D6",
    639    => X"1000" or X"00D6",
    640    => X"1000" or X"00D7",
    641    => X"1000" or X"00D7",
    642    => X"1000" or X"00D7",
    643    => X"1000" or X"00D8",
    644    => X"1000" or X"00D8",
    645    => X"1000" or X"00D9",
    646    => X"1000" or X"00D9",
    647    => X"1000" or X"00DA",
    648    => X"1000" or X"00DA",
    649    => X"1000" or X"00DA",
    650    => X"1000" or X"00DB",
    651    => X"1000" or X"00DB",
    652    => X"1000" or X"00DC",
    653    => X"1000" or X"00DC",
    654    => X"1000" or X"00DC",
    655    => X"1000" or X"00DD",
    656    => X"1000" or X"00DD",
    657    => X"1000" or X"00DD",
    658    => X"1000" or X"00DD",
    659    => X"1000" or X"00DE",
    660    => X"1000" or X"00DE",
    661    => X"1000" or X"00DE",
    662    => X"1000" or X"00DF",
    663    => X"1000" or X"00DF",
    664    => X"1000" or X"00DF",
    665    => X"1000" or X"00DF",
    666    => X"1000" or X"00E0",
    667    => X"1000" or X"00E0",
    668    => X"1000" or X"00E0",
    669    => X"1000" or X"00E0",
    670    => X"1000" or X"00E0",
    671    => X"1000" or X"00E0",
    672    => X"1000" or X"00E1",
    673    => X"1000" or X"00E1",
    674    => X"1000" or X"00E1",
    675    => X"1000" or X"00E1",
    676    => X"1000" or X"00E1",
    677    => X"1000" or X"00E1",
    678    => X"1000" or X"00E1",
    679    => X"1000" or X"00E1",
    680    => X"1000" or X"00E1",
    681    => X"1000" or X"00E2",
    682    => X"1000" or X"00E2",
    683    => X"1000" or X"00E2",
    684    => X"1000" or X"00E2",
    685    => X"1000" or X"00E2",
    686    => X"1000" or X"00E2",
    687    => X"1000" or X"00E2",
    688    => X"1000" or X"00E2",
    689    => X"1000" or X"00E2",
    690    => X"1000" or X"00E2",
    691    => X"1000" or X"00E2",
    692    => X"1000" or X"00E2",
    693    => X"1000" or X"00E1",
    694    => X"1000" or X"00E1",
    695    => X"1000" or X"00E1",
    696    => X"1000" or X"00E1",
    697    => X"1000" or X"00E1",
    698    => X"1000" or X"00E1",
    699    => X"1000" or X"00E1",
    700    => X"1000" or X"00E1",
    701    => X"1000" or X"00E1",
    702    => X"1000" or X"00E0",
    703    => X"1000" or X"00E0",
    704    => X"1000" or X"00E0",
    705    => X"1000" or X"00E0",
    706    => X"1000" or X"00E0",
    707    => X"1000" or X"00E0",
    708    => X"1000" or X"00DF",
    709    => X"1000" or X"00DF",
    710    => X"1000" or X"00DF",
    711    => X"1000" or X"00DF",
    712    => X"1000" or X"00DE",
    713    => X"1000" or X"00DE",
    714    => X"1000" or X"00DE",
    715    => X"1000" or X"00DE",
    716    => X"1000" or X"00DD",
    717    => X"1000" or X"00DD",
    718    => X"1000" or X"00DD",
    719    => X"1000" or X"00DD",
    720    => X"1000" or X"00DC",
    721    => X"1000" or X"00DC",
    722    => X"1000" or X"00DC",
    723    => X"1000" or X"00DB",
    724    => X"1000" or X"00DB",
    725    => X"1000" or X"00DB",
    726    => X"1000" or X"00DA",
    727    => X"1000" or X"00DA",
    728    => X"1000" or X"00DA",
    729    => X"1000" or X"00D9",
    730    => X"1000" or X"00D9",
    731    => X"1000" or X"00D9",
    732    => X"1000" or X"00D8",
    733    => X"1000" or X"00D8",
    734    => X"1000" or X"00D8",
    735    => X"1000" or X"00D7",
    736    => X"1000" or X"00D7",
    737    => X"1000" or X"00D6",
    738    => X"1000" or X"00D6",
    739    => X"1000" or X"00D6",
    740    => X"1000" or X"00D5",
    741    => X"1000" or X"00D5",
    742    => X"1000" or X"00D4",
    743    => X"1000" or X"00D4",
    744    => X"1000" or X"00D4",
    745    => X"1000" or X"00D3",
    746    => X"1000" or X"00D3",
    747    => X"1000" or X"00D2",
    748    => X"1000" or X"00D2",
    749    => X"1000" or X"00D2",
    750    => X"1000" or X"00D1",
    751    => X"1000" or X"00D1",
    752    => X"1000" or X"00D0",
    753    => X"1000" or X"00D0",
    754    => X"1000" or X"00CF",
    755    => X"1000" or X"00CF",
    756    => X"1000" or X"00CF",
    757    => X"1000" or X"00CE",
    758    => X"1000" or X"00CE",
    759    => X"1000" or X"00CD",
    760    => X"1000" or X"00CD",
    761    => X"1000" or X"00CC",
    762    => X"1000" or X"00CC",
    763    => X"1000" or X"00CC",
    764    => X"1000" or X"00CB",
    765    => X"1000" or X"00CB",
    766    => X"1000" or X"00CA",
    767    => X"1000" or X"00CA",
    768    => X"1000" or X"00C9",
    769    => X"1000" or X"00C9",
    770    => X"1000" or X"00C9",
    771    => X"1000" or X"00C8",
    772    => X"1000" or X"00C8",
    773    => X"1000" or X"00C7",
    774    => X"1000" or X"00C7",
    775    => X"1000" or X"00C6",
    776    => X"1000" or X"00C6",
    777    => X"1000" or X"00C6",
    778    => X"1000" or X"00C5",
    779    => X"1000" or X"00C5",
    780    => X"1000" or X"00C4",
    781    => X"1000" or X"00C4",
    782    => X"1000" or X"00C4",
    783    => X"1000" or X"00C3",
    784    => X"1000" or X"00C3",
    785    => X"1000" or X"00C2",
    786    => X"1000" or X"00C2",
    787    => X"1000" or X"00C2",
    788    => X"1000" or X"00C1",
    789    => X"1000" or X"00C1",
    790    => X"1000" or X"00C1",
    791    => X"1000" or X"00C0",
    792    => X"1000" or X"00C0",
    793    => X"1000" or X"00BF",
    794    => X"1000" or X"00BF",
    795    => X"1000" or X"00BF",
    796    => X"1000" or X"00BE",
    797    => X"1000" or X"00BE",
    798    => X"1000" or X"00BE",
    799    => X"1000" or X"00BD",
    800    => X"1000" or X"00BD",
    others => X"1000" or X"0064"
    );

begin
  -- wave form or video-line memory
  -- |------| |-------------------------------------------|
  -- | P  P | |  D  D  D |  D  D  D | D D D D D D D D D D |
  -- |======| |===========================================|
  -- |17 16 | | 15 14 13 | 12 11 10 | 9 8 7 6 5 4 3 2 1 0 |
  -- |======| |===========================================|
  -- | Free | |  Reserv. |  R  G  B |      vert. pos.     |
  -- |------| |-------------------------------------------|
  --


  p_rw0_port : process (i_clockA)
  begin
    if rising_edge(i_clockA) then
      if (true) then
        if (i_WEA = '1') then
          v_ram(conv_integer(i_ADDRA)) := i_DIA;
        end if;
        --o_DOA <= v_ram(conv_integer(i_ADDRA));
      end if;
    end if;
  end process;

  p_rw1_port : process (i_clockB)
  begin
    if rising_edge(i_clockB) then
      if (true) then
        o_DOB <= v_ram(conv_integer(i_ADDRB));
        if (i_WEB = '1') then
          v_ram(conv_integer(i_ADDRB)) := i_DIB;
        end if;
      end if;
    end if;
  end process;

end Behavioral;
