-------------------------------------------------------------------------------
--
-- The Data memory controller.
--
-- $Id: t400_dmem_ctrl-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_dmem_ctrl_rtl_c0 of t400_dmem_ctrl is

  for rtl
  end for;

end t400_dmem_ctrl_rtl_c0;
