-------------------------------------------------------------------------------
--
-- GCpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: gcpad_sampler-c.vhd 41 2009-04-01 19:58:04Z arniml $
--
-------------------------------------------------------------------------------

configuration gcpad_sampler_rtl_c0 of gcpad_sampler is

  for rtl
  end for;

end gcpad_sampler_rtl_c0;
