-- MultiIO enable 
  constant CFG_MULTIIO  : integer := CONFIG_MULTIIO_ENABLE;

