000000 => x"bc0b", -- B
000001 => x"bc04", -- B
000002 => x"bc03", -- B
000003 => x"bc02", -- B
000004 => x"bc01", -- B
000005 => x"be73", -- BL
000006 => x"c578", -- LDIL
000007 => x"c906", -- LDIH
000008 => x"be7f", -- BL
000009 => x"be6f", -- BL
000010 => x"bc00", -- B
000011 => x"c724", -- LDIL
000012 => x"cb07", -- LDIH
000013 => x"c114", -- LDIL
000014 => x"c907", -- LDIH
000015 => x"be78", -- BL
000016 => x"c47f", -- LDIL
000017 => x"ec0b", -- MCR
000018 => x"c002", -- LDIL
000019 => x"ec0c", -- MCR
000020 => x"c400", -- LDIL
000021 => x"c800", -- LDIH
000022 => x"c7e6", -- LDIL
000023 => x"cb82", -- LDIH
000024 => x"3474", -- GTL
000025 => x"6c6a", -- PUSH
000026 => x"c6f8", -- LDIL
000027 => x"ca83", -- LDIH
000028 => x"c578", -- LDIL
000029 => x"c904", -- LDIH
000030 => x"29b3", -- CLR
000031 => x"785a", -- LDR
000032 => x"c080", -- LDIL
000033 => x"526a", -- PEEK
000034 => x"c7c4", -- LDIL
000035 => x"cb82", -- LDIH
000036 => x"3474", -- GTL
000037 => x"01b1", -- INC
000038 => x"c400", -- LDIL
000039 => x"c800", -- LDIH
000040 => x"1838", -- CMP
000041 => x"85f6", -- BNE
000042 => x"586a", -- POP
000043 => x"2ad5", -- CLR
000044 => x"ec5a", -- MCR
000045 => x"c478", -- LDIL
000046 => x"c804", -- LDIH
000047 => x"c480", -- LDIL
000048 => x"c880", -- LDIH
000049 => x"c578", -- LDIL
000050 => x"c902", -- LDIH
000051 => x"be5e", -- BL
000052 => x"ee02", -- MRC
000053 => x"be1a", -- BL
000054 => x"be42", -- BL
000055 => x"c6f8", -- LDIL
000056 => x"ca84", -- LDIH
000057 => x"c580", -- LDIL
000058 => x"c980", -- LDIH
000059 => x"7a5a", -- LDR
000060 => x"be13", -- BL
000061 => x"c0a0", -- LDIL
000062 => x"be07", -- BL
000063 => x"7a5a", -- LDR
000064 => x"be0f", -- BL
000065 => x"be37", -- BL
000066 => x"05b9", -- DECS
000067 => x"85f8", -- BNE
000068 => x"bc00", -- B
000069 => x"ec22", -- MRC
000070 => x"dc05", -- STB
000071 => x"b9fe", -- BTS
000072 => x"ed18", -- MCR
000073 => x"3470", -- RET
000074 => x"ec20", -- MRC
000075 => x"dc8f", -- STBI
000076 => x"b9fe", -- BTS
000077 => x"c800", -- LDIH
000078 => x"3470", -- RET
000079 => x"6c6a", -- PUSH
000080 => x"6cea", -- PUSH
000081 => x"6d6a", -- PUSH
000082 => x"6dea", -- PUSH
000083 => x"6e6a", -- PUSH
000084 => x"6fea", -- PUSH
000085 => x"3d42", -- SFT
000086 => x"3d22", -- SFT
000087 => x"3d22", -- SFT
000088 => x"3d22", -- SFT
000089 => x"be15", -- BL
000090 => x"bfeb", -- BL
000091 => x"3d40", -- SFT
000092 => x"be12", -- BL
000093 => x"bfe8", -- BL
000094 => x"3d45", -- SFT
000095 => x"3d25", -- SFT
000096 => x"3d25", -- SFT
000097 => x"3d25", -- SFT
000098 => x"be0c", -- BL
000099 => x"bfe2", -- BL
000100 => x"0140", -- MOV
000101 => x"be09", -- BL
000102 => x"bfdf", -- BL
000103 => x"5bea", -- POP
000104 => x"5a6a", -- POP
000105 => x"59ea", -- POP
000106 => x"596a", -- POP
000107 => x"58ea", -- POP
000108 => x"586a", -- POP
000109 => x"3470", -- RET
000110 => x"c08f", -- LDIL
000111 => x"2121", -- AND
000112 => x"c089", -- LDIL
000113 => x"181a", -- CMP
000114 => x"8803", -- BCS
000115 => x"c0b0", -- LDIL
000116 => x"bc02", -- B
000117 => x"c0b7", -- LDIL
000118 => x"0892", -- ADD
000119 => x"3470", -- RET
000120 => x"6c6a", -- PUSH
000121 => x"6cea", -- PUSH
000122 => x"6d6a", -- PUSH
000123 => x"6fea", -- PUSH
000124 => x"0170", -- MOV
000125 => x"c08d", -- LDIL
000126 => x"bfc7", -- BL
000127 => x"c08a", -- LDIL
000128 => x"03a0", -- MOV
000129 => x"bfc4", -- BL
000130 => x"5bea", -- POP
000131 => x"596a", -- POP
000132 => x"58ea", -- POP
000133 => x"586a", -- POP
000134 => x"3470", -- RET
000135 => x"0270", -- MOV
000136 => x"7829", -- LDR
000137 => x"c080", -- LDIL
000138 => x"ccff", -- LDIH
000139 => x"2081", -- AND
000140 => x"3c98", -- SFTS
000141 => x"8003", -- BEQ
000142 => x"bfb7", -- BL
000143 => x"bdf9", -- B
000144 => x"3440", -- RET
000145 => x"6eea", -- PUSH
000146 => x"6e6a", -- PUSH
000147 => x"6dea", -- PUSH
000148 => x"6d6a", -- PUSH
000149 => x"6cea", -- PUSH
000150 => x"6c6a", -- PUSH
000151 => x"6fea", -- PUSH
000152 => x"c3b6", -- LDIL
000153 => x"cb82", -- LDIH
000154 => x"447e", -- STR
000155 => x"44fa", -- STR
000156 => x"457c", -- STR
000157 => x"2800", -- CLR
000158 => x"3c95", -- SFT
000159 => x"3419", -- TEQ
000160 => x"8003", -- BEQ
000161 => x"0001", -- INC
000162 => x"bdfc", -- B
000163 => x"c3b6", -- LDIL
000164 => x"cb82", -- LDIH
000165 => x"5478", -- STR
000166 => x"c3b6", -- LDIL
000167 => x"cb82", -- LDIH
000168 => x"c281", -- LDIL
000169 => x"56fa", -- STR
000170 => x"56fc", -- STR
000171 => x"56fe", -- STR
000172 => x"c3be", -- LDIL
000173 => x"cb82", -- LDIH
000174 => x"c280", -- LDIL
000175 => x"56f8", -- STR
000176 => x"c3ba", -- LDIL
000177 => x"cb82", -- LDIH
000178 => x"40fa", -- LDR
000179 => x"5178", -- LDR
000180 => x"0521", -- DEC
000181 => x"c204", -- LDIL
000182 => x"3e44", -- SFT
000183 => x"0499", -- DECS
000184 => x"85fe", -- BNE
000185 => x"f124", -- MUL
000186 => x"557c", -- STR
000187 => x"c3b6", -- LDIL
000188 => x"cb82", -- LDIH
000189 => x"427e", -- LDR
000190 => x"50fa", -- LDR
000191 => x"517e", -- LDR
000192 => x"41fc", -- LDR
000193 => x"0521", -- DEC
000194 => x"3d24", -- SFT
000195 => x"3d24", -- SFT
000196 => x"0932", -- ADD
000197 => x"c3be", -- LDIL
000198 => x"cb82", -- LDIH
000199 => x"5078", -- LDR
000200 => x"0804", -- ADD
000201 => x"c182", -- LDIL
000202 => x"3db4", -- SFT
000203 => x"0499", -- DECS
000204 => x"85fe", -- BNE
000205 => x"0883", -- ADD
000206 => x"c3c0", -- LDIL
000207 => x"cb82", -- LDIH
000208 => x"5478", -- STR
000209 => x"54fa", -- STR
000210 => x"557c", -- STR
000211 => x"0180", -- MOV
000212 => x"0210", -- MOV
000213 => x"02a0", -- MOV
000214 => x"6dea", -- PUSH
000215 => x"6e6a", -- PUSH
000216 => x"5038", -- LDR
000217 => x"50ba", -- LDR
000218 => x"5148", -- LDR
000219 => x"51ca", -- LDR
000220 => x"5258", -- LDR
000221 => x"52da", -- LDR
000222 => x"be45", -- BL
000223 => x"5aea", -- POP
000224 => x"5a6a", -- POP
000225 => x"5558", -- STR
000226 => x"55da", -- STR
000227 => x"5448", -- STR
000228 => x"54ca", -- STR
000229 => x"c3be", -- LDIL
000230 => x"cb82", -- LDIH
000231 => x"5078", -- LDR
000232 => x"c084", -- LDIL
000233 => x"0801", -- ADD
000234 => x"5478", -- STR
000235 => x"c3b6", -- LDIL
000236 => x"cb82", -- LDIH
000237 => x"507a", -- LDR
000238 => x"517e", -- LDR
000239 => x"c081", -- LDIL
000240 => x"0409", -- DECS
000241 => x"8003", -- BEQ
000242 => x"3c94", -- SFT
000243 => x"bdfd", -- B
000244 => x"181a", -- CMP
000245 => x"0121", -- INC
000246 => x"557e", -- STR
000247 => x"85c4", -- BNE
000248 => x"c101", -- LDIL
000249 => x"557e", -- STR
000250 => x"c3b6", -- LDIL
000251 => x"cb82", -- LDIH
000252 => x"407a", -- LDR
000253 => x"50fa", -- LDR
000254 => x"517c", -- LDR
000255 => x"3c05", -- SFT
000256 => x"0499", -- DECS
000257 => x"85fe", -- BNE
000258 => x"180a", -- CMP
000259 => x"0121", -- INC
000260 => x"557c", -- STR
000261 => x"85ab", -- BNE
000262 => x"c101", -- LDIL
000263 => x"557c", -- STR
000264 => x"c3b6", -- LDIL
000265 => x"cb82", -- LDIH
000266 => x"5078", -- LDR
000267 => x"50fa", -- LDR
000268 => x"1809", -- CMP
000269 => x"0091", -- INC
000270 => x"54fa", -- STR
000271 => x"85a1", -- BNE
000272 => x"5bea", -- POP
000273 => x"586a", -- POP
000274 => x"58ea", -- POP
000275 => x"596a", -- POP
000276 => x"59ea", -- POP
000277 => x"5a6a", -- POP
000278 => x"5aea", -- POP
000279 => x"3470", -- RET
000280 => x"0000", -- NOP
000281 => x"0000", -- NOP
000282 => x"0000", -- NOP
000283 => x"0000", -- NOP
000284 => x"0000", -- NOP
000285 => x"0000", -- NOP
000286 => x"0000", -- NOP
000287 => x"0000", -- NOP
000288 => x"0000", -- NOP
000289 => x"0000", -- NOP
000290 => x"0000", -- NOP
000291 => x"6fea", -- PUSH
000292 => x"6c6a", -- PUSH
000293 => x"6cea", -- PUSH
000294 => x"c7bc", -- LDIL
000295 => x"cb82", -- LDIH
000296 => x"f042", -- MUL
000297 => x"f0ca", -- MULH
000298 => x"3c0c", -- SFTS
000299 => x"3c92", -- SFT
000300 => x"3c0c", -- SFTS
000301 => x"3c92", -- SFT
000302 => x"54f8", -- STR
000303 => x"f043", -- MUL
000304 => x"f0cb", -- MULH
000305 => x"3c0c", -- SFTS
000306 => x"3c92", -- SFT
000307 => x"3c0c", -- SFTS
000308 => x"3c92", -- SFT
000309 => x"54fa", -- STR
000310 => x"f052", -- MUL
000311 => x"f0da", -- MULH
000312 => x"3c0c", -- SFTS
000313 => x"3c92", -- SFT
000314 => x"3c0c", -- SFTS
000315 => x"3c92", -- SFT
000316 => x"54fc", -- STR
000317 => x"f053", -- MUL
000318 => x"f0db", -- MULH
000319 => x"3c0c", -- SFTS
000320 => x"3c92", -- SFT
000321 => x"3c0c", -- SFTS
000322 => x"3c92", -- SFT
000323 => x"54fe", -- STR
000324 => x"58ea", -- POP
000325 => x"586a", -- POP
000326 => x"5178", -- LDR
000327 => x"51fe", -- LDR
000328 => x"090a", -- ADDS
000329 => x"15a3", -- SBC
000330 => x"6dea", -- PUSH
000331 => x"517a", -- LDR
000332 => x"51fc", -- LDR
000333 => x"091a", -- ADDS
000334 => x"0da3", -- ADC
000335 => x"6dea", -- PUSH
000336 => x"5178", -- LDR
000337 => x"51fe", -- LDR
000338 => x"110a", -- SUBS
000339 => x"0da3", -- ADC
000340 => x"6dea", -- PUSH
000341 => x"517a", -- LDR
000342 => x"51fc", -- LDR
000343 => x"111a", -- SUBS
000344 => x"15a3", -- SBC
000345 => x"596a", -- POP
000346 => x"58ea", -- POP
000347 => x"586a", -- POP
000348 => x"5bea", -- POP
000349 => x"3470", -- RET
000350 => x"0000", -- NOP
000351 => x"0000", -- NOP
000352 => x"0000", -- NOP
000353 => x"0000", -- NOP
000354 => x"6dea", -- PUSH
000355 => x"6e6a", -- PUSH
000356 => x"6eea", -- PUSH
000357 => x"2ad5", -- CLR
000358 => x"3dbd", -- SFTS
000359 => x"3ed6", -- SFT
000360 => x"0649", -- DECS
000361 => x"85fd", -- BNE
000362 => x"3ed4", -- SFT
000363 => x"3ed4", -- SFT
000364 => x"0aa5", -- ADD
000365 => x"5458", -- STR
000366 => x"54da", -- STR
000367 => x"5aea", -- POP
000368 => x"5a6a", -- POP
000369 => x"59ea", -- POP
000370 => x"3470", -- RET
000371 => x"6cea", -- PUSH
000372 => x"2891", -- CLR
000373 => x"3c0d", -- SFTS
000374 => x"8003", -- BEQ
000375 => x"0091", -- INC
000376 => x"bdfd", -- B
000377 => x"0010", -- MOV
000378 => x"58ea", -- POP
000379 => x"3470", -- RET
000380 => x"4000", -- .DW
000381 => x"0000", -- .DW
000382 => x"3fec", -- .DW
000383 => x"0323", -- .DW
000384 => x"3fb1", -- .DW
000385 => x"0645", -- .DW
000386 => x"3f4e", -- .DW
000387 => x"0964", -- .DW
000388 => x"3ec5", -- .DW
000389 => x"0c7c", -- .DW
000390 => x"3e14", -- .DW
000391 => x"0f8c", -- .DW
000392 => x"3d3e", -- .DW
000393 => x"1294", -- .DW
000394 => x"3c42", -- .DW
000395 => x"158f", -- .DW
000396 => x"3b20", -- .DW
000397 => x"187d", -- .DW
000398 => x"39da", -- .DW
000399 => x"1b5d", -- .DW
000400 => x"3871", -- .DW
000401 => x"1e2b", -- .DW
000402 => x"36e5", -- .DW
000403 => x"20e7", -- .DW
000404 => x"3536", -- .DW
000405 => x"238e", -- .DW
000406 => x"3367", -- .DW
000407 => x"261f", -- .DW
000408 => x"3179", -- .DW
000409 => x"2899", -- .DW
000410 => x"2f6b", -- .DW
000411 => x"2afa", -- .DW
000412 => x"2d41", -- .DW
000413 => x"2d41", -- .DW
000414 => x"2afa", -- .DW
000415 => x"2f6b", -- .DW
000416 => x"2899", -- .DW
000417 => x"3179", -- .DW
000418 => x"261f", -- .DW
000419 => x"3367", -- .DW
000420 => x"238e", -- .DW
000421 => x"3536", -- .DW
000422 => x"20e7", -- .DW
000423 => x"36e5", -- .DW
000424 => x"1e2b", -- .DW
000425 => x"3871", -- .DW
000426 => x"1b5d", -- .DW
000427 => x"39da", -- .DW
000428 => x"187d", -- .DW
000429 => x"3b20", -- .DW
000430 => x"158f", -- .DW
000431 => x"3c42", -- .DW
000432 => x"1294", -- .DW
000433 => x"3d3e", -- .DW
000434 => x"0f8c", -- .DW
000435 => x"3e14", -- .DW
000436 => x"0c7c", -- .DW
000437 => x"3ec5", -- .DW
000438 => x"0964", -- .DW
000439 => x"3f4e", -- .DW
000440 => x"0645", -- .DW
000441 => x"3fb1", -- .DW
000442 => x"0323", -- .DW
000443 => x"3fec", -- .DW
000444 => x"0000", -- .DW
000445 => x"4000", -- .DW
000446 => x"fcdd", -- .DW
000447 => x"3fec", -- .DW
000448 => x"f9bb", -- .DW
000449 => x"3fb1", -- .DW
000450 => x"f69c", -- .DW
000451 => x"3f4e", -- .DW
000452 => x"f384", -- .DW
000453 => x"3ec5", -- .DW
000454 => x"f074", -- .DW
000455 => x"3e14", -- .DW
000456 => x"ed6c", -- .DW
000457 => x"3d3e", -- .DW
000458 => x"ea71", -- .DW
000459 => x"3c42", -- .DW
000460 => x"e783", -- .DW
000461 => x"3b20", -- .DW
000462 => x"e4a3", -- .DW
000463 => x"39da", -- .DW
000464 => x"e1d5", -- .DW
000465 => x"3871", -- .DW
000466 => x"df19", -- .DW
000467 => x"36e5", -- .DW
000468 => x"dc72", -- .DW
000469 => x"3536", -- .DW
000470 => x"d9e1", -- .DW
000471 => x"3367", -- .DW
000472 => x"d767", -- .DW
000473 => x"3179", -- .DW
000474 => x"d506", -- .DW
000475 => x"2f6b", -- .DW
000476 => x"d2bf", -- .DW
000477 => x"2d41", -- .DW
000478 => x"d095", -- .DW
000479 => x"2afa", -- .DW
000480 => x"ce87", -- .DW
000481 => x"2899", -- .DW
000482 => x"cc99", -- .DW
000483 => x"261f", -- .DW
000484 => x"caca", -- .DW
000485 => x"238e", -- .DW
000486 => x"c91b", -- .DW
000487 => x"20e7", -- .DW
000488 => x"c78f", -- .DW
000489 => x"1e2b", -- .DW
000490 => x"c626", -- .DW
000491 => x"1b5d", -- .DW
000492 => x"c4e0", -- .DW
000493 => x"187d", -- .DW
000494 => x"c3be", -- .DW
000495 => x"158f", -- .DW
000496 => x"c2c2", -- .DW
000497 => x"1294", -- .DW
000498 => x"c1ec", -- .DW
000499 => x"0f8c", -- .DW
000500 => x"c13b", -- .DW
000501 => x"0c7c", -- .DW
000502 => x"c0b2", -- .DW
000503 => x"0964", -- .DW
000504 => x"c04f", -- .DW
000505 => x"0645", -- .DW
000506 => x"c014", -- .DW
000507 => x"0323", -- .DW
000508 => x"0400", -- .DW
000509 => x"0000", -- .DW
000510 => x"0000", -- .DW
000511 => x"0000", -- .DW
000512 => x"0400", -- .DW
000513 => x"0000", -- .DW
000514 => x"0000", -- .DW
000515 => x"0000", -- .DW
000516 => x"0400", -- .DW
000517 => x"0000", -- .DW
000518 => x"0000", -- .DW
000519 => x"0000", -- .DW
000520 => x"0400", -- .DW
000521 => x"0000", -- .DW
000522 => x"0000", -- .DW
000523 => x"0000", -- .DW
000524 => x"0400", -- .DW
000525 => x"0000", -- .DW
000526 => x"0000", -- .DW
000527 => x"0000", -- .DW
000528 => x"0400", -- .DW
000529 => x"0000", -- .DW
000530 => x"0000", -- .DW
000531 => x"0000", -- .DW
000532 => x"0400", -- .DW
000533 => x"0000", -- .DW
000534 => x"0000", -- .DW
000535 => x"0000", -- .DW
000536 => x"0400", -- .DW
000537 => x"0000", -- .DW
000538 => x"0000", -- .DW
000539 => x"0000", -- .DW
000540 => x"0400", -- .DW
000541 => x"0000", -- .DW
000542 => x"0000", -- .DW
000543 => x"0000", -- .DW
000544 => x"0400", -- .DW
000545 => x"0000", -- .DW
000546 => x"0000", -- .DW
000547 => x"0000", -- .DW
000548 => x"0400", -- .DW
000549 => x"0000", -- .DW
000550 => x"0000", -- .DW
000551 => x"0000", -- .DW
000552 => x"0400", -- .DW
000553 => x"0000", -- .DW
000554 => x"0000", -- .DW
000555 => x"0000", -- .DW
000556 => x"0400", -- .DW
000557 => x"0000", -- .DW
000558 => x"0000", -- .DW
000559 => x"0000", -- .DW
000560 => x"0400", -- .DW
000561 => x"0000", -- .DW
000562 => x"0000", -- .DW
000563 => x"0000", -- .DW
000564 => x"0400", -- .DW
000565 => x"0000", -- .DW
000566 => x"0000", -- .DW
000567 => x"0000", -- .DW
000568 => x"0400", -- .DW
000569 => x"0000", -- .DW
000570 => x"0000", -- .DW
000571 => x"0000", -- .DW
000572 => x"0400", -- .DW
000573 => x"0000", -- .DW
000574 => x"0000", -- .DW
000575 => x"0000", -- .DW
000576 => x"0400", -- .DW
000577 => x"0000", -- .DW
000578 => x"0000", -- .DW
000579 => x"0000", -- .DW
000580 => x"0400", -- .DW
000581 => x"0000", -- .DW
000582 => x"0000", -- .DW
000583 => x"0000", -- .DW
000584 => x"0400", -- .DW
000585 => x"0000", -- .DW
000586 => x"0000", -- .DW
000587 => x"0000", -- .DW
000588 => x"0400", -- .DW
000589 => x"0000", -- .DW
000590 => x"0000", -- .DW
000591 => x"0000", -- .DW
000592 => x"0400", -- .DW
000593 => x"0000", -- .DW
000594 => x"0000", -- .DW
000595 => x"0000", -- .DW
000596 => x"0400", -- .DW
000597 => x"0000", -- .DW
000598 => x"0000", -- .DW
000599 => x"0000", -- .DW
000600 => x"0400", -- .DW
000601 => x"0000", -- .DW
000602 => x"0000", -- .DW
000603 => x"0000", -- .DW
000604 => x"0400", -- .DW
000605 => x"0000", -- .DW
000606 => x"0000", -- .DW
000607 => x"0000", -- .DW
000608 => x"0400", -- .DW
000609 => x"0000", -- .DW
000610 => x"0000", -- .DW
000611 => x"0000", -- .DW
000612 => x"0400", -- .DW
000613 => x"0000", -- .DW
000614 => x"0000", -- .DW
000615 => x"0000", -- .DW
000616 => x"0400", -- .DW
000617 => x"0000", -- .DW
000618 => x"0000", -- .DW
000619 => x"0000", -- .DW
000620 => x"0400", -- .DW
000621 => x"0000", -- .DW
000622 => x"0000", -- .DW
000623 => x"0000", -- .DW
000624 => x"0400", -- .DW
000625 => x"0000", -- .DW
000626 => x"0000", -- .DW
000627 => x"0000", -- .DW
000628 => x"0400", -- .DW
000629 => x"0000", -- .DW
000630 => x"0000", -- .DW
000631 => x"0000", -- .DW
000632 => x"0400", -- .DW
000633 => x"0000", -- .DW
000634 => x"0000", -- .DW
000635 => x"0000", -- .DW
000636 => x"0000", -- NOP
000637 => x"0000", -- NOP
000638 => x"0000", -- NOP
000639 => x"0000", -- NOP
000640 => x"0000", -- NOP
000641 => x"0000", -- NOP
000642 => x"0000", -- NOP
000643 => x"0000", -- NOP
000644 => x"0000", -- NOP
000645 => x"0000", -- NOP
000646 => x"0000", -- NOP
000647 => x"0000", -- NOP
000648 => x"0000", -- NOP
000649 => x"0000", -- NOP
000650 => x"0000", -- NOP
000651 => x"0000", -- NOP
000652 => x"0000", -- NOP
000653 => x"0000", -- NOP
000654 => x"0000", -- NOP
000655 => x"0000", -- NOP
000656 => x"0000", -- NOP
000657 => x"0000", -- NOP
000658 => x"0000", -- NOP
000659 => x"0000", -- NOP
000660 => x"0000", -- NOP
000661 => x"0000", -- NOP
000662 => x"0000", -- NOP
000663 => x"0000", -- NOP
000664 => x"0000", -- NOP
000665 => x"0000", -- NOP
000666 => x"0000", -- NOP
000667 => x"0000", -- NOP
000668 => x"0000", -- NOP
000669 => x"0000", -- NOP
000670 => x"0000", -- NOP
000671 => x"0000", -- NOP
000672 => x"0000", -- NOP
000673 => x"0000", -- NOP
000674 => x"0000", -- NOP
000675 => x"0000", -- NOP
000676 => x"0000", -- NOP
000677 => x"0000", -- NOP
000678 => x"0000", -- NOP
000679 => x"0000", -- NOP
000680 => x"0000", -- NOP
000681 => x"0000", -- NOP
000682 => x"0000", -- NOP
000683 => x"0000", -- NOP
000684 => x"0000", -- NOP
000685 => x"0000", -- NOP
000686 => x"0000", -- NOP
000687 => x"0000", -- NOP
000688 => x"0000", -- NOP
000689 => x"0000", -- NOP
000690 => x"0000", -- NOP
000691 => x"0000", -- NOP
000692 => x"0000", -- NOP
000693 => x"0000", -- NOP
000694 => x"0000", -- NOP
000695 => x"0000", -- NOP
000696 => x"0000", -- NOP
000697 => x"0000", -- NOP
000698 => x"0000", -- NOP
000699 => x"0000", -- NOP
000700 => x"0000", -- NOP
000701 => x"0000", -- NOP
000702 => x"0000", -- NOP
000703 => x"0000", -- NOP
000704 => x"0000", -- NOP
000705 => x"0000", -- NOP
000706 => x"0000", -- NOP
000707 => x"0000", -- NOP
000708 => x"0000", -- NOP
000709 => x"0000", -- NOP
000710 => x"0000", -- NOP
000711 => x"0000", -- NOP
000712 => x"0000", -- NOP
000713 => x"0000", -- NOP
000714 => x"0000", -- NOP
000715 => x"0000", -- NOP
000716 => x"0000", -- NOP
000717 => x"0000", -- NOP
000718 => x"0000", -- NOP
000719 => x"0000", -- NOP
000720 => x"0000", -- NOP
000721 => x"0000", -- NOP
000722 => x"0000", -- NOP
000723 => x"0000", -- NOP
000724 => x"0000", -- NOP
000725 => x"0000", -- NOP
000726 => x"0000", -- NOP
000727 => x"0000", -- NOP
000728 => x"0000", -- NOP
000729 => x"0000", -- NOP
000730 => x"0000", -- NOP
000731 => x"0000", -- NOP
000732 => x"0000", -- NOP
000733 => x"0000", -- NOP
000734 => x"0000", -- NOP
000735 => x"0000", -- NOP
000736 => x"0000", -- NOP
000737 => x"0000", -- NOP
000738 => x"0000", -- NOP
000739 => x"0000", -- NOP
000740 => x"0000", -- NOP
000741 => x"0000", -- NOP
000742 => x"0000", -- NOP
000743 => x"0000", -- NOP
000744 => x"0000", -- NOP
000745 => x"0000", -- NOP
000746 => x"0000", -- NOP
000747 => x"0000", -- NOP
000748 => x"0000", -- NOP
000749 => x"0000", -- NOP
000750 => x"0000", -- NOP
000751 => x"0000", -- NOP
000752 => x"0000", -- NOP
000753 => x"0000", -- NOP
000754 => x"0000", -- NOP
000755 => x"0000", -- NOP
000756 => x"0000", -- NOP
000757 => x"0000", -- NOP
000758 => x"0000", -- NOP
000759 => x"0000", -- NOP
000760 => x"0000", -- NOP
000761 => x"0000", -- NOP
000762 => x"0000", -- NOP
000763 => x"0000", -- NOP
000764 => x"0000", -- NOP
000765 => x"0000", -- NOP
000766 => x"0000", -- NOP
000767 => x"0000", -- NOP
000768 => x"0000", -- NOP
000769 => x"0000", -- NOP
000770 => x"0000", -- NOP
000771 => x"0000", -- NOP
000772 => x"0000", -- NOP
000773 => x"0000", -- NOP
000774 => x"0000", -- NOP
000775 => x"0000", -- NOP
000776 => x"0000", -- NOP
000777 => x"0000", -- NOP
000778 => x"0000", -- NOP
000779 => x"0000", -- NOP
000780 => x"0000", -- NOP
000781 => x"0000", -- NOP
000782 => x"0000", -- NOP
000783 => x"0000", -- NOP
000784 => x"0000", -- NOP
000785 => x"0000", -- NOP
000786 => x"0000", -- NOP
000787 => x"0000", -- NOP
000788 => x"0000", -- NOP
000789 => x"0000", -- NOP
000790 => x"0000", -- NOP
000791 => x"0000", -- NOP
000792 => x"0000", -- NOP
000793 => x"0000", -- NOP
000794 => x"0000", -- NOP
000795 => x"0000", -- NOP
000796 => x"0000", -- NOP
000797 => x"0000", -- NOP
000798 => x"0000", -- NOP
000799 => x"0000", -- NOP
000800 => x"0000", -- NOP
000801 => x"0000", -- NOP
000802 => x"0000", -- NOP
000803 => x"0000", -- NOP
000804 => x"0000", -- NOP
000805 => x"0000", -- NOP
000806 => x"0000", -- NOP
000807 => x"0000", -- NOP
000808 => x"0000", -- NOP
000809 => x"0000", -- NOP
000810 => x"0000", -- NOP
000811 => x"0000", -- NOP
000812 => x"0000", -- NOP
000813 => x"0000", -- NOP
000814 => x"0000", -- NOP
000815 => x"0000", -- NOP
000816 => x"0000", -- NOP
000817 => x"0000", -- NOP
000818 => x"0000", -- NOP
000819 => x"0000", -- NOP
000820 => x"0000", -- NOP
000821 => x"0000", -- NOP
000822 => x"0000", -- NOP
000823 => x"0000", -- NOP
000824 => x"0000", -- NOP
000825 => x"0000", -- NOP
000826 => x"0000", -- NOP
000827 => x"0000", -- NOP
000828 => x"0000", -- NOP
000829 => x"0000", -- NOP
000830 => x"0000", -- NOP
000831 => x"0000", -- NOP
000832 => x"0000", -- NOP
000833 => x"0000", -- NOP
000834 => x"0000", -- NOP
000835 => x"0000", -- NOP
000836 => x"0000", -- NOP
000837 => x"0000", -- NOP
000838 => x"0000", -- NOP
000839 => x"0000", -- NOP
000840 => x"0000", -- NOP
000841 => x"0000", -- NOP
000842 => x"0000", -- NOP
000843 => x"0000", -- NOP
000844 => x"0000", -- NOP
000845 => x"0000", -- NOP
000846 => x"0000", -- NOP
000847 => x"0000", -- NOP
000848 => x"0000", -- NOP
000849 => x"0000", -- NOP
000850 => x"0000", -- NOP
000851 => x"0000", -- NOP
000852 => x"0000", -- NOP
000853 => x"0000", -- NOP
000854 => x"0000", -- NOP
000855 => x"0000", -- NOP
000856 => x"0000", -- NOP
000857 => x"0000", -- NOP
000858 => x"0000", -- NOP
000859 => x"0000", -- NOP
000860 => x"0000", -- NOP
000861 => x"0000", -- NOP
000862 => x"0000", -- NOP
000863 => x"0000", -- NOP
000864 => x"0000", -- NOP
000865 => x"0000", -- NOP
000866 => x"0000", -- NOP
000867 => x"0000", -- NOP
000868 => x"0000", -- NOP
000869 => x"0000", -- NOP
000870 => x"0000", -- NOP
000871 => x"0000", -- NOP
000872 => x"0000", -- NOP
000873 => x"0000", -- NOP
000874 => x"0000", -- NOP
000875 => x"0000", -- NOP
000876 => x"0000", -- NOP
000877 => x"0000", -- NOP
000878 => x"0000", -- NOP
000879 => x"0000", -- NOP
000880 => x"0000", -- NOP
000881 => x"0000", -- NOP
000882 => x"0000", -- NOP
000883 => x"0000", -- NOP
000884 => x"0000", -- NOP
000885 => x"0000", -- NOP
000886 => x"0000", -- NOP
000887 => x"0000", -- NOP
000888 => x"0000", -- NOP
000889 => x"0000", -- NOP
000890 => x"0000", -- NOP
000891 => x"0000", -- NOP
000892 => x"4578", -- .DW
000893 => x"6365", -- .DW
000894 => x"7074", -- .DW
000895 => x"696f", -- .DW
000896 => x"6e2f", -- .DW
000897 => x"696e", -- .DW
000898 => x"7465", -- .DW
000899 => x"7272", -- .DW
000900 => x"7570", -- .DW
000901 => x"7420", -- .DW
000902 => x"6572", -- .DW
000903 => x"726f", -- .DW
000904 => x"7221", -- .DW
000905 => x"0000", -- .DW
000906 => x"436f", -- .DW
000907 => x"6d70", -- .DW
000908 => x"7574", -- .DW
000909 => x"696e", -- .DW
000910 => x"6720", -- .DW
000911 => x"4646", -- .DW
000912 => x"542e", -- .DW
000913 => x"2e2e", -- .DW
000914 => x"2000", -- .DW
000915 => x"0000", -- NOP
000916 => x"0000", -- NOP
000917 => x"0000", -- NOP
000918 => x"0000", -- NOP
000919 => x"0000", -- NOP
000920 => x"0000", -- NOP
000921 => x"0000", -- NOP
000922 => x"0000", -- NOP
000923 => x"0000", -- NOP
000924 => x"0000", -- NOP
000925 => x"0000", -- NOP
000926 => x"0000", -- NOP
000927 => x"0000", -- NOP
000928 => x"0000", -- NOP
000929 => x"0000", -- NOP
000930 => x"0000", -- NOP
000931 => x"0000", -- NOP
000932 => x"0000", -- NOP
000933 => x"0000", -- NOP
000934 => x"0000", -- NOP
000935 => x"0000", -- NOP
000936 => x"0000", -- NOP
000937 => x"0000", -- NOP
000938 => x"0000", -- NOP
000939 => x"0000", -- NOP
000940 => x"0000", -- NOP
000941 => x"0000", -- NOP
000942 => x"0000", -- NOP
000943 => x"0000", -- NOP
000944 => x"0000", -- NOP
000945 => x"0000", -- NOP
000946 => x"0000", -- NOP
000947 => x"0000", -- NOP
000948 => x"0000", -- NOP
000949 => x"0000", -- NOP
000950 => x"0000", -- NOP
000951 => x"0000", -- NOP
000952 => x"0000", -- NOP
000953 => x"0000", -- NOP
000954 => x"0000", -- NOP
000955 => x"0000", -- NOP
000956 => x"0000", -- NOP
000957 => x"0000", -- NOP
000958 => x"0000", -- NOP
000959 => x"0000", -- NOP
000960 => x"0000", -- NOP
000961 => x"0000", -- NOP
000962 => x"0000", -- NOP
000963 => x"0000", -- NOP
000964 => x"0000", -- NOP
000965 => x"0000", -- NOP
000966 => x"0000", -- NOP
000967 => x"0000", -- NOP
000968 => x"0000", -- NOP
000969 => x"0000", -- NOP
000970 => x"0000", -- NOP
000971 => x"0000", -- NOP
000972 => x"0000", -- NOP
000973 => x"0000", -- NOP
000974 => x"0000", -- NOP
000975 => x"0000", -- NOP
000976 => x"0000", -- NOP
000977 => x"0000", -- NOP
000978 => x"0000", -- NOP
others => x"0000"  -- NOP