000000 => x"bc0b", -- B
000001 => x"bc04", -- B
000002 => x"bc03", -- B
000003 => x"bc02", -- B
000004 => x"bc01", -- B
000005 => x"be30", -- BL
000006 => x"c10e", -- LDIL
000007 => x"c901", -- LDIH
000008 => x"be21", -- BL
000009 => x"be2c", -- BL
000010 => x"bc00", -- B
000011 => x"c12a", -- LDIL
000012 => x"c901", -- LDIH
000013 => x"be19", -- BL
000014 => x"c142", -- LDIL
000015 => x"c901", -- LDIH
000016 => x"be19", -- BL
000017 => x"be33", -- BL
000018 => x"ec4d", -- MCR
000019 => x"be22", -- BL
000020 => x"c15e", -- LDIL
000021 => x"c901", -- LDIH
000022 => x"be13", -- BL
000023 => x"be2d", -- BL
000024 => x"d24f", -- CBR
000025 => x"ec4e", -- MCR
000026 => x"be1b", -- BL
000027 => x"c0b0", -- LDIL
000028 => x"be1e", -- BL
000029 => x"c0f8", -- LDIL
000030 => x"be1c", -- BL
000031 => x"ee05", -- MRC
000032 => x"be49", -- BL
000033 => x"be14", -- BL
000034 => x"ec20", -- MRC
000035 => x"dc0f", -- STB
000036 => x"b9ea", -- BTS
000037 => x"bdf6", -- B
000038 => x"c5ff", -- LDIL
000039 => x"0270", -- MOV
000040 => x"bc03", -- B
000041 => x"29b3", -- CLR
000042 => x"0270", -- MOV
000043 => x"78a9", -- LDR
000044 => x"3c90", -- SFT
000045 => x"c880", -- LDIH
000046 => x"3419", -- TEQ
000047 => x"8003", -- BEQ
000048 => x"be0a", -- BL
000049 => x"bdfa", -- B
000050 => x"03c0", -- MOV
000051 => x"343b", -- TEQ
000052 => x"f707", -- RBAEQ
000053 => x"0170", -- MOV
000054 => x"c08d", -- LDIL
000055 => x"be03", -- BL
000056 => x"c08a", -- LDIL
000057 => x"03a0", -- MOV
000058 => x"ec22", -- MRC
000059 => x"dc05", -- STB
000060 => x"b9fe", -- BTS
000061 => x"ed18", -- MCR
000062 => x"3470", -- RET
000063 => x"ec20", -- MRC
000064 => x"dc8f", -- STBI
000065 => x"b9fe", -- BTS
000066 => x"c800", -- LDIH
000067 => x"3470", -- RET
000068 => x"0170", -- MOV
000069 => x"c200", -- LDIL
000070 => x"c184", -- LDIL
000071 => x"bff8", -- BL
000072 => x"c0c7", -- LDIL
000073 => x"1809", -- CMP
000074 => x"9003", -- BMI
000075 => x"c0a0", -- LDIL
000076 => x"1001", -- SUB
000077 => x"c0b0", -- LDIL
000078 => x"1809", -- CMP
000079 => x"91f8", -- BMI
000080 => x"c0c6", -- LDIL
000081 => x"1818", -- CMP
000082 => x"91f5", -- BMI
000083 => x"c0b9", -- LDIL
000084 => x"1818", -- CMP
000085 => x"a404", -- BLS
000086 => x"c0c1", -- LDIL
000087 => x"1809", -- CMP
000088 => x"a1ef", -- BHI
000089 => x"0080", -- MOV
000090 => x"bfe0", -- BL
000091 => x"c030", -- LDIL
000092 => x"1090", -- SUB
000093 => x"c009", -- LDIL
000094 => x"1809", -- CMP
000095 => x"a402", -- BLS
000096 => x"0497", -- DEC
000097 => x"3e42", -- SFT
000098 => x"3e42", -- SFT
000099 => x"3e42", -- SFT
000100 => x"3e42", -- SFT
000101 => x"2641", -- ORR
000102 => x"05b9", -- DECS
000103 => x"85e0", -- BNE
000104 => x"3420", -- RET
000105 => x"0370", -- MOV
000106 => x"3d42", -- SFT
000107 => x"3d22", -- SFT
000108 => x"3d22", -- SFT
000109 => x"3d22", -- SFT
000110 => x"be0f", -- BL
000111 => x"bfcb", -- BL
000112 => x"3d40", -- SFT
000113 => x"be0c", -- BL
000114 => x"bfc8", -- BL
000115 => x"3d45", -- SFT
000116 => x"3d25", -- SFT
000117 => x"3d25", -- SFT
000118 => x"3d25", -- SFT
000119 => x"be06", -- BL
000120 => x"bfc2", -- BL
000121 => x"0140", -- MOV
000122 => x"be03", -- BL
000123 => x"bfbf", -- BL
000124 => x"3460", -- RET
000125 => x"c08f", -- LDIL
000126 => x"2121", -- AND
000127 => x"c089", -- LDIL
000128 => x"181a", -- CMP
000129 => x"8803", -- BCS
000130 => x"c0b0", -- LDIL
000131 => x"bc02", -- B
000132 => x"c0b7", -- LDIL
000133 => x"0892", -- ADD
000134 => x"3470", -- RET
000135 => x"4578", -- .DW
000136 => x"6365", -- .DW
000137 => x"7074", -- .DW
000138 => x"696f", -- .DW
000139 => x"6e2f", -- .DW
000140 => x"696e", -- .DW
000141 => x"7465", -- .DW
000142 => x"7272", -- .DW
000143 => x"7570", -- .DW
000144 => x"7420", -- .DW
000145 => x"6572", -- .DW
000146 => x"726f", -- .DW
000147 => x"7221", -- .DW
000148 => x"0000", -- .DW
000149 => x"5261", -- .DW
000150 => x"6e64", -- .DW
000151 => x"6f6d", -- .DW
000152 => x"204e", -- .DW
000153 => x"756d", -- .DW
000154 => x"6265", -- .DW
000155 => x"7220", -- .DW
000156 => x"4765", -- .DW
000157 => x"6e65", -- .DW
000158 => x"7261", -- .DW
000159 => x"746f", -- .DW
000160 => x"7200", -- .DW
000161 => x"456e", -- .DW
000162 => x"7465", -- .DW
000163 => x"7220", -- .DW
000164 => x"4c46", -- .DW
000165 => x"5352", -- .DW
000166 => x"2073", -- .DW
000167 => x"6565", -- .DW
000168 => x"6420", -- .DW
000169 => x"2834", -- .DW
000170 => x"6865", -- .DW
000171 => x"7829", -- .DW
000172 => x"3a20", -- .DW
000173 => x"3078", -- .DW
000174 => x"0000", -- .DW
000175 => x"456e", -- .DW
000176 => x"7465", -- .DW
000177 => x"7220", -- .DW
000178 => x"4c46", -- .DW
000179 => x"5352", -- .DW
000180 => x"2074", -- .DW
000181 => x"6170", -- .DW
000182 => x"7320", -- .DW
000183 => x"2834", -- .DW
000184 => x"6865", -- .DW
000185 => x"7829", -- .DW
000186 => x"3a20", -- .DW
000187 => x"3078", -- .DW
000188 => x"0000", -- .DW
others => x"0000"  -- NOP