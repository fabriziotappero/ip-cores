`timescale  1 ns / 1 ps

module glbl ();

    wire GR;
    wire GSR;
    wire GTS;
    wire PRLD;

endmodule
