-- Xilinx VHDL produced by program ngd2vhdl, Version M1.3.7
-- Date: Thu Jun 11 15:24:08 1998
-- Design file: processor.pcf.nga
-- Device: 4013epg223-4
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;
architecture STRUCTURE of PROCESSOR_E is
  signal RST , NET4 , N126 , N308 , N309 , N310 , N311 , N312 , N313 , N314 , 
  N315 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 
  , N85 , N86 , N87 , N88 , N316 , N317 , N318 , N319 , N320 , N321 , N322 , 
  N323 , N324 , N325 , N326 , N327 , N328 , N329 , N330 , N331 , N332 , N333 , 
  N334 , N335 , N336 , N337 , N338 , N339 , N340 , N341 , N342 , N343 , N344 , 
  N345 , N346 , N347 , N348 , N349 , N350 , N351 , N125 , N127 , N128 , 
  IFU_N135 , JDEC , IFU_N136 , EN , SEC_B , IDU_N62 , IDU_N61 , IDU_N60 , 
  IDU_N64 , IDU_N66 , IDU_N67 , IDU_N68 , IDU_N65 , IDU_N69 , IDU_N71 , IDU_N90 
  , IDU_N89 , IDU_N93 , IDU_N92 , IDU_N97 , IDU_N100 , IDU_N99 , IDU_N98 , 
  IDU_N101 , IDU_N102 , IDU_N103 , IDU_N104 , IDU_N105 , PSU_STEP1 , PSU_N91 , 
  PSU_GO_A , PSU_EN_1 , PSU_GO_A29 , PSU_STEP2 , ALU_N474 , ALU_N575 , 
  ALU_N_2432 , ALU_N491 , ALU_N_2164 , ALU_N492 , ALU_N493 , ALU_N494 , 
  ALU_N496 , ALU_N495 , ALU_N497 , ALU_N498 , ALU_N499 , ALU_N500 , ALU_N501 , 
  ALU_N502 , ALU_N503 , ALU_N504 , ALU_N505 , ALU_N507 , ALU_N508 , ALU_N509 , 
  ALU_N511 , ALU_N512 , ALU_N513 , ALU_N515 , ALU_N516 , ALU_N517 , ALU_N519 , 
  ALU_N520 , ALU_N521 , ALU_N523 , ALU_N524 , ALU_N525 , ALU_N527 , ALU_N528 , 
  ALU_N529 , ALU_N531 , ALU_N532 , ALU_N533 , ALU_N534 , ALU_N535 , ALU_N536 , 
  ALU_N538 , ALU_N539 , ALU_N540 , ALU_N541 , ALU_N542 , ALU_N543 , ALU_N544 , 
  ALU_N545 , ALU_N547 , ALU_N549 , ALU_N550 , ALU_N551 , ALU_N552 , ALU_N553 , 
  ALU_N554 , ALU_N556 , ALU_N558 , ALU_N559 , ALU_N560 , ALU_N561 , ALU_N562 , 
  ALU_N563 , ALU_N565 , ALU_N566 , ALU_N568 , ALU_N569 , ALU_N570 , ALU_N571 , 
  ALU_N572 , ALU_N573 , ALU_N574 , MAU_N_2809 , MAU_N229 , MAU_N228 , MAU_N231 
  , MAU_N232 , MAU_N230 , IFU_ADD_59_PLUS_PLUS_N19 , ALU_ADD_111_PLUS_N25 , 
  ALU_ADD_111_PLUS_N27 , IFU_TPC_REG_7_GSR_OR , IFU_TPC_REG_6_GSR_OR , 
  IFU_TPC_REG_5_GSR_OR , IFU_TPC_REG_4_GSR_OR , IFU_TPC_REG_3_GSR_OR , 
  IFU_TPC_REG_2_GSR_OR , IFU_TPC_REG_1_GSR_OR , IFU_TPC_REG_0_GSR_OR , 
  IDU_I_REG_6_GSR_OR , IDU_I_REG_5_GSR_OR , IDU_I_REG_4_GSR_OR , 
  IDU_I_REG_3_GSR_OR , IDU_I_REG_2_GSR_OR , IDU_I_REG_1_GSR_OR , 
  IDU_I_REG_0_GSR_OR , ALU_F_REG_1_GSR_OR , ALU_F_REG_0_GSR_OR , 
  ALU_OP2_REG_7_GSR_OR , ALU_OP2_REG_6_GSR_OR , ALU_OP2_REG_5_GSR_OR , 
  ALU_OP2_REG_4_GSR_OR , ALU_OP2_REG_3_GSR_OR , ALU_OP2_REG_2_GSR_OR , 
  ALU_OP2_REG_1_GSR_OR , ALU_OP2_REG_0_GSR_OR , ALU_I2_INT_REG_7_GSR_OR , 
  ALU_I2_INT_REG_6_GSR_OR , ALU_I2_INT_REG_5_GSR_OR , ALU_I2_INT_REG_4_GSR_OR , 
  ALU_I2_INT_REG_3_GSR_OR , ALU_I2_INT_REG_2_GSR_OR , ALU_I2_INT_REG_1_GSR_OR , 
  ALU_I2_INT_REG_0_GSR_OR , ALU_CTR_ALU_REG_10_GSR_OR , 
  ALU_CTR_ALU_REG_7_GSR_OR , MAU_ADR_OUT_REG_7_GSR_OR , 
  MAU_ADR_OUT_REG_6_GSR_OR , MAU_ADR_OUT_REG_5_GSR_OR , 
  MAU_ADR_OUT_REG_4_GSR_OR , MAU_ADR_OUT_REG_3_GSR_OR , 
  MAU_ADR_OUT_REG_2_GSR_OR , MAU_ADR_OUT_REG_1_GSR_OR , 
  MAU_ADR_OUT_REG_0_GSR_OR , MAU_CTR_MAU_REG_1_GSR_OR , 
  MAU_CTR_MAU_REG_0_GSR_OR , MAU_REG_CTR_REG_1_GSR_OR , 
  MAU_REG_CTR_REG_0_GSR_OR , STU_1_INV , ALU_U218_GATE2 , ALU_U218_O_2_0 , 
  ALU_U196_GATE1 , ALU_U196_GATE2 , ALU_U196_GATE3 , ALU_U196_O_2_0 , 
  ALU_A_IN_6_3_INV , ALU_U208_GATE2 , ALU_U208_O_2_0 , ALU_A_IN_5_1_INV , 
  ALU_U228_GATE2 , ALU_U228_O_2_0 , ALU_A_IN_4_3_INV , ALU_U187_GATE1 , 
  ALU_U187_GATE2 , ALU_U187_GATE3 , ALU_U187_O_2_0 , ALU_A_IN_3_0_INV , 
  ALU_U238_GATE2 , ALU_U238_O_2_0 , ALU_A_IN_2_3_INV , ALU_U178_GATE1 , 
  ALU_U178_GATE2 , ALU_U178_GATE3 , ALU_U178_O_2_0 , ALU_A_IN_1_1_INV , 
  ALU_U242_GATE2 , ALU_U242_GATE3 , ALU_U242_O_2_0 , ALU_A_IN_0_9_INV , 
  ALU_A_IN_0_11_INV , ALU_A_IN_0_12_INV , IDU_N71_2_INV , IDU_N71_4_INV , 
  IDU_U76_GATE1 , ALU_CTR_ALU_9_1_INV , ALU_CTR_ALU_9_4_INV , 
  ALU_CTR_ALU_9_5_INV , ALU_CTR_ALU_9_12_INV , IDU_N96 , CTR_1_0_4299 , 
  U134_1I20_GTS_TRI , U135_1I20_GTS_TRI , U136_1I20_GTS_TRI , U137_1I20_GTS_TRI 
  , U138_1I20_GTS_TRI , U139_1I20_GTS_TRI , U140_1I20_GTS_TRI , 
  U141_1I20_GTS_TRI , U158_1I20_GTS_TRI , U159_1I20_GTS_TRI , U160_1I20_GTS_TRI 
  , U161_1I20_GTS_TRI , U162_1I20_GTS_TRI , U163_1I20_GTS_TRI , 
  U164_1I20_GTS_TRI , U165_1I20_GTS_TRI , U166_1I20_GTS_TRI , U167_1I20_GTS_TRI 
  , U168_1I20_GTS_TRI , U169_1I20_GTS_TRI , U170_1I20_GTS_TRI , 
  U171_1I20_GTS_TRI , U172_1I20_GTS_TRI , U173_1I20_GTS_TRI , U174_1I20_GTS_TRI 
  , U175_1I20_GTS_TRI , U176_1I20_GTS_TRI , U177_1I20_GTS_TRI , 
  U178_1I20_GTS_TRI , U179_1I20_GTS_TRI , U180_1I20_GTS_TRI , U181_1I20_GTS_TRI 
  , U182_1I20_GTS_TRI , U183_1I20_GTS_TRI , U184_1I20_GTS_TRI , 
  U185_1I20_GTS_TRI , U186_1I20_GTS_TRI , U187_1I20_GTS_TRI , U188_1I20_GTS_TRI 
  , U189_1I20_GTS_TRI , U190_1I20_GTS_TRI , U191_1I20_GTS_TRI , 
  U192_1I20_GTS_TRI , U193_1I20_GTS_TRI , IFU_U44_GATE1 , IFU_U44_GATE2 , 
  IFU_U44_GATE1_2_0 , IFU_U44_GATE2_2_0 , IFU_U45_GATE1 , IFU_U45_GATE2 , 
  IFU_U45_GATE1_2_0 , IFU_U45_GATE2_2_0 , IFU_U46_GATE1 , IFU_U46_GATE2 , 
  IFU_U46_GATE1_2_0 , IFU_U46_GATE2_2_0 , IFU_U47_GATE1 , IFU_U47_GATE2 , 
  IFU_U47_GATE1_2_0 , IFU_U47_GATE2_2_0 , IFU_U48_GATE1 , IFU_U48_GATE2 , 
  IFU_U48_GATE1_2_0 , IFU_U48_GATE2_2_0 , IFU_U49_GATE1 , IFU_U49_GATE2 , 
  IFU_U49_GATE1_2_0 , IFU_U49_GATE2_2_0 , IFU_U50_GATE1 , IFU_U50_GATE2 , 
  IFU_U50_GATE1_2_0 , IFU_U50_GATE2_2_0 , IFU_U51_GATE1 , IFU_U51_GATE2 , 
  IFU_U51_GATE1_2_0 , IFU_U51_GATE2_2_0 , IDU_U35_GATE1 , IDU_U35_GATE2 , 
  IDU_U35_GATE1_2_0 , IDU_U35_GATE2_2_0 , PSU_U33_GATE1 , 
  PSU_STEP2_REG_1I13_GSR_OR , PSU_GO_A_REG_1I13_GSR_OR , PSU_EN_REG_1I13_GSR_OR 
  , PSU_STEP1_REG_1I13_GSR_OR , ALU_U129_GATE1 , ALU_U129_GATE2 , 
  ALU_U129_GATE1_2_0 , ALU_U129_GATE2_2_0 , ALU_U130_GATE1 , ALU_U130_GATE2 , 
  ALU_U130_GATE1_2_0 , ALU_U130_GATE2_2_0 , ALU_U131_GATE1 , ALU_U131_GATE2 , 
  ALU_U131_GATE1_2_0 , ALU_U131_GATE2_2_0 , ALU_U132_GATE1 , ALU_U132_GATE2 , 
  ALU_U132_GATE1_2_0 , ALU_U132_GATE2_2_0 , ALU_U133_GATE1 , ALU_U133_GATE2 , 
  ALU_U133_GATE1_2_0 , ALU_U133_GATE2_2_0 , ALU_U134_GATE1 , ALU_U134_GATE2 , 
  ALU_U134_GATE1_2_0 , ALU_U134_GATE2_2_0 , ALU_U135_GATE1 , ALU_U135_GATE2 , 
  ALU_U135_GATE1_2_0 , ALU_U135_GATE2_2_0 , ALU_U136_GATE1 , ALU_U136_GATE2 , 
  ALU_U136_GATE1_2_0 , ALU_U136_GATE2_2_0 , ALU_U137_GATE1 , ALU_U137_GATE2 , 
  ALU_U137_GATE1_2_0 , ALU_U137_GATE2_2_0 , ALU_U138_GATE1 , ALU_U138_GATE2 , 
  ALU_U138_GATE1_2_0 , ALU_U138_GATE2_2_0 , ALU_U156_GATE1 , ALU_U156_GATE2 , 
  ALU_U157_GATE1 , ALU_U157_GATE2 , ALU_U158_GATE1 , ALU_U158_GATE2 , 
  ALU_U158_GATE3 , ALU_U158_O_2_0 , ALU_U172_GATE1 , ALU_U172_GATE1_2_0 , 
  ALU_U173_GATE1 , ALU_U173_GATE2 , ALU_U177_GATE1 , ALU_U179_GATE1 , 
  ALU_U179_GATE2 , ALU_U180_GATE1 , ALU_U182_GATE1 , ALU_U182_GATE2 , 
  ALU_U186_GATE1 , ALU_U188_GATE1 , ALU_U188_GATE2 , ALU_U189_GATE1 , 
  ALU_U191_GATE1 , ALU_U191_GATE2 , ALU_U195_GATE1 , ALU_U197_GATE1 , 
  ALU_U197_GATE2 , ALU_U198_GATE1 , ALU_U200_GATE1 , ALU_U200_GATE2 , 
  ALU_U203_GATE1 , ALU_U204_GATE1 , ALU_U204_GATE2 , ALU_U206_GATE1 , 
  ALU_U210_GATE1 , ALU_U210_GATE2 , ALU_U211_GATE1 , ALU_U211_GATE1_2_0 , 
  ALU_U213_GATE1 , ALU_U214_GATE1 , ALU_U214_GATE2 , ALU_U216_GATE1 , 
  ALU_U220_GATE1 , ALU_U220_GATE2 , ALU_U223_GATE1 , ALU_U224_GATE1 , 
  ALU_U224_GATE2 , ALU_U226_GATE1 , ALU_U230_GATE1 , ALU_U230_GATE2 , 
  ALU_U233_GATE1 , ALU_U234_GATE1 , ALU_U234_GATE2 , ALU_U236_GATE1 , 
  ALU_U244_GATE1 , ALU_U244_GATE2 , ALU_U244_GATE1_2_0 , ALU_U246_GATE1 , 
  ALU_U246_GATE2 , ALU_U247_GATE1 , ALU_U247_GATE2 , ALU_U247_GATE1_2_0 , 
  ALU_U248_GATE1 , ALU_U248_O_2_0 , MAU_U94_GATE1 , MAU_U94_GATE2 , 
  MAU_U94_GATE3 , MAU_U94_O_2_0 , MAU_U95_GATE1 , MAU_U95_GATE2 , MAU_U95_GATE3 
  , MAU_U95_O_2_0 , MAU_NRD_REG_1I13_GSR_OR , MAU_NWR_REG_1I13_GSR_OR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_7 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_6 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_5 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_4 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_3 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_2 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_1 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C1 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C2 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C3 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C4 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C5 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C6 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C7 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_COUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_C , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C3_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXB_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_CIN_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C0 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C1 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C2 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C3 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C4 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C5 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C6 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C7 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_C , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C3_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXB_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_CIN_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ZERO , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C0 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C1 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C2 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C3 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C4 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C5 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C6 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C7 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_C , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C3_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXB_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_CIN_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ZERO , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C0 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C1 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C2 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C3 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C4 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C5 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C6 , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C7 
  , IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_C , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C3_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXB_OUT , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_CIN_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_XOR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT0_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_2_0 , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_CO_8 , ALU_ADD_111_PLUS_U10_S0_1_CO_7 , 
  ALU_ADD_111_PLUS_U10_S0_1_CO_6 , ALU_ADD_111_PLUS_U10_S0_1_CO_5 , 
  ALU_ADD_111_PLUS_U10_S0_1_CO_4 , ALU_ADD_111_PLUS_U10_S0_1_CO_3 , 
  ALU_ADD_111_PLUS_U10_S0_1_CO_2 , ALU_ADD_111_PLUS_U10_S0_1_CO_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_CO_9 , ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C0 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C1 , ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C2 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C3 , ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C4 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C5 , ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C6 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C7 , ALU_ADD_111_PLUS_U10_S0_1_CY4_5_COUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_C , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C3_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXB_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_CIN_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ZERO , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C0 , ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C1 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C2 , ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C3 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C4 , ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C5 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C6 , ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C7 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_C , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C3_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXB_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_CIN_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ZERO , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C0 , ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C1 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C2 , ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C3 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C4 , ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C5 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C6 , ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C7 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_C , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C3_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXB_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_CIN_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ZERO , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C0 , ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C1 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C2 , ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C3 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C4 , ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C5 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C6 , ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C7 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_C , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C3_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXB_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_CIN_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ZERO , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C0 , ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C1 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C2 , ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C3 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C4 , ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C5 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C6 , ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C7 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_COUT0 , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_C , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C3_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXB_OUT , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_CIN_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_XOR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT0_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ONE , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_1 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_2_0 , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_N25_1 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_G , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_COUT0 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_1N8 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A0BUF , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A1BUF , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B0BUF , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B1BUF , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR3 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR1 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND2 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND4 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV1 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR2 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV0 , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR0 , 
  U194_CLKIO_BUFSIG , IDU_U33_2_0 , IDU_U45_2_0 , IDU_U45_2_1 , IDU_U55_2_0 , 
  IDU_U56_2_0 , IDU_U58_2_0 , IDU_U68_2_0 , IDU_U70_2_0 , ALU_U162_2_0 , 
  ALU_U162_2_1 , ALU_U165_2_0 , ALU_U166_2_0 , ALU_U168_2_0 , ALU_U168_2_1 , 
  ALU_U169_2_0 , ALU_U250_2_0 , ALU_U250_2_1 , ALU_U251_4_0 , 
  ALU_U251_ALU_F_IN_1_4_0_2_0 , ALU_U251_ALU_F_IN_1_4_0_2_1 , MAU_U90_2_0 , 
  ALU_N491_F , ALU_N491_G , ALU_N491_H1 , ALU_N491_H , ALU_N491_H0 , 
  ALU_N491_FGBLOCK_1N8 , ALU_N491_FGBLOCK_1N7 , 
  ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0 , ALU_N491_HLUT_AND0 , ALU_A_IN_6_F , 
  ALU_A_IN_6_G , ALU_A_IN_6_H1 , ALU_A_IN_6_H , ALU_A_IN_6_H0 , 
  ALU_A_IN_6_FGBLOCK_1N8 , ALU_A_IN_6_FGBLOCK_1N18 , ALU_A_IN_6_FGBLOCK_1N7 , 
  ALU_A_IN_6_FGBLOCK_LUTRAM_FLUT_OR0 , ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_6_HLUT_AND0 , ALU_A_IN_5_F , 
  ALU_A_IN_5_G , ALU_A_IN_5_H1 , ALU_A_IN_5_H , ALU_A_IN_5_H0 , 
  ALU_A_IN_5_FGBLOCK_1N8 , ALU_A_IN_5_FGBLOCK_1N18 , ALU_A_IN_5_FGBLOCK_1N7 , 
  ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0 , ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_5_HLUT_AND0 , ALU_A_IN_4_F , 
  ALU_A_IN_4_G , ALU_A_IN_4_H1 , ALU_A_IN_4_H , ALU_A_IN_4_H0 , 
  ALU_A_IN_4_FGBLOCK_1N8 , ALU_A_IN_4_FGBLOCK_1N18 , ALU_A_IN_4_FGBLOCK_1N7 , 
  ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0 , ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_4_HLUT_AND0 , ALU_A_IN_3_F , 
  ALU_A_IN_3_G , ALU_A_IN_3_H1 , ALU_A_IN_3_H , ALU_A_IN_3_H0 , 
  ALU_A_IN_3_FGBLOCK_1N8 , ALU_A_IN_3_FGBLOCK_1N7 , 
  ALU_A_IN_3_FGBLOCK_LUTRAM_FLUT_OR0 , ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_3_HLUT_AND0 , ALU_A_IN_2_F , 
  ALU_A_IN_2_G , ALU_A_IN_2_H1 , ALU_A_IN_2_H , ALU_A_IN_2_H0 , 
  ALU_A_IN_2_FGBLOCK_1N8 , ALU_A_IN_2_FGBLOCK_1N18 , ALU_A_IN_2_FGBLOCK_1N7 , 
  ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0 , ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_2_HLUT_AND0 , ALU_A_IN_1_F , 
  ALU_A_IN_1_G , ALU_A_IN_1_H1 , ALU_A_IN_1_H , ALU_A_IN_1_H0 , 
  ALU_A_IN_1_FGBLOCK_1N8 , ALU_A_IN_1_FGBLOCK_1N18 , ALU_A_IN_1_FGBLOCK_1N7 , 
  ALU_A_IN_1_FGBLOCK_LUTRAM_FLUT_OR0 , ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND0 , 
  ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND1 , ALU_A_IN_1_HLUT_AND0 , ALU_A_IN_0_F , 
  ALU_A_IN_0_G , ALU_A_IN_0_H1 , ALU_A_IN_0_H , ALU_A_IN_0_H0 , 
  ALU_A_IN_0_FGBLOCK_1N8 , ALU_A_IN_0_FGBLOCK_1N18 , ALU_A_IN_0_FGBLOCK_1N7 , 
  ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0 , ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_OR1 , 
  ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0 , ALU_A_IN_0_HLUT_AND0 , IDU_N71_F , 
  IDU_N71_G , IDU_N71_H , IDU_N71_H0 , IDU_N71_FGBLOCK_1N8 , 
  IDU_N71_FGBLOCK_1N7 , IDU_N71_FGBLOCK_LUTRAM_FLUT_AND0 , 
  IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1 , IDU_N71_FGBLOCK_LUTRAM_FLUT_AND2 , 
  IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3 , IDU_N71_FGBLOCK_LUTRAM_GLUT_AND0 , 
  IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1 , IDU_N71_FGBLOCK_LUTRAM_GLUT_OR2 , 
  IDU_N71_FGBLOCK_LUTRAM_GLUT_AND3 , CTR_1_9_F , CTR_1_9_H1 , CTR_1_9_H , 
  CTR_1_9_FGBLOCK_1N18 , CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND0 , IDU_U76_O_2_0 , 
  IDU_N96_F , IDU_N96_G , IDU_N96_H1 , IDU_N96_H , IDU_N96_H0 , 
  IDU_N96_FGBLOCK_1N8 , IDU_N96_FGBLOCK_1N18 , IDU_N96_FGBLOCK_1N7 , 
  IDU_N96_FGBLOCK_LUTRAM_FLUT_AND0 , IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0 , 
  IDU_N96_HLUT_AND0 , ALU_CTR_ALU_4_F , ALU_CTR_ALU_4_H1 , ALU_CTR_ALU_4_H , 
  ALU_CTR_ALU_4_FGBLOCK_1N18 , ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0 , 
  ALU_CTR_ALU_2_F , ALU_CTR_ALU_2_G , ALU_CTR_ALU_2_FGBLOCK_1N18 , 
  ALU_CTR_ALU_2_FGBLOCK_1N7 , ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND0 , 
  ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1 , 
  ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0 , CTR_1_0_F , CTR_1_0_G , CTR_1_0_H , 
  CTR_1_0_H0 , CTR_1_0_FGBLOCK_1N8 , CTR_1_0_FGBLOCK_1N18 , CTR_1_0_FGBLOCK_1N7 
  , CTR_1_0_FGBLOCK_LUTRAM_FLUT_AND0 , CTR_1_0_FGBLOCK_LUTRAM_GLUT_AND0 , 
  IDU_N105_F , IDU_N105_G , IDU_N105_FGBLOCK_1N8 , IDU_N105_FGBLOCK_1N18 , 
  IDU_N105_FGBLOCK_1N7 , IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0 , 
  IDU_N105_FGBLOCK_LUTRAM_GLUT_AND0 , IDU_N105_FGBLOCK_LUTRAM_GLUT_AND1 , 
  IDU_N105_FGBLOCK_LUTRAM_GLUT_AND2 , CTR_1_4_F , CTR_1_4_G , CTR_1_4_H1 , 
  CTR_1_4_H , CTR_1_4_H0 , CTR_1_4_FGBLOCK_1N8 , CTR_1_4_FGBLOCK_1N18 , 
  CTR_1_4_FGBLOCK_1N7 , CTR_1_4_FGBLOCK_LUTRAM_GLUT_AND0 , CTR_1_4_HLUT_AND0 , 
  IFU_U61_2_INV , ALU_U167_2_INV , ALU_U178_GATE1_0_INV , ALU_U187_GATE1_0_INV 
  , ALU_U196_GATE1_0_INV , MAU_U94_GATE1_0_INV , MAU_U95_GATE1_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT_2_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT_2_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND_1_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND_1_INV , 
  IFU_U44_GATE1_IFU_U44_GATE1_1_INV , IFU_U45_GATE1_IFU_U45_GATE1_1_INV , 
  IFU_U46_GATE1_IFU_U46_GATE1_1_INV , IFU_U47_GATE1_IFU_U47_GATE1_1_INV , 
  IFU_U48_GATE1_IFU_U48_GATE1_1_INV , IFU_U49_GATE1_IFU_U49_GATE1_1_INV , 
  IFU_U50_GATE1_IFU_U50_GATE1_1_INV , IFU_U51_GATE1_IFU_U51_GATE1_1_INV , 
  ALU_U129_GATE1_ALU_U129_GATE1_1_INV , ALU_U130_GATE1_ALU_U130_GATE1_1_INV , 
  ALU_U131_GATE1_ALU_U131_GATE1_1_INV , ALU_U132_GATE1_ALU_U132_GATE1_1_INV , 
  ALU_U133_GATE1_ALU_U133_GATE1_1_INV , ALU_U134_GATE1_ALU_U134_GATE1_1_INV , 
  ALU_U135_GATE1_ALU_U135_GATE1_1_INV , ALU_U136_GATE1_ALU_U136_GATE1_1_INV , 
  ALU_U137_GATE1_ALU_U137_GATE1_1_INV , ALU_U138_GATE1_ALU_U138_GATE1_1_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_2_0_0_INV , 
  IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_0_0_INV , 
  ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_2_0_0_INV , 
  IDU_U58_IDU_N66_2_INV , IDU_U68_IDU_N67_2_INV , IDU_U70_IDU_N68_2_INV , 
  ALU_U251_ALU_F_IN_1_2_INV , U134_1I20_GTS_TRI_2_INV , U135_1I20_GTS_TRI_2_INV 
  , U136_1I20_GTS_TRI_2_INV , U137_1I20_GTS_TRI_2_INV , U138_1I20_GTS_TRI_2_INV 
  , U139_1I20_GTS_TRI_2_INV , U140_1I20_GTS_TRI_2_INV , U141_1I20_GTS_TRI_2_INV 
  , U158_1I20_GTS_TRI_2_INV , U159_1I20_GTS_TRI_2_INV , U160_1I20_GTS_TRI_2_INV 
  , U161_1I20_GTS_TRI_2_INV , U162_1I20_GTS_TRI_2_INV , U163_1I20_GTS_TRI_2_INV 
  , U164_1I20_GTS_TRI_2_INV , U165_1I20_GTS_TRI_2_INV , U166_1I20_GTS_TRI_2_INV 
  , U167_1I20_GTS_TRI_2_INV , U168_1I20_GTS_TRI_2_INV , U169_1I20_GTS_TRI_2_INV 
  , U170_1I20_GTS_TRI_2_INV , U171_1I20_GTS_TRI_2_INV , U172_1I20_GTS_TRI_2_INV 
  , U173_1I20_GTS_TRI_2_INV , U174_1I20_GTS_TRI_2_INV , U175_1I20_GTS_TRI_2_INV 
  , U176_1I20_GTS_TRI_2_INV , U177_1I20_GTS_TRI_2_INV , U178_1I20_GTS_TRI_2_INV 
  , U179_1I20_GTS_TRI_2_INV , U180_1I20_GTS_TRI_2_INV , U181_1I20_GTS_TRI_2_INV 
  , U182_1I20_GTS_TRI_2_INV , U183_1I20_GTS_TRI_2_INV , U184_1I20_GTS_TRI_2_INV 
  , U185_1I20_GTS_TRI_2_INV , U186_1I20_GTS_TRI_2_INV , U187_1I20_GTS_TRI_2_INV 
  , U188_1I20_GTS_TRI_2_INV , U189_1I20_GTS_TRI_2_INV , U190_1I20_GTS_TRI_2_INV 
  , U191_1I20_GTS_TRI_2_INV , U192_1I20_GTS_TRI_2_INV , U193_1I20_GTS_TRI_2_INV 
  , ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3_0_INV , 
  ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5_0_INV , 
  ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0_0_INV , ALU_N491_HLUT_AND0_0_INV , 
  ALU_A_IN_6_HLUT_AND0_0_INV , ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
  ALU_A_IN_5_HLUT_AND0_0_INV , ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
  ALU_A_IN_4_HLUT_AND0_0_INV , ALU_A_IN_3_HLUT_AND0_0_INV , 
  ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , ALU_A_IN_2_HLUT_AND0_0_INV , 
  ALU_A_IN_1_HLUT_AND0_0_INV , ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
  ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0_1_INV , 
  ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_1_INV , 
  ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_2_INV , 
  IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_0_INV , 
  IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
  IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3_1_INV , 
  IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1_0_INV , IDU_N71_HLUT_AND0_2_INV , 
  CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
  CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_2_INV , CTR_1_9_HLUT_AND0_0_INV , 
  CTR_1_9_HLUT_AND0_2_INV , IDU_N96_FGBLOCK_LUTRAM_FLUT_AND1_2_INV , 
  IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0_0_INV , 
  IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_0_INV , 
  IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_1_INV , 
  IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_2_INV , IDU_N96_HLUT_AND1_1_INV , 
  ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
  ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND1_0_INV , ALU_CTR_ALU_4_HLUT_AND0_1_INV 
  , ALU_CTR_ALU_4_HLUT_AND0_2_INV , 
  ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
  ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0_1_INV , CTR_1_0_HLUT_AND0_0_INV , 
  CTR_1_0_HLUT_AND0_1_INV , CTR_1_0_HLUT_AND0_2_INV , 
  IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
  IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_1_INV , VCC , GND , GSR , GTS : STD_LOGIC ;
  signal JUMP_ADR : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal IFU_RETURN89 : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal IFU_TPC35 : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal INS : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal IFU_N36 : STD_LOGIC_VECTOR ( 0 downto 0 );
  signal CTR_1 : STD_LOGIC_VECTOR ( 14 downto 0 );
  signal IDU_I : STD_LOGIC_VECTOR ( 6 downto 0 );
  signal ALU_CTR_ALU : STD_LOGIC_VECTOR ( 10 downto 0 );
  signal ALU_B_IN : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal ALU_ADD : STD_LOGIC_VECTOR ( 8 downto 0 );
  signal ALU_F_IN : STD_LOGIC_VECTOR ( 1 downto 0 );
  signal ADR : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal REG_CTR : STD_LOGIC_VECTOR ( 1 downto 0 );
  signal ALU_A_IN : STD_LOGIC_VECTOR ( 7 downto 0 );
  signal CTR_2 : STD_LOGIC_VECTOR ( 3 downto 0 );
  signal MAU_CTR_MAU : STD_LOGIC_VECTOR ( 1 downto 0 );
  begin
    U132 : X_ZERO 
      port map ( O => NET4 ) ;
    U142 : X_BUF 
      port map ( I => PROG_DATA(7) , O => N73 ) ;
    U143 : X_BUF 
      port map ( I => PROG_DATA(6) , O => N74 ) ;
    U144 : X_BUF 
      port map ( I => PROG_DATA(5) , O => N75 ) ;
    U145 : X_BUF 
      port map ( I => PROG_DATA(4) , O => N76 ) ;
    U146 : X_BUF 
      port map ( I => PROG_DATA(3) , O => N77 ) ;
    U147 : X_BUF 
      port map ( I => PROG_DATA(2) , O => N78 ) ;
    U148 : X_BUF 
      port map ( I => PROG_DATA(1) , O => N79 ) ;
    U149 : X_BUF 
      port map ( I => PROG_DATA(0) , O => N80 ) ;
    U150 : X_BUF 
      port map ( I => DATMEM_DATA_IN(7) , O => N81 ) ;
    U151 : X_BUF 
      port map ( I => DATMEM_DATA_IN(6) , O => N82 ) ;
    U152 : X_BUF 
      port map ( I => DATMEM_DATA_IN(5) , O => N83 ) ;
    U153 : X_BUF 
      port map ( I => DATMEM_DATA_IN(4) , O => N84 ) ;
    U154 : X_BUF 
      port map ( I => DATMEM_DATA_IN(3) , O => N85 ) ;
    U155 : X_BUF 
      port map ( I => DATMEM_DATA_IN(2) , O => N86 ) ;
    U156 : X_BUF 
      port map ( I => DATMEM_DATA_IN(1) , O => N87 ) ;
    U157 : X_BUF 
      port map ( I => DATMEM_DATA_IN(0) , O => N88 ) ;
    U195 : X_BUF 
      port map ( I => NRESET , O => N126 ) ;
    U196 : X_BUF 
      port map ( I => GO_STEP , O => N127 ) ;
    U197 : X_BUF 
      port map ( I => ONE_STEP , O => N128 ) ;
    IFU_U43 : X_ONE 
      port map ( O => IFU_N135 ) ;
    IFU_U52 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N73 , O => INS(7) ) ;
    IFU_U53 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N74 , O => INS(6) ) ;
    IFU_U54 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N75 , O => INS(5) ) ;
    IFU_U56 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N77 , O => INS(3) ) ;
    IFU_U57 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N78 , O => INS(2) ) ;
    IFU_U58 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N79 , O => INS(1) ) ;
    IFU_U59 : X_AND2 
      port map ( I0 => IFU_N136 , I1 => N80 , O => INS(0) ) ;
    IFU_U60 : X_OR2 
      port map ( I0 => JDEC , I1 => EN , O => IFU_N36(0) ) ;
    IFU_U61 : X_OR2 
      port map ( I0 => JDEC , I1 => SEC_B , O => IFU_U61_2_INV ) ;
    IFU_TPC_REG_7_Q : X_FF 
      port map ( I => IFU_TPC35(7) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_7_GSR_OR , O => N308 ) ;
    IFU_TPC_REG_6_Q : X_FF 
      port map ( I => IFU_TPC35(6) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_6_GSR_OR , O => N309 ) ;
    IFU_TPC_REG_5_Q : X_FF 
      port map ( I => IFU_TPC35(5) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_5_GSR_OR , O => N310 ) ;
    IFU_TPC_REG_4_Q : X_FF 
      port map ( I => IFU_TPC35(4) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_4_GSR_OR , O => N311 ) ;
    IFU_TPC_REG_3_Q : X_FF 
      port map ( I => IFU_TPC35(3) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_3_GSR_OR , O => N312 ) ;
    IFU_TPC_REG_2_Q : X_FF 
      port map ( I => IFU_TPC35(2) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_2_GSR_OR , O => N313 ) ;
    IFU_TPC_REG_1_Q : X_FF 
      port map ( I => IFU_TPC35(1) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_1_GSR_OR , O => N314 ) ;
    IFU_TPC_REG_0_Q : X_FF 
      port map ( I => IFU_TPC35(0) , CLK => N125 , CE => IFU_N36(0) , 
      SET => GND , RST => IFU_TPC_REG_0_GSR_OR , O => N315 ) ;
    IDU_U57 : X_AND2 
      port map ( I0 => IDU_N92 , I1 => IDU_I(0) , O => IDU_N60 ) ;
    IDU_U74 : X_INV 
      port map ( I => IDU_N60 , O => IDU_N103 ) ;
    IDU_I_REG_6_Q : X_FF 
      port map ( I => INS(7) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_6_GSR_OR , O => IDU_I(6) ) ;
    IDU_I_REG_5_Q : X_FF 
      port map ( I => INS(6) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_5_GSR_OR , O => IDU_I(5) ) ;
    IDU_I_REG_4_Q : X_FF 
      port map ( I => INS(5) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_4_GSR_OR , O => IDU_I(4) ) ;
    IDU_I_REG_3_Q : X_FF 
      port map ( I => INS(3) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_3_GSR_OR , O => IDU_I(3) ) ;
    IDU_I_REG_2_Q : X_FF 
      port map ( I => INS(2) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_2_GSR_OR , O => IDU_I(2) ) ;
    IDU_I_REG_1_Q : X_FF 
      port map ( I => INS(1) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_1_GSR_OR , O => IDU_I(1) ) ;
    IDU_I_REG_0_Q : X_FF 
      port map ( I => INS(0) , CLK => N125 , CE => EN , SET => GND , 
      RST => IDU_I_REG_0_GSR_OR , O => IDU_I(0) ) ;
    ALU_U128 : X_ONE 
      port map ( O => ALU_N474 ) ;
    ALU_U164 : X_AND2 
      port map ( I0 => ALU_N492 , I1 => ALU_N496 , O => ALU_N497 ) ;
    ALU_U167 : X_OR2 
      port map ( I0 => ALU_N495 , I1 => ALU_CTR_ALU(3) , O => ALU_U167_2_INV ) ;
    ALU_U176 : X_AND2 
      port map ( I0 => ALU_N507 , I1 => ALU_N494 , O => ALU_N508 ) ;
    ALU_U185 : X_AND2 
      port map ( I0 => ALU_N515 , I1 => ALU_N494 , O => ALU_N516 ) ;
    ALU_U194 : X_AND2 
      port map ( I0 => ALU_N523 , I1 => ALU_N494 , O => ALU_N524 ) ;
    ALU_U207 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(3) , I1 => JUMP_ADR(5) , O => ALU_N536 ) ;
    ALU_U217 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(3) , I1 => JUMP_ADR(7) , O => ALU_N545 ) ;
    ALU_U227 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(3) , I1 => JUMP_ADR(4) , O => ALU_N554 ) ;
    ALU_U237 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(3) , I1 => JUMP_ADR(2) , O => ALU_N563 ) ;
    ALU_U241 : X_AND2 
      port map ( I0 => ALU_N565 , I1 => ALU_N494 , O => ALU_N566 ) ;
    ALU_U245 : X_AND2 
      port map ( I0 => N349 , I1 => N341 , O => ALU_N570 ) ;
    ALU_F_REG_1_Q : X_FF 
      port map ( I => ALU_F_IN(1) , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_F_REG_1_GSR_OR , O => N351 ) ;
    ALU_F_REG_0_Q : X_FF 
      port map ( I => ALU_F_IN(0) , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_F_REG_0_GSR_OR , O => N350 ) ;
    ALU_OP2_REG_7_Q : X_FF 
      port map ( I => ALU_B_IN(7) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_7_GSR_OR , O => N342 ) ;
    ALU_OP2_REG_6_Q : X_FF 
      port map ( I => ALU_B_IN(6) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_6_GSR_OR , O => N343 ) ;
    ALU_OP2_REG_5_Q : X_FF 
      port map ( I => ALU_B_IN(5) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_5_GSR_OR , O => N344 ) ;
    ALU_OP2_REG_4_Q : X_FF 
      port map ( I => ALU_B_IN(4) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_4_GSR_OR , O => N345 ) ;
    ALU_OP2_REG_3_Q : X_FF 
      port map ( I => ALU_B_IN(3) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_3_GSR_OR , O => N346 ) ;
    ALU_OP2_REG_2_Q : X_FF 
      port map ( I => ALU_B_IN(2) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_2_GSR_OR , O => N347 ) ;
    ALU_OP2_REG_1_Q : X_FF 
      port map ( I => ALU_B_IN(1) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_1_GSR_OR , O => N348 ) ;
    ALU_OP2_REG_0_Q : X_FF 
      port map ( I => ALU_B_IN(0) , CLK => N125 , CE => ALU_N_2432 , SET => GND 
      , RST => ALU_OP2_REG_0_GSR_OR , O => N349 ) ;
    ALU_I2_INT_REG_7_Q : X_FF 
      port map ( I => N73 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_7_GSR_OR , O => JUMP_ADR(7) ) ;
    ALU_I2_INT_REG_6_Q : X_FF 
      port map ( I => N74 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_6_GSR_OR , O => JUMP_ADR(6) ) ;
    ALU_I2_INT_REG_5_Q : X_FF 
      port map ( I => N75 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_5_GSR_OR , O => JUMP_ADR(5) ) ;
    ALU_I2_INT_REG_4_Q : X_FF 
      port map ( I => N76 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_4_GSR_OR , O => JUMP_ADR(4) ) ;
    ALU_I2_INT_REG_3_Q : X_FF 
      port map ( I => N77 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_3_GSR_OR , O => JUMP_ADR(3) ) ;
    ALU_I2_INT_REG_2_Q : X_FF 
      port map ( I => N78 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_2_GSR_OR , O => JUMP_ADR(2) ) ;
    ALU_I2_INT_REG_1_Q : X_FF 
      port map ( I => N79 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_1_GSR_OR , O => JUMP_ADR(1) ) ;
    ALU_I2_INT_REG_0_Q : X_FF 
      port map ( I => N80 , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_I2_INT_REG_0_GSR_OR , O => JUMP_ADR(0) ) ;
    ALU_CTR_ALU_REG_10_Q : X_FF 
      port map ( I => CTR_1(14) , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_CTR_ALU_REG_10_GSR_OR , O => ALU_CTR_ALU(10) ) ;
    ALU_CTR_ALU_REG_7_Q : X_FF 
      port map ( I => CTR_1(11) , CLK => N125 , CE => EN , SET => GND , 
      RST => ALU_CTR_ALU_REG_7_GSR_OR , O => ALU_CTR_ALU(7) ) ;
    MAU_ADR_OUT_REG_7_Q : X_FF 
      port map ( I => ADR(7) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_7_GSR_OR , O => N326 ) ;
    MAU_ADR_OUT_REG_6_Q : X_FF 
      port map ( I => ADR(6) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_6_GSR_OR , O => N327 ) ;
    MAU_ADR_OUT_REG_5_Q : X_FF 
      port map ( I => ADR(5) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_5_GSR_OR , O => N328 ) ;
    MAU_ADR_OUT_REG_4_Q : X_FF 
      port map ( I => ADR(4) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_4_GSR_OR , O => N329 ) ;
    MAU_ADR_OUT_REG_3_Q : X_FF 
      port map ( I => ADR(3) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_3_GSR_OR , O => N330 ) ;
    MAU_ADR_OUT_REG_2_Q : X_FF 
      port map ( I => ADR(2) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_2_GSR_OR , O => N331 ) ;
    MAU_ADR_OUT_REG_1_Q : X_FF 
      port map ( I => ADR(1) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_1_GSR_OR , O => N332 ) ;
    MAU_ADR_OUT_REG_0_Q : X_FF 
      port map ( I => ADR(0) , CLK => N125 , CE => MAU_N_2809 , SET => GND , 
      RST => MAU_ADR_OUT_REG_0_GSR_OR , O => N333 ) ;
    MAU_CTR_MAU_REG_1_Q : X_FF 
      port map ( I => CTR_2(3) , CLK => N125 , CE => EN , SET => GND , 
      RST => MAU_CTR_MAU_REG_1_GSR_OR , O => MAU_CTR_MAU(1) ) ;
    MAU_CTR_MAU_REG_0_Q : X_FF 
      port map ( I => CTR_2(2) , CLK => N125 , CE => EN , SET => GND , 
      RST => MAU_CTR_MAU_REG_0_GSR_OR , O => MAU_CTR_MAU(0) ) ;
    MAU_REG_CTR_REG_1_Q : X_FF 
      port map ( I => CTR_2(1) , CLK => N125 , CE => EN , SET => GND , 
      RST => MAU_REG_CTR_REG_1_GSR_OR , O => REG_CTR(1) ) ;
    MAU_REG_CTR_REG_0_Q : X_FF 
      port map ( I => CTR_2(0) , CLK => N125 , CE => EN , SET => GND , 
      RST => MAU_REG_CTR_REG_0_GSR_OR , O => REG_CTR(0) ) ;
    IFU_ADD_59_PLUS_PLUS_U6 : X_ONE 
      port map ( O => IFU_ADD_59_PLUS_PLUS_N19 ) ;
    ALU_ADD_111_PLUS_U6 : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_N27 ) ;
    ALU_ADD_111_PLUS_U7 : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_N25 ) ;
    IFU_TPC_REG_7_GSR_OR_1394 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_7_GSR_OR ) ;
    IFU_TPC_REG_6_GSR_OR_1395 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_6_GSR_OR ) ;
    IFU_TPC_REG_5_GSR_OR_1396 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_5_GSR_OR ) ;
    IFU_TPC_REG_4_GSR_OR_1397 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_4_GSR_OR ) ;
    IFU_TPC_REG_3_GSR_OR_1398 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_3_GSR_OR ) ;
    IFU_TPC_REG_2_GSR_OR_1399 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_2_GSR_OR ) ;
    IFU_TPC_REG_1_GSR_OR_1400 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_1_GSR_OR ) ;
    IFU_TPC_REG_0_GSR_OR_1401 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IFU_TPC_REG_0_GSR_OR ) ;
    IDU_I_REG_6_GSR_OR_1402 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_6_GSR_OR ) ;
    IDU_I_REG_5_GSR_OR_1403 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_5_GSR_OR ) ;
    IDU_I_REG_4_GSR_OR_1404 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_4_GSR_OR ) ;
    IDU_I_REG_3_GSR_OR_1405 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_3_GSR_OR ) ;
    IDU_I_REG_2_GSR_OR_1406 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_2_GSR_OR ) ;
    IDU_I_REG_1_GSR_OR_1407 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_1_GSR_OR ) ;
    IDU_I_REG_0_GSR_OR_1408 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => IDU_I_REG_0_GSR_OR ) ;
    ALU_F_REG_1_GSR_OR_1417 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_F_REG_1_GSR_OR ) ;
    ALU_F_REG_0_GSR_OR_1418 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_F_REG_0_GSR_OR ) ;
    ALU_OP2_REG_7_GSR_OR_1419 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_7_GSR_OR ) ;
    ALU_OP2_REG_6_GSR_OR_1420 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_6_GSR_OR ) ;
    ALU_OP2_REG_5_GSR_OR_1421 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_5_GSR_OR ) ;
    ALU_OP2_REG_4_GSR_OR_1422 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_4_GSR_OR ) ;
    ALU_OP2_REG_3_GSR_OR_1423 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_3_GSR_OR ) ;
    ALU_OP2_REG_2_GSR_OR_1424 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_2_GSR_OR ) ;
    ALU_OP2_REG_1_GSR_OR_1425 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_1_GSR_OR ) ;
    ALU_OP2_REG_0_GSR_OR_1426 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_OP2_REG_0_GSR_OR ) ;
    ALU_I2_INT_REG_7_GSR_OR_1427 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_7_GSR_OR ) ;
    ALU_I2_INT_REG_6_GSR_OR_1428 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_6_GSR_OR ) ;
    ALU_I2_INT_REG_5_GSR_OR_1429 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_5_GSR_OR ) ;
    ALU_I2_INT_REG_4_GSR_OR_1430 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_4_GSR_OR ) ;
    ALU_I2_INT_REG_3_GSR_OR_1431 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_3_GSR_OR ) ;
    ALU_I2_INT_REG_2_GSR_OR_1432 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_2_GSR_OR ) ;
    ALU_I2_INT_REG_1_GSR_OR_1433 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_1_GSR_OR ) ;
    ALU_I2_INT_REG_0_GSR_OR_1434 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_I2_INT_REG_0_GSR_OR ) ;
    ALU_CTR_ALU_REG_10_GSR_OR_1435 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_CTR_ALU_REG_10_GSR_OR ) ;
    ALU_CTR_ALU_REG_7_GSR_OR_1438 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => ALU_CTR_ALU_REG_7_GSR_OR ) ;
    MAU_ADR_OUT_REG_7_GSR_OR_1450 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_7_GSR_OR ) ;
    MAU_ADR_OUT_REG_6_GSR_OR_1451 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_6_GSR_OR ) ;
    MAU_ADR_OUT_REG_5_GSR_OR_1452 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_5_GSR_OR ) ;
    MAU_ADR_OUT_REG_4_GSR_OR_1453 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_4_GSR_OR ) ;
    MAU_ADR_OUT_REG_3_GSR_OR_1454 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_3_GSR_OR ) ;
    MAU_ADR_OUT_REG_2_GSR_OR_1455 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_2_GSR_OR ) ;
    MAU_ADR_OUT_REG_1_GSR_OR_1456 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_1_GSR_OR ) ;
    MAU_ADR_OUT_REG_0_GSR_OR_1457 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_ADR_OUT_REG_0_GSR_OR ) ;
    MAU_CTR_MAU_REG_1_GSR_OR_1458 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_CTR_MAU_REG_1_GSR_OR ) ;
    MAU_CTR_MAU_REG_0_GSR_OR_1459 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_CTR_MAU_REG_0_GSR_OR ) ;
    MAU_REG_CTR_REG_1_GSR_OR_1460 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_REG_CTR_REG_1_GSR_OR ) ;
    MAU_REG_CTR_REG_0_GSR_OR_1461 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_REG_CTR_REG_0_GSR_OR ) ;
    STU_1_INV_1509 : X_INV 
      port map ( I => RST , O => STU_1_INV ) ;
    ALU_U218_GATE2_607 : X_AND2 
      port map ( I0 => N334 , I1 => ALU_N544 , O => ALU_U218_GATE2 ) ;
    ALU_U218_O_ALU_N546_2_0 : X_OR2 
      port map ( I0 => ALU_N545 , I1 => ALU_U218_GATE2 , O => ALU_U218_O_2_0 ) ;
    ALU_U196_GATE1_562 : X_AND2 
      port map ( I0 => ALU_U196_GATE1_0_INV , I1 => ALU_N525 , 
      O => ALU_U196_GATE1 ) ;
    ALU_U196_GATE2_563 : X_AND2 
      port map ( I0 => ALU_N524 , I1 => N335 , O => ALU_U196_GATE2 ) ;
    ALU_U196_GATE3_564 : X_AND2 
      port map ( I0 => ALU_N502 , I1 => N335 , O => ALU_U196_GATE3 ) ;
    ALU_U196_O_ALU_N526_2_0 : X_OR2 
      port map ( I0 => ALU_U196_GATE3 , I1 => ALU_U196_GATE2 , 
      O => ALU_U196_O_2_0 ) ;
    ALU_A_IN_6_3_INV_1572 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_6_3_INV ) ;
    ALU_U208_GATE2_588 : X_AND2 
      port map ( I0 => N336 , I1 => ALU_N535 , O => ALU_U208_GATE2 ) ;
    ALU_U208_O_ALU_N537_2_0 : X_OR2 
      port map ( I0 => ALU_N536 , I1 => ALU_U208_GATE2 , O => ALU_U208_O_2_0 ) ;
    ALU_A_IN_5_1_INV_1593 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_5_1_INV ) ;
    ALU_U228_GATE2_626 : X_AND2 
      port map ( I0 => N337 , I1 => ALU_N553 , O => ALU_U228_GATE2 ) ;
    ALU_U228_O_ALU_N555_2_0 : X_OR2 
      port map ( I0 => ALU_N554 , I1 => ALU_U228_GATE2 , O => ALU_U228_O_2_0 ) ;
    ALU_A_IN_4_3_INV_1614 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_4_3_INV ) ;
    ALU_U187_GATE1_543 : X_AND2 
      port map ( I0 => ALU_U187_GATE1_0_INV , I1 => ALU_N517 , 
      O => ALU_U187_GATE1 ) ;
    ALU_U187_GATE2_544 : X_AND2 
      port map ( I0 => ALU_N516 , I1 => N338 , O => ALU_U187_GATE2 ) ;
    ALU_U187_GATE3_545 : X_AND2 
      port map ( I0 => ALU_N502 , I1 => N338 , O => ALU_U187_GATE3 ) ;
    ALU_U187_O_ALU_N518_2_0 : X_OR2 
      port map ( I0 => ALU_U187_GATE3 , I1 => ALU_U187_GATE2 , 
      O => ALU_U187_O_2_0 ) ;
    ALU_A_IN_3_0_INV_1634 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_3_0_INV ) ;
    ALU_U238_GATE2_645 : X_AND2 
      port map ( I0 => N339 , I1 => ALU_N562 , O => ALU_U238_GATE2 ) ;
    ALU_U238_O_ALU_N564_2_0 : X_OR2 
      port map ( I0 => ALU_N563 , I1 => ALU_U238_GATE2 , O => ALU_U238_O_2_0 ) ;
    ALU_A_IN_2_3_INV_1655 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_2_3_INV ) ;
    ALU_U178_GATE1_524 : X_AND2 
      port map ( I0 => ALU_U178_GATE1_0_INV , I1 => ALU_N509 , 
      O => ALU_U178_GATE1 ) ;
    ALU_U178_GATE2_525 : X_AND2 
      port map ( I0 => ALU_N508 , I1 => N340 , O => ALU_U178_GATE2 ) ;
    ALU_U178_GATE3_526 : X_AND2 
      port map ( I0 => ALU_N502 , I1 => N340 , O => ALU_U178_GATE3 ) ;
    ALU_U178_O_ALU_N510_2_0 : X_OR2 
      port map ( I0 => ALU_U178_GATE3 , I1 => ALU_U178_GATE2 , 
      O => ALU_U178_O_2_0 ) ;
    ALU_A_IN_1_1_INV_1676 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_1_1_INV ) ;
    ALU_U242_GATE2_651 : X_AND2 
      port map ( I0 => ALU_N502 , I1 => N341 , O => ALU_U242_GATE2 ) ;
    ALU_U242_GATE3_652 : X_AND2 
      port map ( I0 => ALU_N566 , I1 => N341 , O => ALU_U242_GATE3 ) ;
    ALU_U242_O_ALU_N567_2_0 : X_OR2 
      port map ( I0 => ALU_U242_GATE3 , I1 => ALU_U242_GATE2 , 
      O => ALU_U242_O_2_0 ) ;
    ALU_A_IN_0_9_INV_1698 : X_INV 
      port map ( I => ALU_N495 , O => ALU_A_IN_0_9_INV ) ;
    ALU_A_IN_0_11_INV_1699 : X_INV 
      port map ( I => ALU_N496 , O => ALU_A_IN_0_11_INV ) ;
    ALU_A_IN_0_12_INV_1700 : X_INV 
      port map ( I => ALU_N493 , O => ALU_A_IN_0_12_INV ) ;
    IDU_N71_2_INV_1737 : X_INV 
      port map ( I => IDU_N103 , O => IDU_N71_2_INV ) ;
    IDU_N71_4_INV_1738 : X_INV 
      port map ( I => IDU_N92 , O => IDU_N71_4_INV ) ;
    ALU_CTR_ALU_9_1_INV_1840 : X_INV 
      port map ( I => IDU_N97 , O => ALU_CTR_ALU_9_1_INV ) ;
    ALU_CTR_ALU_9_4_INV_1841 : X_INV 
      port map ( I => IDU_N64 , O => ALU_CTR_ALU_9_4_INV ) ;
    ALU_CTR_ALU_9_5_INV_1842 : X_INV 
      port map ( I => IDU_N104 , O => ALU_CTR_ALU_9_5_INV ) ;
    ALU_CTR_ALU_9_12_INV_1843 : X_INV 
      port map ( I => IDU_N65 , O => ALU_CTR_ALU_9_12_INV ) ;
    U133_O : X_INV 
      port map ( I => N126 , O => RST ) ;
    U134_1I20 : X_BUF 
      port map ( I => N308 , O => U134_1I20_GTS_TRI ) ;
    U134_1I20_GTS_TRI_1462 : X_TRI 
      port map ( I => U134_1I20_GTS_TRI , O => PROG_ADR(7) , 
      CTL => U134_1I20_GTS_TRI_2_INV ) ;
    U135_1I20 : X_BUF 
      port map ( I => N309 , O => U135_1I20_GTS_TRI ) ;
    U135_1I20_GTS_TRI_1463 : X_TRI 
      port map ( I => U135_1I20_GTS_TRI , O => PROG_ADR(6) , 
      CTL => U135_1I20_GTS_TRI_2_INV ) ;
    U136_1I20 : X_BUF 
      port map ( I => N310 , O => U136_1I20_GTS_TRI ) ;
    U136_1I20_GTS_TRI_1464 : X_TRI 
      port map ( I => U136_1I20_GTS_TRI , O => PROG_ADR(5) , 
      CTL => U136_1I20_GTS_TRI_2_INV ) ;
    U137_1I20 : X_BUF 
      port map ( I => N311 , O => U137_1I20_GTS_TRI ) ;
    U137_1I20_GTS_TRI_1465 : X_TRI 
      port map ( I => U137_1I20_GTS_TRI , O => PROG_ADR(4) , 
      CTL => U137_1I20_GTS_TRI_2_INV ) ;
    U138_1I20 : X_BUF 
      port map ( I => N312 , O => U138_1I20_GTS_TRI ) ;
    U138_1I20_GTS_TRI_1466 : X_TRI 
      port map ( I => U138_1I20_GTS_TRI , O => PROG_ADR(3) , 
      CTL => U138_1I20_GTS_TRI_2_INV ) ;
    U139_1I20 : X_BUF 
      port map ( I => N313 , O => U139_1I20_GTS_TRI ) ;
    U139_1I20_GTS_TRI_1467 : X_TRI 
      port map ( I => U139_1I20_GTS_TRI , O => PROG_ADR(2) , 
      CTL => U139_1I20_GTS_TRI_2_INV ) ;
    U140_1I20 : X_BUF 
      port map ( I => N314 , O => U140_1I20_GTS_TRI ) ;
    U140_1I20_GTS_TRI_1468 : X_TRI 
      port map ( I => U140_1I20_GTS_TRI , O => PROG_ADR(1) , 
      CTL => U140_1I20_GTS_TRI_2_INV ) ;
    U141_1I20 : X_BUF 
      port map ( I => N315 , O => U141_1I20_GTS_TRI ) ;
    U141_1I20_GTS_TRI_1469 : X_TRI 
      port map ( I => U141_1I20_GTS_TRI , O => PROG_ADR(0) , 
      CTL => U141_1I20_GTS_TRI_2_INV ) ;
    U158_1I20 : X_BUF 
      port map ( I => N316 , O => U158_1I20_GTS_TRI ) ;
    U158_1I20_GTS_TRI_1470 : X_TRI 
      port map ( I => U158_1I20_GTS_TRI , O => DATMEM_DATA_OUT(7) , 
      CTL => U158_1I20_GTS_TRI_2_INV ) ;
    U159_1I20 : X_BUF 
      port map ( I => N317 , O => U159_1I20_GTS_TRI ) ;
    U159_1I20_GTS_TRI_1471 : X_TRI 
      port map ( I => U159_1I20_GTS_TRI , O => DATMEM_DATA_OUT(6) , 
      CTL => U159_1I20_GTS_TRI_2_INV ) ;
    U160_1I20 : X_BUF 
      port map ( I => N318 , O => U160_1I20_GTS_TRI ) ;
    U160_1I20_GTS_TRI_1472 : X_TRI 
      port map ( I => U160_1I20_GTS_TRI , O => DATMEM_DATA_OUT(5) , 
      CTL => U160_1I20_GTS_TRI_2_INV ) ;
    U161_1I20 : X_BUF 
      port map ( I => N319 , O => U161_1I20_GTS_TRI ) ;
    U161_1I20_GTS_TRI_1473 : X_TRI 
      port map ( I => U161_1I20_GTS_TRI , O => DATMEM_DATA_OUT(4) , 
      CTL => U161_1I20_GTS_TRI_2_INV ) ;
    U162_1I20 : X_BUF 
      port map ( I => N320 , O => U162_1I20_GTS_TRI ) ;
    U162_1I20_GTS_TRI_1474 : X_TRI 
      port map ( I => U162_1I20_GTS_TRI , O => DATMEM_DATA_OUT(3) , 
      CTL => U162_1I20_GTS_TRI_2_INV ) ;
    U163_1I20 : X_BUF 
      port map ( I => N321 , O => U163_1I20_GTS_TRI ) ;
    U163_1I20_GTS_TRI_1475 : X_TRI 
      port map ( I => U163_1I20_GTS_TRI , O => DATMEM_DATA_OUT(2) , 
      CTL => U163_1I20_GTS_TRI_2_INV ) ;
    U164_1I20 : X_BUF 
      port map ( I => N322 , O => U164_1I20_GTS_TRI ) ;
    U164_1I20_GTS_TRI_1476 : X_TRI 
      port map ( I => U164_1I20_GTS_TRI , O => DATMEM_DATA_OUT(1) , 
      CTL => U164_1I20_GTS_TRI_2_INV ) ;
    U165_1I20 : X_BUF 
      port map ( I => N323 , O => U165_1I20_GTS_TRI ) ;
    U165_1I20_GTS_TRI_1477 : X_TRI 
      port map ( I => U165_1I20_GTS_TRI , O => DATMEM_DATA_OUT(0) , 
      CTL => U165_1I20_GTS_TRI_2_INV ) ;
    U166_1I20 : X_BUF 
      port map ( I => N324 , O => U166_1I20_GTS_TRI ) ;
    U166_1I20_GTS_TRI_1478 : X_TRI 
      port map ( I => U166_1I20_GTS_TRI , O => DATMEM_NRD , 
      CTL => U166_1I20_GTS_TRI_2_INV ) ;
    U167_1I20 : X_BUF 
      port map ( I => N325 , O => U167_1I20_GTS_TRI ) ;
    U167_1I20_GTS_TRI_1479 : X_TRI 
      port map ( I => U167_1I20_GTS_TRI , O => DATMEM_NWR , 
      CTL => U167_1I20_GTS_TRI_2_INV ) ;
    U168_1I20 : X_BUF 
      port map ( I => N326 , O => U168_1I20_GTS_TRI ) ;
    U168_1I20_GTS_TRI_1480 : X_TRI 
      port map ( I => U168_1I20_GTS_TRI , O => DATMEM_ADR(7) , 
      CTL => U168_1I20_GTS_TRI_2_INV ) ;
    U169_1I20 : X_BUF 
      port map ( I => N327 , O => U169_1I20_GTS_TRI ) ;
    U169_1I20_GTS_TRI_1481 : X_TRI 
      port map ( I => U169_1I20_GTS_TRI , O => DATMEM_ADR(6) , 
      CTL => U169_1I20_GTS_TRI_2_INV ) ;
    U170_1I20 : X_BUF 
      port map ( I => N328 , O => U170_1I20_GTS_TRI ) ;
    U170_1I20_GTS_TRI_1482 : X_TRI 
      port map ( I => U170_1I20_GTS_TRI , O => DATMEM_ADR(5) , 
      CTL => U170_1I20_GTS_TRI_2_INV ) ;
    U171_1I20 : X_BUF 
      port map ( I => N329 , O => U171_1I20_GTS_TRI ) ;
    U171_1I20_GTS_TRI_1483 : X_TRI 
      port map ( I => U171_1I20_GTS_TRI , O => DATMEM_ADR(4) , 
      CTL => U171_1I20_GTS_TRI_2_INV ) ;
    U172_1I20 : X_BUF 
      port map ( I => N330 , O => U172_1I20_GTS_TRI ) ;
    U172_1I20_GTS_TRI_1484 : X_TRI 
      port map ( I => U172_1I20_GTS_TRI , O => DATMEM_ADR(3) , 
      CTL => U172_1I20_GTS_TRI_2_INV ) ;
    U173_1I20 : X_BUF 
      port map ( I => N331 , O => U173_1I20_GTS_TRI ) ;
    U173_1I20_GTS_TRI_1485 : X_TRI 
      port map ( I => U173_1I20_GTS_TRI , O => DATMEM_ADR(2) , 
      CTL => U173_1I20_GTS_TRI_2_INV ) ;
    U174_1I20 : X_BUF 
      port map ( I => N332 , O => U174_1I20_GTS_TRI ) ;
    U174_1I20_GTS_TRI_1486 : X_TRI 
      port map ( I => U174_1I20_GTS_TRI , O => DATMEM_ADR(1) , 
      CTL => U174_1I20_GTS_TRI_2_INV ) ;
    U175_1I20 : X_BUF 
      port map ( I => N333 , O => U175_1I20_GTS_TRI ) ;
    U175_1I20_GTS_TRI_1487 : X_TRI 
      port map ( I => U175_1I20_GTS_TRI , O => DATMEM_ADR(0) , 
      CTL => U175_1I20_GTS_TRI_2_INV ) ;
    U176_1I20 : X_BUF 
      port map ( I => N334 , O => U176_1I20_GTS_TRI ) ;
    U176_1I20_GTS_TRI_1488 : X_TRI 
      port map ( I => U176_1I20_GTS_TRI , O => A(7) , 
      CTL => U176_1I20_GTS_TRI_2_INV ) ;
    U177_1I20 : X_BUF 
      port map ( I => N335 , O => U177_1I20_GTS_TRI ) ;
    U177_1I20_GTS_TRI_1489 : X_TRI 
      port map ( I => U177_1I20_GTS_TRI , O => A(6) , 
      CTL => U177_1I20_GTS_TRI_2_INV ) ;
    U178_1I20 : X_BUF 
      port map ( I => N336 , O => U178_1I20_GTS_TRI ) ;
    U178_1I20_GTS_TRI_1490 : X_TRI 
      port map ( I => U178_1I20_GTS_TRI , O => A(5) , 
      CTL => U178_1I20_GTS_TRI_2_INV ) ;
    U179_1I20 : X_BUF 
      port map ( I => N337 , O => U179_1I20_GTS_TRI ) ;
    U179_1I20_GTS_TRI_1491 : X_TRI 
      port map ( I => U179_1I20_GTS_TRI , O => A(4) , 
      CTL => U179_1I20_GTS_TRI_2_INV ) ;
    U180_1I20 : X_BUF 
      port map ( I => N338 , O => U180_1I20_GTS_TRI ) ;
    U180_1I20_GTS_TRI_1492 : X_TRI 
      port map ( I => U180_1I20_GTS_TRI , O => A(3) , 
      CTL => U180_1I20_GTS_TRI_2_INV ) ;
    U181_1I20 : X_BUF 
      port map ( I => N339 , O => U181_1I20_GTS_TRI ) ;
    U181_1I20_GTS_TRI_1493 : X_TRI 
      port map ( I => U181_1I20_GTS_TRI , O => A(2) , 
      CTL => U181_1I20_GTS_TRI_2_INV ) ;
    U182_1I20 : X_BUF 
      port map ( I => N340 , O => U182_1I20_GTS_TRI ) ;
    U182_1I20_GTS_TRI_1494 : X_TRI 
      port map ( I => U182_1I20_GTS_TRI , O => A(1) , 
      CTL => U182_1I20_GTS_TRI_2_INV ) ;
    U183_1I20 : X_BUF 
      port map ( I => N341 , O => U183_1I20_GTS_TRI ) ;
    U183_1I20_GTS_TRI_1495 : X_TRI 
      port map ( I => U183_1I20_GTS_TRI , O => A(0) , 
      CTL => U183_1I20_GTS_TRI_2_INV ) ;
    U184_1I20 : X_BUF 
      port map ( I => N342 , O => U184_1I20_GTS_TRI ) ;
    U184_1I20_GTS_TRI_1496 : X_TRI 
      port map ( I => U184_1I20_GTS_TRI , O => B(7) , 
      CTL => U184_1I20_GTS_TRI_2_INV ) ;
    U185_1I20 : X_BUF 
      port map ( I => N343 , O => U185_1I20_GTS_TRI ) ;
    U185_1I20_GTS_TRI_1497 : X_TRI 
      port map ( I => U185_1I20_GTS_TRI , O => B(6) , 
      CTL => U185_1I20_GTS_TRI_2_INV ) ;
    U186_1I20 : X_BUF 
      port map ( I => N344 , O => U186_1I20_GTS_TRI ) ;
    U186_1I20_GTS_TRI_1498 : X_TRI 
      port map ( I => U186_1I20_GTS_TRI , O => B(5) , 
      CTL => U186_1I20_GTS_TRI_2_INV ) ;
    U187_1I20 : X_BUF 
      port map ( I => N345 , O => U187_1I20_GTS_TRI ) ;
    U187_1I20_GTS_TRI_1499 : X_TRI 
      port map ( I => U187_1I20_GTS_TRI , O => B(4) , 
      CTL => U187_1I20_GTS_TRI_2_INV ) ;
    U188_1I20 : X_BUF 
      port map ( I => N346 , O => U188_1I20_GTS_TRI ) ;
    U188_1I20_GTS_TRI_1500 : X_TRI 
      port map ( I => U188_1I20_GTS_TRI , O => B(3) , 
      CTL => U188_1I20_GTS_TRI_2_INV ) ;
    U189_1I20 : X_BUF 
      port map ( I => N347 , O => U189_1I20_GTS_TRI ) ;
    U189_1I20_GTS_TRI_1501 : X_TRI 
      port map ( I => U189_1I20_GTS_TRI , O => B(2) , 
      CTL => U189_1I20_GTS_TRI_2_INV ) ;
    U190_1I20 : X_BUF 
      port map ( I => N348 , O => U190_1I20_GTS_TRI ) ;
    U190_1I20_GTS_TRI_1502 : X_TRI 
      port map ( I => U190_1I20_GTS_TRI , O => B(1) , 
      CTL => U190_1I20_GTS_TRI_2_INV ) ;
    U191_1I20 : X_BUF 
      port map ( I => N349 , O => U191_1I20_GTS_TRI ) ;
    U191_1I20_GTS_TRI_1503 : X_TRI 
      port map ( I => U191_1I20_GTS_TRI , O => B(0) , 
      CTL => U191_1I20_GTS_TRI_2_INV ) ;
    U192_1I20 : X_BUF 
      port map ( I => N350 , O => U192_1I20_GTS_TRI ) ;
    U192_1I20_GTS_TRI_1504 : X_TRI 
      port map ( I => U192_1I20_GTS_TRI , O => CFLAG , 
      CTL => U192_1I20_GTS_TRI_2_INV ) ;
    U193_1I20 : X_BUF 
      port map ( I => N351 , O => U193_1I20_GTS_TRI ) ;
    U193_1I20_GTS_TRI_1505 : X_TRI 
      port map ( I => U193_1I20_GTS_TRI , O => ZFLAG , 
      CTL => U193_1I20_GTS_TRI_2_INV ) ;
    IFU_U44_O : X_OR2 
      port map ( I0 => IFU_U44_GATE1 , I1 => IFU_U44_GATE2 , O => IFU_TPC35(7) 
      ) ;
    IFU_U44_GATE1_IFU_U44_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(7) , 
      O => IFU_U44_GATE1_2_0 ) ;
    IFU_U44_GATE1_IFU_U44_GATE1 : X_AND2 
      port map ( I0 => IFU_U44_GATE1_2_0 , 
      I1 => IFU_U44_GATE1_IFU_U44_GATE1_1_INV , O => IFU_U44_GATE1 ) ;
    IFU_U44_GATE2_IFU_U44_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(7) , O => IFU_U44_GATE2_2_0 ) ;
    IFU_U44_GATE2_IFU_U44_GATE2 : X_AND2 
      port map ( I0 => IFU_U44_GATE2_2_0 , I1 => JDEC , O => IFU_U44_GATE2 ) ;
    IFU_U45_O : X_OR2 
      port map ( I0 => IFU_U45_GATE1 , I1 => IFU_U45_GATE2 , O => IFU_TPC35(6) 
      ) ;
    IFU_U45_GATE1_IFU_U45_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(6) , 
      O => IFU_U45_GATE1_2_0 ) ;
    IFU_U45_GATE1_IFU_U45_GATE1 : X_AND2 
      port map ( I0 => IFU_U45_GATE1_2_0 , 
      I1 => IFU_U45_GATE1_IFU_U45_GATE1_1_INV , O => IFU_U45_GATE1 ) ;
    IFU_U45_GATE2_IFU_U45_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(6) , O => IFU_U45_GATE2_2_0 ) ;
    IFU_U45_GATE2_IFU_U45_GATE2 : X_AND2 
      port map ( I0 => IFU_U45_GATE2_2_0 , I1 => JDEC , O => IFU_U45_GATE2 ) ;
    IFU_U46_O : X_OR2 
      port map ( I0 => IFU_U46_GATE1 , I1 => IFU_U46_GATE2 , O => IFU_TPC35(5) 
      ) ;
    IFU_U46_GATE1_IFU_U46_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(5) , 
      O => IFU_U46_GATE1_2_0 ) ;
    IFU_U46_GATE1_IFU_U46_GATE1 : X_AND2 
      port map ( I0 => IFU_U46_GATE1_2_0 , 
      I1 => IFU_U46_GATE1_IFU_U46_GATE1_1_INV , O => IFU_U46_GATE1 ) ;
    IFU_U46_GATE2_IFU_U46_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(5) , O => IFU_U46_GATE2_2_0 ) ;
    IFU_U46_GATE2_IFU_U46_GATE2 : X_AND2 
      port map ( I0 => IFU_U46_GATE2_2_0 , I1 => JDEC , O => IFU_U46_GATE2 ) ;
    IFU_U47_O : X_OR2 
      port map ( I0 => IFU_U47_GATE1 , I1 => IFU_U47_GATE2 , O => IFU_TPC35(4) 
      ) ;
    IFU_U47_GATE1_IFU_U47_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(4) , 
      O => IFU_U47_GATE1_2_0 ) ;
    IFU_U47_GATE1_IFU_U47_GATE1 : X_AND2 
      port map ( I0 => IFU_U47_GATE1_2_0 , 
      I1 => IFU_U47_GATE1_IFU_U47_GATE1_1_INV , O => IFU_U47_GATE1 ) ;
    IFU_U47_GATE2_IFU_U47_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(4) , O => IFU_U47_GATE2_2_0 ) ;
    IFU_U47_GATE2_IFU_U47_GATE2 : X_AND2 
      port map ( I0 => IFU_U47_GATE2_2_0 , I1 => JDEC , O => IFU_U47_GATE2 ) ;
    IFU_U48_O : X_OR2 
      port map ( I0 => IFU_U48_GATE1 , I1 => IFU_U48_GATE2 , O => IFU_TPC35(3) 
      ) ;
    IFU_U48_GATE1_IFU_U48_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(3) , 
      O => IFU_U48_GATE1_2_0 ) ;
    IFU_U48_GATE1_IFU_U48_GATE1 : X_AND2 
      port map ( I0 => IFU_U48_GATE1_2_0 , 
      I1 => IFU_U48_GATE1_IFU_U48_GATE1_1_INV , O => IFU_U48_GATE1 ) ;
    IFU_U48_GATE2_IFU_U48_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(3) , O => IFU_U48_GATE2_2_0 ) ;
    IFU_U48_GATE2_IFU_U48_GATE2 : X_AND2 
      port map ( I0 => IFU_U48_GATE2_2_0 , I1 => JDEC , O => IFU_U48_GATE2 ) ;
    IFU_U49_O : X_OR2 
      port map ( I0 => IFU_U49_GATE1 , I1 => IFU_U49_GATE2 , O => IFU_TPC35(2) 
      ) ;
    IFU_U49_GATE1_IFU_U49_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(2) , 
      O => IFU_U49_GATE1_2_0 ) ;
    IFU_U49_GATE1_IFU_U49_GATE1 : X_AND2 
      port map ( I0 => IFU_U49_GATE1_2_0 , 
      I1 => IFU_U49_GATE1_IFU_U49_GATE1_1_INV , O => IFU_U49_GATE1 ) ;
    IFU_U49_GATE2_IFU_U49_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(2) , O => IFU_U49_GATE2_2_0 ) ;
    IFU_U49_GATE2_IFU_U49_GATE2 : X_AND2 
      port map ( I0 => IFU_U49_GATE2_2_0 , I1 => JDEC , O => IFU_U49_GATE2 ) ;
    IFU_U50_O : X_OR2 
      port map ( I0 => IFU_U50_GATE1 , I1 => IFU_U50_GATE2 , O => IFU_TPC35(1) 
      ) ;
    IFU_U50_GATE1_IFU_U50_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(1) , 
      O => IFU_U50_GATE1_2_0 ) ;
    IFU_U50_GATE1_IFU_U50_GATE1 : X_AND2 
      port map ( I0 => IFU_U50_GATE1_2_0 , 
      I1 => IFU_U50_GATE1_IFU_U50_GATE1_1_INV , O => IFU_U50_GATE1 ) ;
    IFU_U50_GATE2_IFU_U50_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(1) , O => IFU_U50_GATE2_2_0 ) ;
    IFU_U50_GATE2_IFU_U50_GATE2 : X_AND2 
      port map ( I0 => IFU_U50_GATE2_2_0 , I1 => JDEC , O => IFU_U50_GATE2 ) ;
    IFU_U51_O : X_OR2 
      port map ( I0 => IFU_U51_GATE1 , I1 => IFU_U51_GATE2 , O => IFU_TPC35(0) 
      ) ;
    IFU_U51_GATE1_IFU_U51_GATE1_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => IFU_RETURN89(0) , 
      O => IFU_U51_GATE1_2_0 ) ;
    IFU_U51_GATE1_IFU_U51_GATE1 : X_AND2 
      port map ( I0 => IFU_U51_GATE1_2_0 , 
      I1 => IFU_U51_GATE1_IFU_U51_GATE1_1_INV , O => IFU_U51_GATE1 ) ;
    IFU_U51_GATE2_IFU_U51_GATE2_2_0 : X_AND2 
      port map ( I0 => IFU_N135 , I1 => JUMP_ADR(0) , O => IFU_U51_GATE2_2_0 ) ;
    IFU_U51_GATE2_IFU_U51_GATE2 : X_AND2 
      port map ( I0 => IFU_U51_GATE2_2_0 , I1 => JDEC , O => IFU_U51_GATE2 ) ;
    IDU_U35_O : X_OR2 
      port map ( I0 => IDU_U35_GATE1 , I1 => IDU_U35_GATE2 , O => IDU_N65 ) ;
    IDU_U35_GATE1_IDU_U35_GATE1_2_0 : X_AND2 
      port map ( I0 => IDU_N68 , I1 => IDU_N67 , O => IDU_U35_GATE1_2_0 ) ;
    IDU_U35_GATE1_IDU_U35_GATE1 : X_AND2 
      port map ( I0 => IDU_U35_GATE1_2_0 , I1 => IDU_I(0) , O => IDU_U35_GATE1 
      ) ;
    IDU_U35_GATE2_IDU_U35_GATE2_2_0 : X_AND2 
      port map ( I0 => IDU_N68 , I1 => IDU_N67 , O => IDU_U35_GATE2_2_0 ) ;
    IDU_U35_GATE2_IDU_U35_GATE2 : X_AND2 
      port map ( I0 => IDU_U35_GATE2_2_0 , I1 => IDU_N66 , O => IDU_U35_GATE2 
      ) ;
    IDU_U44_O : X_INV 
      port map ( I => IDU_I(5) , O => IDU_N97 ) ;
    IDU_U46_O : X_INV 
      port map ( I => IDU_I(4) , O => IDU_N61 ) ;
    IDU_U48_O : X_INV 
      port map ( I => IDU_I(1) , O => IDU_N92 ) ;
    IDU_U49_O : X_INV 
      port map ( I => IDU_I(6) , O => IDU_N98 ) ;
    IDU_U50_O : X_INV 
      port map ( I => IDU_I(3) , O => IDU_N99 ) ;
    IDU_U51_O : X_INV 
      port map ( I => IDU_I(2) , O => IDU_N100 ) ;
    IDU_U52_O : X_INV 
      port map ( I => IDU_I(0) , O => IDU_N93 ) ;
    IDU_U63_O : X_INV 
      port map ( I => IDU_N89 , O => CTR_1(1) ) ;
    IDU_U65_O : X_INV 
      port map ( I => IDU_N90 , O => CTR_1(0) ) ;
    IDU_U69_O : X_INV 
      port map ( I => CTR_1(9) , O => IDU_N69 ) ;
    IDU_U71_O : X_INV 
      port map ( I => IDU_N66 , O => IDU_N104 ) ;
    IDU_U72_O : X_INV 
      port map ( I => IDU_N65 , O => CTR_1(11) ) ;
    IDU_U73_O : X_INV 
      port map ( I => CTR_1(10) , O => IDU_N64 ) ;
    PSU_U33_GATE1_446 : X_AND2 
      port map ( I0 => PSU_STEP1 , I1 => PSU_N91 , O => PSU_U33_GATE1 ) ;
    PSU_U33_O : X_OR2 
      port map ( I0 => PSU_U33_GATE1 , I1 => PSU_GO_A , O => PSU_EN_1 ) ;
    PSU_U34_O : X_INV 
      port map ( I => N127 , O => PSU_GO_A29 ) ;
    PSU_U35_O : X_INV 
      port map ( I => PSU_STEP2 , O => PSU_N91 ) ;
    PSU_STEP2_REG_1I13 : X_FF 
      port map ( I => PSU_STEP1 , CLK => N125 , CE => VCC , SET => GND , 
      RST => PSU_STEP2_REG_1I13_GSR_OR , O => PSU_STEP2 ) ;
    PSU_STEP2_REG_1I13_GSR_OR_1388 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => PSU_STEP2_REG_1I13_GSR_OR ) ;
    PSU_GO_A_REG_1I13 : X_FF 
      port map ( I => PSU_GO_A29 , CLK => N125 , CE => VCC , SET => GND , 
      RST => PSU_GO_A_REG_1I13_GSR_OR , O => PSU_GO_A ) ;
    PSU_GO_A_REG_1I13_GSR_OR_1389 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => PSU_GO_A_REG_1I13_GSR_OR ) ;
    PSU_EN_REG_1I13 : X_FF 
      port map ( I => PSU_EN_1 , CLK => N125 , CE => VCC , SET => GND , 
      RST => PSU_EN_REG_1I13_GSR_OR , O => EN ) ;
    PSU_EN_REG_1I13_GSR_OR_1390 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => PSU_EN_REG_1I13_GSR_OR ) ;
    PSU_STEP1_REG_1I13 : X_FF 
      port map ( I => N128 , CLK => N125 , CE => VCC , SET => GND , 
      RST => PSU_STEP1_REG_1I13_GSR_OR , O => PSU_STEP1 ) ;
    PSU_STEP1_REG_1I13_GSR_OR_1391 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => PSU_STEP1_REG_1I13_GSR_OR ) ;
    ALU_U129_O : X_OR2 
      port map ( I0 => ALU_U129_GATE1 , I1 => ALU_U129_GATE2 , O => ALU_B_IN(7) 
      ) ;
    ALU_U129_GATE1_ALU_U129_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N81 , O => ALU_U129_GATE1_2_0 ) ;
    ALU_U129_GATE1_ALU_U129_GATE1 : X_AND2 
      port map ( I0 => ALU_U129_GATE1_2_0 , 
      I1 => ALU_U129_GATE1_ALU_U129_GATE1_1_INV , O => ALU_U129_GATE1 ) ;
    ALU_U129_GATE2_ALU_U129_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(7) , O => ALU_U129_GATE2_2_0 
      ) ;
    ALU_U129_GATE2_ALU_U129_GATE2 : X_AND2 
      port map ( I0 => ALU_U129_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U129_GATE2 ) ;
    ALU_U130_O : X_OR2 
      port map ( I0 => ALU_U130_GATE1 , I1 => ALU_U130_GATE2 , O => ALU_B_IN(6) 
      ) ;
    ALU_U130_GATE1_ALU_U130_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N82 , O => ALU_U130_GATE1_2_0 ) ;
    ALU_U130_GATE1_ALU_U130_GATE1 : X_AND2 
      port map ( I0 => ALU_U130_GATE1_2_0 , 
      I1 => ALU_U130_GATE1_ALU_U130_GATE1_1_INV , O => ALU_U130_GATE1 ) ;
    ALU_U130_GATE2_ALU_U130_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(6) , O => ALU_U130_GATE2_2_0 
      ) ;
    ALU_U130_GATE2_ALU_U130_GATE2 : X_AND2 
      port map ( I0 => ALU_U130_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U130_GATE2 ) ;
    ALU_U131_O : X_OR2 
      port map ( I0 => ALU_U131_GATE1 , I1 => ALU_U131_GATE2 , O => ALU_B_IN(5) 
      ) ;
    ALU_U131_GATE1_ALU_U131_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N83 , O => ALU_U131_GATE1_2_0 ) ;
    ALU_U131_GATE1_ALU_U131_GATE1 : X_AND2 
      port map ( I0 => ALU_U131_GATE1_2_0 , 
      I1 => ALU_U131_GATE1_ALU_U131_GATE1_1_INV , O => ALU_U131_GATE1 ) ;
    ALU_U131_GATE2_ALU_U131_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(5) , O => ALU_U131_GATE2_2_0 
      ) ;
    ALU_U131_GATE2_ALU_U131_GATE2 : X_AND2 
      port map ( I0 => ALU_U131_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U131_GATE2 ) ;
    ALU_U132_O : X_OR2 
      port map ( I0 => ALU_U132_GATE1 , I1 => ALU_U132_GATE2 , O => ALU_B_IN(4) 
      ) ;
    ALU_U132_GATE1_ALU_U132_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N84 , O => ALU_U132_GATE1_2_0 ) ;
    ALU_U132_GATE1_ALU_U132_GATE1 : X_AND2 
      port map ( I0 => ALU_U132_GATE1_2_0 , 
      I1 => ALU_U132_GATE1_ALU_U132_GATE1_1_INV , O => ALU_U132_GATE1 ) ;
    ALU_U132_GATE2_ALU_U132_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(4) , O => ALU_U132_GATE2_2_0 
      ) ;
    ALU_U132_GATE2_ALU_U132_GATE2 : X_AND2 
      port map ( I0 => ALU_U132_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U132_GATE2 ) ;
    ALU_U133_O : X_OR2 
      port map ( I0 => ALU_U133_GATE1 , I1 => ALU_U133_GATE2 , O => ALU_B_IN(3) 
      ) ;
    ALU_U133_GATE1_ALU_U133_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N85 , O => ALU_U133_GATE1_2_0 ) ;
    ALU_U133_GATE1_ALU_U133_GATE1 : X_AND2 
      port map ( I0 => ALU_U133_GATE1_2_0 , 
      I1 => ALU_U133_GATE1_ALU_U133_GATE1_1_INV , O => ALU_U133_GATE1 ) ;
    ALU_U133_GATE2_ALU_U133_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(3) , O => ALU_U133_GATE2_2_0 
      ) ;
    ALU_U133_GATE2_ALU_U133_GATE2 : X_AND2 
      port map ( I0 => ALU_U133_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U133_GATE2 ) ;
    ALU_U134_O : X_OR2 
      port map ( I0 => ALU_U134_GATE1 , I1 => ALU_U134_GATE2 , O => ALU_B_IN(2) 
      ) ;
    ALU_U134_GATE1_ALU_U134_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N86 , O => ALU_U134_GATE1_2_0 ) ;
    ALU_U134_GATE1_ALU_U134_GATE1 : X_AND2 
      port map ( I0 => ALU_U134_GATE1_2_0 , 
      I1 => ALU_U134_GATE1_ALU_U134_GATE1_1_INV , O => ALU_U134_GATE1 ) ;
    ALU_U134_GATE2_ALU_U134_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(2) , O => ALU_U134_GATE2_2_0 
      ) ;
    ALU_U134_GATE2_ALU_U134_GATE2 : X_AND2 
      port map ( I0 => ALU_U134_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U134_GATE2 ) ;
    ALU_U135_O : X_OR2 
      port map ( I0 => ALU_U135_GATE1 , I1 => ALU_U135_GATE2 , O => ALU_B_IN(1) 
      ) ;
    ALU_U135_GATE1_ALU_U135_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N87 , O => ALU_U135_GATE1_2_0 ) ;
    ALU_U135_GATE1_ALU_U135_GATE1 : X_AND2 
      port map ( I0 => ALU_U135_GATE1_2_0 , 
      I1 => ALU_U135_GATE1_ALU_U135_GATE1_1_INV , O => ALU_U135_GATE1 ) ;
    ALU_U135_GATE2_ALU_U135_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(1) , O => ALU_U135_GATE2_2_0 
      ) ;
    ALU_U135_GATE2_ALU_U135_GATE2 : X_AND2 
      port map ( I0 => ALU_U135_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U135_GATE2 ) ;
    ALU_U136_O : X_OR2 
      port map ( I0 => ALU_U136_GATE1 , I1 => ALU_U136_GATE2 , O => ALU_B_IN(0) 
      ) ;
    ALU_U136_GATE1_ALU_U136_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N88 , O => ALU_U136_GATE1_2_0 ) ;
    ALU_U136_GATE1_ALU_U136_GATE1 : X_AND2 
      port map ( I0 => ALU_U136_GATE1_2_0 , 
      I1 => ALU_U136_GATE1_ALU_U136_GATE1_1_INV , O => ALU_U136_GATE1 ) ;
    ALU_U136_GATE2_ALU_U136_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => JUMP_ADR(0) , O => ALU_U136_GATE2_2_0 
      ) ;
    ALU_U136_GATE2_ALU_U136_GATE2 : X_AND2 
      port map ( I0 => ALU_U136_GATE2_2_0 , I1 => ALU_CTR_ALU(2) , 
      O => ALU_U136_GATE2 ) ;
    ALU_U137_O : X_OR2 
      port map ( I0 => ALU_U137_GATE1 , I1 => ALU_U137_GATE2 , O => ALU_N575 ) ;
    ALU_U137_GATE1_ALU_U137_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => ALU_ADD(8) , O => ALU_U137_GATE1_2_0 ) ;
    ALU_U137_GATE1_ALU_U137_GATE1 : X_AND2 
      port map ( I0 => ALU_U137_GATE1_2_0 , 
      I1 => ALU_U137_GATE1_ALU_U137_GATE1_1_INV , O => ALU_U137_GATE1 ) ;
    ALU_U137_GATE2_ALU_U137_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N334 , O => ALU_U137_GATE2_2_0 ) ;
    ALU_U137_GATE2_ALU_U137_GATE2 : X_AND2 
      port map ( I0 => ALU_U137_GATE2_2_0 , I1 => ALU_CTR_ALU(5) , 
      O => ALU_U137_GATE2 ) ;
    ALU_U138_O : X_OR2 
      port map ( I0 => ALU_U138_GATE1 , I1 => ALU_U138_GATE2 , O => ALU_F_IN(0) 
      ) ;
    ALU_U138_GATE1_ALU_U138_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => N350 , O => ALU_U138_GATE1_2_0 ) ;
    ALU_U138_GATE1_ALU_U138_GATE1 : X_AND2 
      port map ( I0 => ALU_U138_GATE1_2_0 , 
      I1 => ALU_U138_GATE1_ALU_U138_GATE1_1_INV , O => ALU_U138_GATE1 ) ;
    ALU_U138_GATE2_ALU_U138_GATE2_2_0 : X_AND2 
      port map ( I0 => ALU_N474 , I1 => ALU_N575 , O => ALU_U138_GATE2_2_0 ) ;
    ALU_U138_GATE2_ALU_U138_GATE2 : X_AND2 
      port map ( I0 => ALU_U138_GATE2_2_0 , I1 => ALU_CTR_ALU(6) , 
      O => ALU_U138_GATE2 ) ;
    ALU_U139_O : X_BUF 
      port map ( I => N336 , O => N318 ) ;
    ALU_U140_O : X_BUF 
      port map ( I => N340 , O => N322 ) ;
    ALU_U141_O : X_BUF 
      port map ( I => N338 , O => N320 ) ;
    ALU_U142_O : X_BUF 
      port map ( I => N334 , O => N316 ) ;
    ALU_U143_O : X_BUF 
      port map ( I => JUMP_ADR(0) , O => ADR(0) ) ;
    ALU_U144_O : X_BUF 
      port map ( I => JUMP_ADR(4) , O => ADR(4) ) ;
    ALU_U145_O : X_BUF 
      port map ( I => JUMP_ADR(6) , O => ADR(6) ) ;
    ALU_U146_O : X_BUF 
      port map ( I => JUMP_ADR(2) , O => ADR(2) ) ;
    ALU_U147_O : X_BUF 
      port map ( I => JUMP_ADR(3) , O => ADR(3) ) ;
    ALU_U148_O : X_BUF 
      port map ( I => JUMP_ADR(7) , O => ADR(7) ) ;
    ALU_U149_O : X_BUF 
      port map ( I => JUMP_ADR(5) , O => ADR(5) ) ;
    ALU_U150_O : X_BUF 
      port map ( I => N335 , O => N317 ) ;
    ALU_U151_O : X_BUF 
      port map ( I => JUMP_ADR(1) , O => ADR(1) ) ;
    ALU_U152_O : X_BUF 
      port map ( I => N341 , O => N323 ) ;
    ALU_U153_O : X_BUF 
      port map ( I => N339 , O => N321 ) ;
    ALU_U154_O : X_BUF 
      port map ( I => N337 , O => N319 ) ;
    ALU_U156_GATE1_500 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(2) , I1 => EN , O => ALU_U156_GATE1 ) ;
    ALU_U156_GATE2_501 : X_AND2 
      port map ( I0 => REG_CTR(1) , I1 => EN , O => ALU_U156_GATE2 ) ;
    ALU_U156_O : X_OR2 
      port map ( I0 => ALU_U156_GATE1 , I1 => ALU_U156_GATE2 , O => ALU_N_2432 
      ) ;
    ALU_U157_GATE1_503 : X_AND2 
      port map ( I0 => ALU_N491 , I1 => EN , O => ALU_U157_GATE1 ) ;
    ALU_U157_GATE2_504 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(4) , I1 => EN , O => ALU_U157_GATE2 ) ;
    ALU_U157_O : X_OR2 
      port map ( I0 => ALU_U157_GATE1 , I1 => ALU_U157_GATE2 , O => ALU_N_2164 
      ) ;
    ALU_U158_GATE1_506 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(1) , I1 => ALU_CTR_ALU(0) , 
      O => ALU_U158_GATE1 ) ;
    ALU_U158_GATE2_507 : X_AND2 
      port map ( I0 => N350 , I1 => ALU_CTR_ALU(0) , O => ALU_U158_GATE2 ) ;
    ALU_U158_GATE3_508 : X_AND2 
      port map ( I0 => N351 , I1 => ALU_CTR_ALU(1) , O => ALU_U158_GATE3 ) ;
    ALU_U158_O_JDEC_2_0 : X_OR2 
      port map ( I0 => ALU_U158_GATE3 , I1 => ALU_U158_GATE2 , 
      O => ALU_U158_O_2_0 ) ;
    ALU_U158_O_JDEC : X_OR2 
      port map ( I0 => ALU_U158_O_2_0 , I1 => ALU_U158_GATE1 , O => JDEC ) ;
    ALU_U160_O : X_INV 
      port map ( I => ALU_CTR_ALU(7) , O => ALU_N492 ) ;
    ALU_U161_O : X_INV 
      port map ( I => ALU_CTR_ALU(8) , O => ALU_N493 ) ;
    ALU_U163_O : X_INV 
      port map ( I => ALU_CTR_ALU(9) , O => ALU_N496 ) ;
    ALU_U171_O : X_INV 
      port map ( I => ALU_N491 , O => ALU_N495 ) ;
    ALU_U172_O : X_OR2 
      port map ( I0 => ALU_U172_GATE1 , I1 => ALU_N498 , O => ALU_N504 ) ;
    ALU_U172_GATE1_ALU_U172_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(9) , I1 => ALU_N493 , 
      O => ALU_U172_GATE1_2_0 ) ;
    ALU_U172_GATE1_ALU_U172_GATE1 : X_AND2 
      port map ( I0 => ALU_U172_GATE1_2_0 , I1 => ALU_CTR_ALU(7) , 
      O => ALU_U172_GATE1 ) ;
    ALU_U173_GATE1_516 : X_AND2 
      port map ( I0 => ALU_ADD(1) , I1 => ALU_N499 , O => ALU_U173_GATE1 ) ;
    ALU_U173_GATE2_517 : X_AND2 
      port map ( I0 => N341 , I1 => ALU_N504 , O => ALU_U173_GATE2 ) ;
    ALU_U173_O : X_OR2 
      port map ( I0 => ALU_U173_GATE1 , I1 => ALU_U173_GATE2 , O => ALU_N505 ) ;
    ALU_U175_O : X_INV 
      port map ( I => N348 , O => ALU_N507 ) ;
    ALU_U177_GATE1_522 : X_AND2 
      port map ( I0 => N348 , I1 => ALU_N494 , O => ALU_U177_GATE1 ) ;
    ALU_U177_O : X_OR2 
      port map ( I0 => ALU_U177_GATE1 , I1 => ALU_N503 , O => ALU_N509 ) ;
    ALU_U179_GATE1_528 : X_AND2 
      port map ( I0 => N348 , I1 => ALU_N501 , O => ALU_U179_GATE1 ) ;
    ALU_U179_GATE2_529 : X_AND2 
      port map ( I0 => N87 , I1 => ALU_N500 , O => ALU_U179_GATE2 ) ;
    ALU_U179_O : X_OR2 
      port map ( I0 => ALU_U179_GATE1 , I1 => ALU_U179_GATE2 , O => ALU_N511 ) ;
    ALU_U180_GATE1_531 : X_AND2 
      port map ( I0 => JUMP_ADR(1) , I1 => ALU_CTR_ALU(3) , O => ALU_U180_GATE1 
      ) ;
    ALU_U180_O : X_OR2 
      port map ( I0 => ALU_U180_GATE1 , I1 => ALU_N511 , O => ALU_N512 ) ;
    ALU_U182_GATE1_535 : X_AND2 
      port map ( I0 => ALU_ADD(3) , I1 => ALU_N499 , O => ALU_U182_GATE1 ) ;
    ALU_U182_GATE2_536 : X_AND2 
      port map ( I0 => N339 , I1 => ALU_N504 , O => ALU_U182_GATE2 ) ;
    ALU_U182_O : X_OR2 
      port map ( I0 => ALU_U182_GATE1 , I1 => ALU_U182_GATE2 , O => ALU_N513 ) ;
    ALU_U184_O : X_INV 
      port map ( I => N346 , O => ALU_N515 ) ;
    ALU_U186_GATE1_541 : X_AND2 
      port map ( I0 => N346 , I1 => ALU_N494 , O => ALU_U186_GATE1 ) ;
    ALU_U186_O : X_OR2 
      port map ( I0 => ALU_U186_GATE1 , I1 => ALU_N503 , O => ALU_N517 ) ;
    ALU_U188_GATE1_547 : X_AND2 
      port map ( I0 => N346 , I1 => ALU_N501 , O => ALU_U188_GATE1 ) ;
    ALU_U188_GATE2_548 : X_AND2 
      port map ( I0 => N85 , I1 => ALU_N500 , O => ALU_U188_GATE2 ) ;
    ALU_U188_O : X_OR2 
      port map ( I0 => ALU_U188_GATE1 , I1 => ALU_U188_GATE2 , O => ALU_N519 ) ;
    ALU_U189_GATE1_550 : X_AND2 
      port map ( I0 => JUMP_ADR(3) , I1 => ALU_CTR_ALU(3) , O => ALU_U189_GATE1 
      ) ;
    ALU_U189_O : X_OR2 
      port map ( I0 => ALU_U189_GATE1 , I1 => ALU_N519 , O => ALU_N520 ) ;
    ALU_U191_GATE1_554 : X_AND2 
      port map ( I0 => ALU_ADD(6) , I1 => ALU_N499 , O => ALU_U191_GATE1 ) ;
    ALU_U191_GATE2_555 : X_AND2 
      port map ( I0 => N336 , I1 => ALU_N504 , O => ALU_U191_GATE2 ) ;
    ALU_U191_O : X_OR2 
      port map ( I0 => ALU_U191_GATE1 , I1 => ALU_U191_GATE2 , O => ALU_N521 ) ;
    ALU_U193_O : X_INV 
      port map ( I => N343 , O => ALU_N523 ) ;
    ALU_U195_GATE1_560 : X_AND2 
      port map ( I0 => N343 , I1 => ALU_N494 , O => ALU_U195_GATE1 ) ;
    ALU_U195_O : X_OR2 
      port map ( I0 => ALU_U195_GATE1 , I1 => ALU_N503 , O => ALU_N525 ) ;
    ALU_U197_GATE1_566 : X_AND2 
      port map ( I0 => ALU_N501 , I1 => N343 , O => ALU_U197_GATE1 ) ;
    ALU_U197_GATE2_567 : X_AND2 
      port map ( I0 => N82 , I1 => ALU_N500 , O => ALU_U197_GATE2 ) ;
    ALU_U197_O : X_OR2 
      port map ( I0 => ALU_U197_GATE1 , I1 => ALU_U197_GATE2 , O => ALU_N527 ) ;
    ALU_U198_GATE1_569 : X_AND2 
      port map ( I0 => JUMP_ADR(6) , I1 => ALU_CTR_ALU(3) , O => ALU_U198_GATE1 
      ) ;
    ALU_U198_O : X_OR2 
      port map ( I0 => ALU_U198_GATE1 , I1 => ALU_N527 , O => ALU_N528 ) ;
    ALU_U200_GATE1_573 : X_AND2 
      port map ( I0 => ALU_ADD(5) , I1 => ALU_N499 , O => ALU_U200_GATE1 ) ;
    ALU_U200_GATE2_574 : X_AND2 
      port map ( I0 => N337 , I1 => ALU_N504 , O => ALU_U200_GATE2 ) ;
    ALU_U200_O : X_OR2 
      port map ( I0 => ALU_U200_GATE1 , I1 => ALU_U200_GATE2 , O => ALU_N529 ) ;
    ALU_U202_O : X_INV 
      port map ( I => N336 , O => ALU_N531 ) ;
    ALU_U203_GATE1_579 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N531 , O => ALU_U203_GATE1 ) ;
    ALU_U203_O : X_OR2 
      port map ( I0 => ALU_U203_GATE1 , I1 => ALU_N501 , O => ALU_N532 ) ;
    ALU_U204_GATE1_581 : X_AND2 
      port map ( I0 => N83 , I1 => ALU_N500 , O => ALU_U204_GATE1 ) ;
    ALU_U204_GATE2_582 : X_AND2 
      port map ( I0 => N344 , I1 => ALU_N532 , O => ALU_U204_GATE2 ) ;
    ALU_U204_O : X_OR2 
      port map ( I0 => ALU_U204_GATE1 , I1 => ALU_U204_GATE2 , O => ALU_N533 ) ;
    ALU_U205_O : X_INV 
      port map ( I => N344 , O => ALU_N534 ) ;
    ALU_U206_GATE1_585 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N534 , O => ALU_U206_GATE1 ) ;
    ALU_U206_O : X_OR2 
      port map ( I0 => ALU_U206_GATE1 , I1 => ALU_N502 , O => ALU_N535 ) ;
    ALU_U210_GATE1_592 : X_AND2 
      port map ( I0 => ALU_ADD(7) , I1 => ALU_N499 , O => ALU_U210_GATE1 ) ;
    ALU_U210_GATE2_593 : X_AND2 
      port map ( I0 => N335 , I1 => ALU_N504 , O => ALU_U210_GATE2 ) ;
    ALU_U210_O : X_OR2 
      port map ( I0 => ALU_U210_GATE1 , I1 => ALU_U210_GATE2 , O => ALU_N538 ) ;
    ALU_U211_O : X_OR2 
      port map ( I0 => ALU_U211_GATE1 , I1 => ALU_N538 , O => ALU_N539 ) ;
    ALU_U211_GATE1_ALU_U211_GATE1_2_0 : X_AND2 
      port map ( I0 => N342 , I1 => ALU_N497 , O => ALU_U211_GATE1_2_0 ) ;
    ALU_U211_GATE1_ALU_U211_GATE1 : X_AND2 
      port map ( I0 => ALU_U211_GATE1_2_0 , I1 => N334 , O => ALU_U211_GATE1 ) ;
    ALU_U212_O : X_INV 
      port map ( I => N334 , O => ALU_N540 ) ;
    ALU_U213_GATE1_598 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N540 , O => ALU_U213_GATE1 ) ;
    ALU_U213_O : X_OR2 
      port map ( I0 => ALU_U213_GATE1 , I1 => ALU_N501 , O => ALU_N541 ) ;
    ALU_U214_GATE1_600 : X_AND2 
      port map ( I0 => N81 , I1 => ALU_N500 , O => ALU_U214_GATE1 ) ;
    ALU_U214_GATE2_601 : X_AND2 
      port map ( I0 => N342 , I1 => ALU_N541 , O => ALU_U214_GATE2 ) ;
    ALU_U214_O : X_OR2 
      port map ( I0 => ALU_U214_GATE1 , I1 => ALU_U214_GATE2 , O => ALU_N542 ) ;
    ALU_U215_O : X_INV 
      port map ( I => N342 , O => ALU_N543 ) ;
    ALU_U216_GATE1_604 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N543 , O => ALU_U216_GATE1 ) ;
    ALU_U216_O : X_OR2 
      port map ( I0 => ALU_U216_GATE1 , I1 => ALU_N502 , O => ALU_N544 ) ;
    ALU_U220_GATE1_611 : X_AND2 
      port map ( I0 => ALU_ADD(4) , I1 => ALU_N499 , O => ALU_U220_GATE1 ) ;
    ALU_U220_GATE2_612 : X_AND2 
      port map ( I0 => N338 , I1 => ALU_N504 , O => ALU_U220_GATE2 ) ;
    ALU_U220_O : X_OR2 
      port map ( I0 => ALU_U220_GATE1 , I1 => ALU_U220_GATE2 , O => ALU_N547 ) ;
    ALU_U222_O : X_INV 
      port map ( I => N337 , O => ALU_N549 ) ;
    ALU_U223_GATE1_617 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N549 , O => ALU_U223_GATE1 ) ;
    ALU_U223_O : X_OR2 
      port map ( I0 => ALU_U223_GATE1 , I1 => ALU_N501 , O => ALU_N550 ) ;
    ALU_U224_GATE1_619 : X_AND2 
      port map ( I0 => N84 , I1 => ALU_N500 , O => ALU_U224_GATE1 ) ;
    ALU_U224_GATE2_620 : X_AND2 
      port map ( I0 => N345 , I1 => ALU_N550 , O => ALU_U224_GATE2 ) ;
    ALU_U224_O : X_OR2 
      port map ( I0 => ALU_U224_GATE1 , I1 => ALU_U224_GATE2 , O => ALU_N551 ) ;
    ALU_U225_O : X_INV 
      port map ( I => N345 , O => ALU_N552 ) ;
    ALU_U226_GATE1_623 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N552 , O => ALU_U226_GATE1 ) ;
    ALU_U226_O : X_OR2 
      port map ( I0 => ALU_U226_GATE1 , I1 => ALU_N502 , O => ALU_N553 ) ;
    ALU_U230_GATE1_630 : X_AND2 
      port map ( I0 => ALU_ADD(2) , I1 => ALU_N499 , O => ALU_U230_GATE1 ) ;
    ALU_U230_GATE2_631 : X_AND2 
      port map ( I0 => N340 , I1 => ALU_N504 , O => ALU_U230_GATE2 ) ;
    ALU_U230_O : X_OR2 
      port map ( I0 => ALU_U230_GATE1 , I1 => ALU_U230_GATE2 , O => ALU_N556 ) ;
    ALU_U232_O : X_INV 
      port map ( I => N339 , O => ALU_N558 ) ;
    ALU_U233_GATE1_636 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N558 , O => ALU_U233_GATE1 ) ;
    ALU_U233_O : X_OR2 
      port map ( I0 => ALU_U233_GATE1 , I1 => ALU_N501 , O => ALU_N559 ) ;
    ALU_U234_GATE1_638 : X_AND2 
      port map ( I0 => N86 , I1 => ALU_N500 , O => ALU_U234_GATE1 ) ;
    ALU_U234_GATE2_639 : X_AND2 
      port map ( I0 => N347 , I1 => ALU_N559 , O => ALU_U234_GATE2 ) ;
    ALU_U234_O : X_OR2 
      port map ( I0 => ALU_U234_GATE1 , I1 => ALU_U234_GATE2 , O => ALU_N560 ) ;
    ALU_U235_O : X_INV 
      port map ( I => N347 , O => ALU_N561 ) ;
    ALU_U236_GATE1_642 : X_AND2 
      port map ( I0 => ALU_N494 , I1 => ALU_N561 , O => ALU_U236_GATE1 ) ;
    ALU_U236_O : X_OR2 
      port map ( I0 => ALU_U236_GATE1 , I1 => ALU_N502 , O => ALU_N562 ) ;
    ALU_U240_O : X_INV 
      port map ( I => N349 , O => ALU_N565 ) ;
    ALU_U243_O : X_INV 
      port map ( I => N341 , O => ALU_N568 ) ;
    ALU_U244_GATE2_656 : X_AND2 
      port map ( I0 => ALU_N501 , I1 => N349 , O => ALU_U244_GATE2 ) ;
    ALU_U244_O : X_OR2 
      port map ( I0 => ALU_U244_GATE1 , I1 => ALU_U244_GATE2 , O => ALU_N569 ) ;
    ALU_U244_GATE1_ALU_U244_GATE1_2_0 : X_AND2 
      port map ( I0 => N349 , I1 => ALU_N568 , O => ALU_U244_GATE1_2_0 ) ;
    ALU_U244_GATE1_ALU_U244_GATE1 : X_AND2 
      port map ( I0 => ALU_U244_GATE1_2_0 , I1 => ALU_N494 , 
      O => ALU_U244_GATE1 ) ;
    ALU_U246_GATE1_658 : X_AND2 
      port map ( I0 => N350 , I1 => ALU_N498 , O => ALU_U246_GATE1 ) ;
    ALU_U246_GATE2_659 : X_AND2 
      port map ( I0 => ALU_N570 , I1 => ALU_N497 , O => ALU_U246_GATE2 ) ;
    ALU_U246_O : X_OR2 
      port map ( I0 => ALU_U246_GATE1 , I1 => ALU_U246_GATE2 , O => ALU_N571 ) ;
    ALU_U247_GATE2_662 : X_AND2 
      port map ( I0 => ALU_N571 , I1 => ALU_N495 , O => ALU_U247_GATE2 ) ;
    ALU_U247_O : X_OR2 
      port map ( I0 => ALU_U247_GATE1 , I1 => ALU_U247_GATE2 , O => ALU_N572 ) ;
    ALU_U247_GATE1_ALU_U247_GATE1_2_0 : X_AND2 
      port map ( I0 => ALU_N495 , I1 => ALU_N499 , O => ALU_U247_GATE1_2_0 ) ;
    ALU_U247_GATE1_ALU_U247_GATE1 : X_AND2 
      port map ( I0 => ALU_U247_GATE1_2_0 , I1 => ALU_ADD(0) , 
      O => ALU_U247_GATE1 ) ;
    ALU_U248_GATE1_664 : X_AND2 
      port map ( I0 => N88 , I1 => ALU_N500 , O => ALU_U248_GATE1 ) ;
    ALU_U248_O_ALU_N573_2_0 : X_OR2 
      port map ( I0 => ALU_N569 , I1 => ALU_N572 , O => ALU_U248_O_2_0 ) ;
    ALU_U248_O_ALU_N573 : X_OR2 
      port map ( I0 => ALU_U248_O_2_0 , I1 => ALU_U248_GATE1 , O => ALU_N573 ) ;
    MAU_U91_O : X_INV 
      port map ( I => N125 , O => MAU_N231 ) ;
    MAU_U92_O : X_INV 
      port map ( I => MAU_CTR_MAU(1) , O => MAU_N229 ) ;
    MAU_U93_O : X_INV 
      port map ( I => MAU_CTR_MAU(0) , O => MAU_N228 ) ;
    MAU_U94_GATE1_671 : X_AND2 
      port map ( I0 => MAU_U94_GATE1_0_INV , I1 => N325 , O => MAU_U94_GATE1 ) ;
    MAU_U94_GATE2_672 : X_AND2 
      port map ( I0 => MAU_N229 , I1 => EN , O => MAU_U94_GATE2 ) ;
    MAU_U94_GATE3_673 : X_AND2 
      port map ( I0 => MAU_CTR_MAU(0) , I1 => EN , O => MAU_U94_GATE3 ) ;
    MAU_U94_O_MAU_N232_2_0 : X_OR2 
      port map ( I0 => MAU_U94_GATE3 , I1 => MAU_U94_GATE2 , O => MAU_U94_O_2_0 
      ) ;
    MAU_U94_O_MAU_N232 : X_OR2 
      port map ( I0 => MAU_U94_O_2_0 , I1 => MAU_U94_GATE1 , O => MAU_N232 ) ;
    MAU_U95_GATE1_675 : X_AND2 
      port map ( I0 => MAU_U95_GATE1_0_INV , I1 => N324 , O => MAU_U95_GATE1 ) ;
    MAU_U95_GATE2_676 : X_AND2 
      port map ( I0 => MAU_N228 , I1 => EN , O => MAU_U95_GATE2 ) ;
    MAU_U95_GATE3_677 : X_AND2 
      port map ( I0 => MAU_CTR_MAU(1) , I1 => EN , O => MAU_U95_GATE3 ) ;
    MAU_U95_O_MAU_N230_2_0 : X_OR2 
      port map ( I0 => MAU_U95_GATE3 , I1 => MAU_U95_GATE2 , O => MAU_U95_O_2_0 
      ) ;
    MAU_U95_O_MAU_N230 : X_OR2 
      port map ( I0 => MAU_U95_O_2_0 , I1 => MAU_U95_GATE1 , O => MAU_N230 ) ;
    MAU_NRD_REG_1I13 : X_FF 
      port map ( I => MAU_N230 , CLK => MAU_N231 , CE => VCC , 
      SET => MAU_NRD_REG_1I13_GSR_OR , RST => GND , O => N324 ) ;
    MAU_NRD_REG_1I13_GSR_OR_1392 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_NRD_REG_1I13_GSR_OR ) ;
    MAU_NWR_REG_1I13 : X_FF 
      port map ( I => MAU_N232 , CLK => MAU_N231 , CE => VCC , 
      SET => MAU_NWR_REG_1I13_GSR_OR , RST => GND , O => N325 ) ;
    MAU_NWR_REG_1I13_GSR_OR_1393 : X_OR2 
      port map ( I0 => RST , I1 => GSR , O => MAU_NWR_REG_1I13_GSR_OR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_INV1_F_SUM_0 : X_INV 
      port map ( I => N315 , O => IFU_RETURN89(0) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_702 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C7 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_1_INV , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_703 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_C_704 : X_AND3 
      port map ( I0 => N309 , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_C ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_OUT_705 : X_OR3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_C , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND_706 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C1 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C0_AND_707 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C0 , 
      I1 => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT_708 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_AND_709 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_XOR_710 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F1_XOR_711 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F2_XOR , 
      I1 => N309 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND_712 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C2 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C3_AND_713 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C3 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_F1_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C3_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXB_OUT_714 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C3_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXB_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_CIN_AND_715 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_6 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_CIN_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND_716 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_OUT , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT0 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_CIN_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_7 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_AND_718 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_XOR_719 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_XOR_720 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G1_XOR , 
      I1 => GND , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_AND_721 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C6 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR_722 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT0_AND_723 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_7 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND_724 : X_AND2 
      port map ( I0 => VCC , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_COUT0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_COUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C0BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C1BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C1 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C2BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C2 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C3BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C3 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C4BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C4 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C5BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C5 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C6BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C6 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_C7BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C7 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_X_ZERO : X_ZERO 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ZERO ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_X_ONE : X_ONE 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_31_ONE ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_738 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C7 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_1_INV , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_739 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_C_740 : X_AND3 
      port map ( I0 => N311 , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_C ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_OUT_741 : X_OR3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_C , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND_742 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C1 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C0_AND_743 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C0 , 
      I1 => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT_744 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_AND_745 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_XOR_746 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F1_XOR_747 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F2_XOR , 
      I1 => N311 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND_748 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C2 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C3_AND_749 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C3 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_F1_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C3_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXB_OUT_750 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C3_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXB_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_CIN_AND_751 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_4 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_CIN_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND_752 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_OUT , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT0 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_CIN_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_5 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_AND_754 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_XOR_755 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_XOR_756 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G1_XOR , 
      I1 => N310 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_AND_757 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C6 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR_758 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT0_AND_759 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_5 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND_760 : X_AND2 
      port map ( I0 => N310 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_COUT0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_6 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C0BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C1BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C1 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C2BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C2 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C3BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C3 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C4BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C4 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C5BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C5 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C6BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C6 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_C7BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C7 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_X_ZERO : X_ZERO 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ZERO ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_X_ONE : X_ONE 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_32_ONE ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_774 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C7 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_1_INV , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_775 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_C_776 : X_AND3 
      port map ( I0 => N313 , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_C ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_OUT_777 : X_OR3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_C , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND_778 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C1 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C0_AND_779 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C0 , 
      I1 => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT_780 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_AND_781 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_XOR_782 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F1_XOR_783 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F2_XOR , 
      I1 => N313 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND_784 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C2 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C3_AND_785 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C3 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_F1_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C3_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXB_OUT_786 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C3_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXB_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_CIN_AND_787 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_2 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_CIN_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND_788 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_OUT , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT0 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_CIN_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_3 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_AND_790 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_XOR_791 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_XOR_792 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G1_XOR , 
      I1 => N312 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_AND_793 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C6 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR_794 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT0_AND_795 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_3 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND_796 : X_AND2 
      port map ( I0 => N312 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_COUT0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_4 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C0BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C1BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C1 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C2BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C2 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C3BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C3 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C4BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C4 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C5BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C5 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C6BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C6 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_C7BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C7 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_X_ZERO : X_ZERO 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ZERO ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_X_ONE : X_ONE 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_32_ONE ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_810 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C7 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_1_INV , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_811 : X_AND3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_C_812 : X_AND3 
      port map ( I0 => N315 , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C5 , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_C ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_OUT_813 : X_OR3 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B , 
      I2 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_C , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND_814 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C1 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C0_AND_815 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C0 , 
      I1 => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT_816 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_AND_817 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_XOR_818 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F1_XOR_819 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F2_XOR , 
      I1 => N315 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND_820 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C2 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C3_AND_821 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C3 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_F1_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C3_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXB_OUT_822 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C3_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXB_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_CIN_AND_823 : X_AND2 
      port map ( I0 => VCC , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_CIN_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND_824 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_OUT , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT0 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_CIN_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_1 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_AND_826 : X_AND2 
      port map ( I0 => VCC , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_XOR_827 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_XOR_828 : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G1_XOR , 
      I1 => N314 , O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_XOR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_AND_829 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C6 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_XOR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR_830 : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR_0_INV , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT0_AND_831 : X_AND2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_1 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT0_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND_832 : X_AND2 
      port map ( I0 => N314 , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND_1_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT : X_OR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_COUT0_AND , 
      I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_2 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C0BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C1BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C1 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C2BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C2 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C3BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C3 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C4BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C4 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C5BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C5 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C6BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C6 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_C7BUF : X_BUF 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C7 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_X_ZERO : X_ZERO 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ZERO ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_X_ONE : X_ONE 
      port map ( O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_33_ONE ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_7 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_2_0 , 
      I1 => N308 , O => IFU_RETURN89(7) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_6 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_2_0 , 
      I1 => N309 , O => IFU_RETURN89(6) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_5 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_2_0 , 
      I1 => N310 , O => IFU_RETURN89(5) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_2_0 , 
      I1 => N311 , O => IFU_RETURN89(4) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_3 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_2_0 , 
      I1 => N312 , O => IFU_RETURN89(3) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_2 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_2_0 , 
      I1 => N313 , O => IFU_RETURN89(2) ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_2_0 : X_XOR2 
      port map ( 
      I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_2_0_0_INV 
      , I1 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CO_1 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_2_0 ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_Q : X_XOR2 
      port map ( I0 => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_2_0 , 
      I1 => N314 , O => IFU_RETURN89(1) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_872 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_1_INV , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_873 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_C_874 : X_AND3 
      port map ( I0 => N334 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_C ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_OUT_875 : X_OR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_C , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND_876 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C1 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C0_AND_877 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C0 , 
      I1 => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT_878 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_AND_879 : X_AND2 
      port map ( I0 => N342 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_XOR_880 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F1_XOR_881 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F2_XOR , I1 => N334 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND_882 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C3_AND_883 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_F1_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C3_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXB_OUT_884 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C3_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXB_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_CIN_AND_885 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_8 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_CIN_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND_886 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_OUT , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT0 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_CIN_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_9 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_AND_888 : X_AND2 
      port map ( I0 => VCC , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_XOR_889 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_XOR_890 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G1_XOR , I1 => GND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_AND_891 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR_892 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT0_AND_893 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_9 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND_894 : X_AND2 
      port map ( I0 => VCC , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_COUT0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_COUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C0BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C1BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C2BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C2 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C3BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C4BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C5BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C6BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_C7BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_X_ZERO : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ZERO ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_X_ONE : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_12_ONE ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_908 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_1_INV , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_909 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_C_910 : X_AND3 
      port map ( I0 => N336 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_C ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_OUT_911 : X_OR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_C , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND_912 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C1 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C0_AND_913 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C0 , 
      I1 => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT_914 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_AND_915 : X_AND2 
      port map ( I0 => N344 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_XOR_916 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F1_XOR_917 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F2_XOR , I1 => N336 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND_918 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C3_AND_919 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_F1_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C3_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXB_OUT_920 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C3_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXB_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_CIN_AND_921 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_CIN_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND_922 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_OUT , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT0 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_CIN_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_AND_924 : X_AND2 
      port map ( I0 => N343 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_XOR_925 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_XOR_926 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G1_XOR , I1 => N335 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_AND_927 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR_928 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT0_AND_929 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND_930 : X_AND2 
      port map ( I0 => N335 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_COUT0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_8 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C0BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C1BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C2BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C2 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C3BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C4BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C5BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C6BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_C7BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_X_ZERO : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ZERO ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_X_ONE : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_13_ONE ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_944 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_1_INV , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_945 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_C_946 : X_AND3 
      port map ( I0 => N338 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_C ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_OUT_947 : X_OR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_C , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND_948 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C1 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C0_AND_949 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C0 , 
      I1 => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT_950 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_AND_951 : X_AND2 
      port map ( I0 => N346 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_XOR_952 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F1_XOR_953 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F2_XOR , I1 => N338 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND_954 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C3_AND_955 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_F1_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C3_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXB_OUT_956 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C3_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXB_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_CIN_AND_957 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_4 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_CIN_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND_958 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_OUT , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT0 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_CIN_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_AND_960 : X_AND2 
      port map ( I0 => N345 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_XOR_961 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_XOR_962 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G1_XOR , I1 => N337 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_AND_963 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR_964 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT0_AND_965 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_5 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND_966 : X_AND2 
      port map ( I0 => N337 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_COUT0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C0BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C1BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C2BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C2 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C3BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C4BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C5BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C6BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_C7BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_X_ZERO : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ZERO ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_X_ONE : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_13_ONE ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_980 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_1_INV , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_981 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_C_982 : X_AND3 
      port map ( I0 => N340 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_C ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_OUT_983 : X_OR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_C , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND_984 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C1 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C0_AND_985 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C0 , 
      I1 => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT_986 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_AND_987 : X_AND2 
      port map ( I0 => N348 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_XOR_988 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F1_XOR_989 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F2_XOR , I1 => N340 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND_990 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C3_AND_991 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_F1_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C3_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXB_OUT_992 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C3_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXB_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_CIN_AND_993 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_CIN_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND_994 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_OUT , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT0 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_CIN_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_AND_996 : X_AND2 
      port map ( I0 => N347 , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_XOR_997 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_XOR_998 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G1_XOR , I1 => N339 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_AND_999 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR_1000 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT0_AND_1001 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND_1002 : X_AND2 
      port map ( I0 => N339 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_COUT0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C0BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C1BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C2BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C2 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C3BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C4BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C5BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C6BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_C7BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_X_ZERO : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ZERO ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_X_ONE : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_13_ONE ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_1052 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C7 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_1_INV , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B_1053 : X_AND3 
      port map ( I0 => VCC , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_C_1054 : X_AND3 
      port map ( I0 => ALU_ADD_111_PLUS_N25 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C5 , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_C ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_OUT_1055 : X_OR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B , 
      I2 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_C , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND_1056 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C1 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C0_AND_1057 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C0 , I1 => VCC , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT_1058 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_AND_1059 : X_AND2 
      port map ( I0 => VCC , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_XOR_1060 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F1_XOR_1061 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F2_XOR , 
      I1 => ALU_ADD_111_PLUS_N25 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND_1062 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C2 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C3_AND_1063 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C3 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_F1_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C3_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXB_OUT_1064 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C3_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXB_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_CIN_AND_1065 : X_AND2 
      port map ( I0 => VCC , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXB_OUT 
      , O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_CIN_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND_1066 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_OUT , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT0 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_CIN_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_COUT0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_AND_1068 : X_AND2 
      port map ( I0 => VCC , I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_XOR_1069 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_XOR_1070 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G1_XOR , I1 => GND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_XOR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_AND_1071 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C6 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_XOR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR_1072 : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT0_AND_1073 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_COUT0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT0_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND_1074 : X_AND2 
      port map ( I0 => VCC , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND_1_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT : X_OR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_COUT0_AND , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C0BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C1BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C2BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C2 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C3BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C3 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C4BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C4 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C5BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ONE , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C5 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C6BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C6 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_C7BUF : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C7 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_X_ZERO : X_ZERO 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ZERO ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_X_ONE : X_ONE 
      port map ( O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_39_ONE ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_8 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_1 : X_XOR2 
      port map ( I0 => N342 , I1 => N334 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_2_1 , O => ALU_ADD(7) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_7 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_1 : X_XOR2 
      port map ( I0 => N343 , I1 => N335 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_2_1 , O => ALU_ADD(6) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_1 : X_XOR2 
      port map ( I0 => N344 , I1 => N336 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_2_1 , O => ALU_ADD(5) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_1 : X_XOR2 
      port map ( I0 => N345 , I1 => N337 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_2_1 , O => ALU_ADD(4) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_1 : X_XOR2 
      port map ( I0 => N346 , I1 => N338 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_2_1 , O => ALU_ADD(3) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_1 : X_XOR2 
      port map ( I0 => N347 , I1 => N339 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_2_1 , O => ALU_ADD(2) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_2 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_1 : X_XOR2 
      port map ( I0 => N348 , I1 => N340 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_1 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_2_1 , O => ALU_ADD(1) ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_2_0 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_2_0_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_CO_9 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_2_0 ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_Q : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_2_0 , 
      I1 => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_N25_1 , O => ALU_ADD(8) ) ;
    
    ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_N25_1 : X_XOR2 
      port map ( I0 => ALU_ADD_111_PLUS_N25 , I1 => ALU_ADD_111_PLUS_N25 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_N25_1 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_ALU_ADD_0_G , O => ALU_ADD(0) ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_COUT0 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_1N8 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A0BUF_1514 : X_BUF 
      port map ( I => N350 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A0BUF ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A1BUF_1515 : X_BUF 
      port map ( I => N341 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A1BUF ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B0BUF_1516 : X_BUF 
      port map ( I => ALU_CTR_ALU(10) , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B0BUF ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B1BUF_1517 : X_BUF 
      port map ( I => N349 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B1BUF ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND2_1518 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_S0_1_CO_0 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR1 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND2 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3_1519 : X_AND2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A0BUF , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_OR0 : X_OR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND2 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_COUT0 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_OR1 : X_OR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND4 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CO_2 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR2_1522 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV1 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B1BUF , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR2 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND4_1523 : X_AND2 
      port map ( I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_COUT0 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR3 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND4 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV1_1524 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV1 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5_1525 : X_AND2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5_0_INV , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A1BUF , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR3_1526 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR2 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A1BUF , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR3 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV0_1527 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV0 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR0_1528 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_INV0 , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_B0BUF , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR0 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR1_1529 : X_XOR2 
      port map ( 
      I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_A0BUF , 
      I1 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR0 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR1 ) ;
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_GLUT_XOR0 : X_XOR3 
      port map ( I0 => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_1N8 , I1 => N349 
      , I2 => N341 , O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_G ) ;
    U194_CLKBUF : X_CKBUF 
      port map ( I => U194_CLKIO_BUFSIG , O => N125 ) ;
    U194_CLKIO_BUF : X_BUF 
      port map ( I => CLK , O => U194_CLKIO_BUFSIG ) ;
    IDU_U33_CTR_1_14_2_0 : X_AND2 
      port map ( I0 => IDU_N60 , I1 => IDU_N61 , O => IDU_U33_2_0 ) ;
    IDU_U33_CTR_1_14_Q : X_AND2 
      port map ( I0 => IDU_U33_2_0 , I1 => IDU_N62 , O => CTR_1(14) ) ;
    IDU_U45_IDU_N62_2_0 : X_AND2 
      port map ( I0 => IDU_I(5) , I1 => IDU_N98 , O => IDU_U45_2_0 ) ;
    IDU_U45_IDU_N62_2_1 : X_AND2 
      port map ( I0 => IDU_N99 , I1 => IDU_N100 , O => IDU_U45_2_1 ) ;
    IDU_U45_IDU_N62 : X_AND2 
      port map ( I0 => IDU_U45_2_0 , I1 => IDU_U45_2_1 , O => IDU_N62 ) ;
    IDU_U55_IDU_N101_2_0 : X_AND2 
      port map ( I0 => IDU_N97 , I1 => IDU_N98 , O => IDU_U55_2_0 ) ;
    IDU_U55_IDU_N101 : X_AND2 
      port map ( I0 => IDU_U55_2_0 , I1 => IDU_I(4) , O => IDU_N101 ) ;
    IDU_U56_IDU_N102_2_0 : X_AND2 
      port map ( I0 => IDU_I(3) , I1 => IDU_N100 , O => IDU_U56_2_0 ) ;
    IDU_U56_IDU_N102 : X_AND2 
      port map ( I0 => IDU_U56_2_0 , I1 => IDU_N101 , O => IDU_N102 ) ;
    IDU_U58_IDU_N66_2_0 : X_AND2 
      port map ( I0 => IDU_I(2) , I1 => IDU_N99 , O => IDU_U58_2_0 ) ;
    IDU_U58_IDU_N66 : X_AND2 
      port map ( I0 => IDU_U58_2_0 , I1 => IDU_N101 , 
      O => IDU_U58_IDU_N66_2_INV ) ;
    IDU_U68_IDU_N67_2_0 : X_AND2 
      port map ( I0 => IDU_N92 , I1 => IDU_N93 , O => IDU_U68_2_0 ) ;
    IDU_U68_IDU_N67 : X_AND2 
      port map ( I0 => IDU_U68_2_0 , I1 => IDU_N102 , 
      O => IDU_U68_IDU_N67_2_INV ) ;
    IDU_U70_IDU_N68_2_0 : X_AND2 
      port map ( I0 => IDU_N61 , I1 => IDU_N92 , O => IDU_U70_2_0 ) ;
    IDU_U70_IDU_N68 : X_AND2 
      port map ( I0 => IDU_U70_2_0 , I1 => IDU_N62 , O => IDU_U70_IDU_N68_2_INV 
      ) ;
    ALU_U162_ALU_N494_2_0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(8) , I1 => ALU_CTR_ALU(7) , 
      O => ALU_U162_2_0 ) ;
    ALU_U162_ALU_N494_2_1 : X_AND2 
      port map ( I0 => ALU_N495 , I1 => ALU_N496 , O => ALU_U162_2_1 ) ;
    ALU_U162_ALU_N494 : X_AND2 
      port map ( I0 => ALU_U162_2_0 , I1 => ALU_U162_2_1 , O => ALU_N494 ) ;
    ALU_U165_ALU_N498_2_0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(8) , I1 => ALU_N492 , O => ALU_U165_2_0 ) ;
    ALU_U165_ALU_N498 : X_AND2 
      port map ( I0 => ALU_U165_2_0 , I1 => ALU_CTR_ALU(9) , O => ALU_N498 ) ;
    ALU_U166_ALU_N499_2_0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(8) , I1 => ALU_CTR_ALU(7) , 
      O => ALU_U166_2_0 ) ;
    ALU_U166_ALU_N499 : X_AND2 
      port map ( I0 => ALU_U166_2_0 , I1 => ALU_CTR_ALU(9) , O => ALU_N499 ) ;
    ALU_U168_ALU_N501_2_0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU(9) , I1 => ALU_N495 , O => ALU_U168_2_0 ) ;
    ALU_U168_ALU_N501_2_1 : X_AND2 
      port map ( I0 => ALU_N492 , I1 => ALU_N493 , O => ALU_U168_2_1 ) ;
    ALU_U168_ALU_N501 : X_AND2 
      port map ( I0 => ALU_U168_2_0 , I1 => ALU_U168_2_1 , O => ALU_N501 ) ;
    ALU_U169_ALU_N502_2_0 : X_AND2 
      port map ( I0 => ALU_N492 , I1 => ALU_N493 , O => ALU_U169_2_0 ) ;
    ALU_U169_ALU_N502 : X_AND2 
      port map ( I0 => ALU_U169_2_0 , I1 => ALU_N495 , O => ALU_N502 ) ;
    ALU_U250_ALU_N574_2_0 : X_OR2 
      port map ( I0 => ALU_A_IN(2) , I1 => ALU_A_IN(0) , O => ALU_U250_2_0 ) ;
    ALU_U250_ALU_N574_2_1 : X_OR2 
      port map ( I0 => ALU_A_IN(7) , I1 => ALU_A_IN(4) , O => ALU_U250_2_1 ) ;
    ALU_U250_ALU_N574 : X_OR2 
      port map ( I0 => ALU_U250_2_0 , I1 => ALU_U250_2_1 , O => ALU_N574 ) ;
    ALU_U251_ALU_F_IN_1_Q : X_OR2 
      port map ( I0 => ALU_U251_4_0 , I1 => ALU_A_IN(5) , 
      O => ALU_U251_ALU_F_IN_1_2_INV ) ;
    ALU_U251_ALU_F_IN_1_4_0_ALU_F_IN_1_4_0_2_0 : X_OR2 
      port map ( I0 => ALU_A_IN(6) , I1 => ALU_A_IN(3) , 
      O => ALU_U251_ALU_F_IN_1_4_0_2_0 ) ;
    ALU_U251_ALU_F_IN_1_4_0_ALU_F_IN_1_4_0_2_1 : X_OR2 
      port map ( I0 => ALU_A_IN(1) , I1 => ALU_N574 , 
      O => ALU_U251_ALU_F_IN_1_4_0_2_1 ) ;
    ALU_U251_ALU_F_IN_1_4_0_ALU_F_IN_1_4_0 : X_OR2 
      port map ( I0 => ALU_U251_ALU_F_IN_1_4_0_2_0 , 
      I1 => ALU_U251_ALU_F_IN_1_4_0_2_1 , O => ALU_U251_4_0 ) ;
    MAU_U90_MAU_N_2809_2_0 : X_AND2 
      port map ( I0 => MAU_N228 , I1 => MAU_N229 , O => MAU_U90_2_0 ) ;
    MAU_U90_MAU_N_2809 : X_AND2 
      port map ( I0 => MAU_U90_2_0 , I1 => EN , O => MAU_N_2809 ) ;
    STU_GSR_BUF : X_INV 
      port map ( I => STU_1_INV , O => GSR ) ;
    STU_GTS_BUF : X_BUF 
      port map ( I => NET4 , O => GTS ) ;
    ALU_N491_H0_1547 : X_BUF 
      port map ( I => ALU_N491_G , O => ALU_N491_H0 ) ;
    ALU_N491_H1_1548 : X_BUF 
      port map ( I => ALU_N539 , O => ALU_N491_H1 ) ;
    ALU_N491_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_N491_H , CLK => N125 , CE => ALU_N_2164 , SET => GND 
      , RST => GSR , O => N334 ) ;
    ALU_N491_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_N491_H , O => ALU_A_IN(7) ) ;
    ALU_N491_DFF_OUT_XMUX : X_BUF 
      port map ( I => ALU_N491_F , O => ALU_N491 ) ;
    ALU_N491_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_N542 , O => ALU_N491_FGBLOCK_1N8 ) ;
    ALU_N491_FGBLOCK_G3MUX : X_BUF 
      port map ( I => N334 , O => ALU_N491_FGBLOCK_1N7 ) ;
    ALU_N491_FGBLOCK_LUTRAM_FLUT_OR0 : X_OR2 
      port map ( I0 => ALU_CTR_ALU(3) , I1 => REG_CTR(0) , O => ALU_N491_F ) ;
    ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0_1540 : X_AND2 
      port map ( I0 => ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0_0_INV , I1 => ALU_N503 
      , O => ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_N491_FGBLOCK_LUTRAM_GLUT_OR1 : X_OR3 
      port map ( I0 => ALU_N491_FGBLOCK_1N8 , I1 => ALU_U218_O_2_0 , 
      I2 => ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0 , O => ALU_N491_G ) ;
    ALU_N491_HLUT_AND0_1545 : X_AND2 
      port map ( I0 => ALU_N491_HLUT_AND0_0_INV , I1 => ALU_N491_H1 , 
      O => ALU_N491_HLUT_AND0 ) ;
    ALU_N491_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_N491_H0 , I1 => ALU_N491_HLUT_AND0 , O => ALU_N491_H 
      ) ;
    ALU_A_IN_6_H0_1568 : X_BUF 
      port map ( I => ALU_A_IN_6_G , O => ALU_A_IN_6_H0 ) ;
    ALU_A_IN_6_H1_1569 : X_BUF 
      port map ( I => ALU_A_IN_6_3_INV , O => ALU_A_IN_6_H1 ) ;
    ALU_A_IN_6_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_A_IN_6_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N335 ) ;
    ALU_A_IN_6_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_A_IN_6_H , O => ALU_A_IN(6) ) ;
    ALU_A_IN_6_FGBLOCK_G2MUX : X_BUF 
      port map ( I => N343 , O => ALU_A_IN_6_FGBLOCK_1N8 ) ;
    ALU_A_IN_6_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_U196_GATE1 , O => ALU_A_IN_6_FGBLOCK_1N18 ) ;
    ALU_A_IN_6_FGBLOCK_G3MUX : X_BUF 
      port map ( I => N335 , O => ALU_A_IN_6_FGBLOCK_1N7 ) ;
    ALU_A_IN_6_FGBLOCK_LUTRAM_FLUT_OR0_1556 : X_OR2 
      port map ( I0 => ALU_U196_O_2_0 , I1 => ALU_A_IN_6_FGBLOCK_1N18 , 
      O => ALU_A_IN_6_FGBLOCK_LUTRAM_FLUT_OR0 ) ;
    ALU_A_IN_6_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_6_FGBLOCK_LUTRAM_FLUT_OR0 , I1 => ALU_N528 , 
      O => ALU_A_IN_6_F ) ;
    ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND0_1559 : X_AND2 
      port map ( I0 => ALU_A_IN_6_FGBLOCK_1N7 , I1 => ALU_N497 , 
      O => ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND1_1560 : X_AND2 
      port map ( I0 => ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => ALU_A_IN_6_FGBLOCK_1N8 , O => ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND1 
      ) ;
    ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_6_FGBLOCK_LUTRAM_GLUT_AND1 , I1 => ALU_N521 , 
      O => ALU_A_IN_6_G ) ;
    ALU_A_IN_6_HLUT_AND0_1566 : X_AND2 
      port map ( I0 => ALU_A_IN_6_HLUT_AND0_0_INV , I1 => ALU_A_IN_6_H0 , 
      O => ALU_A_IN_6_HLUT_AND0 ) ;
    ALU_A_IN_6_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_6_F , I1 => ALU_A_IN_6_HLUT_AND0 , 
      O => ALU_A_IN_6_H ) ;
    ALU_A_IN_5_H0_1589 : X_BUF 
      port map ( I => ALU_A_IN_5_G , O => ALU_A_IN_5_H0 ) ;
    ALU_A_IN_5_H1_1590 : X_BUF 
      port map ( I => ALU_A_IN_5_1_INV , O => ALU_A_IN_5_H1 ) ;
    ALU_A_IN_5_DFF_OUT_FFX : X_FF 
      port map ( I => ALU_A_IN_5_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N336 ) ;
    ALU_A_IN_5_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_A_IN_5_H , O => ALU_A_IN(5) ) ;
    ALU_A_IN_5_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_N497 , O => ALU_A_IN_5_FGBLOCK_1N8 ) ;
    ALU_A_IN_5_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_N533 , O => ALU_A_IN_5_FGBLOCK_1N18 ) ;
    ALU_A_IN_5_FGBLOCK_G3MUX : X_BUF 
      port map ( I => ALU_N529 , O => ALU_A_IN_5_FGBLOCK_1N7 ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0_1577 : X_AND2 
      port map ( I0 => ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => ALU_N503 , O => ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR3 
      port map ( I0 => ALU_A_IN_5_FGBLOCK_1N18 , I1 => ALU_U208_O_2_0 , 
      I2 => ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0 , O => ALU_A_IN_5_F ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND0_1580 : X_AND2 
      port map ( I0 => N344 , I1 => ALU_A_IN_5_FGBLOCK_1N8 , 
      O => ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND1_1581 : X_AND2 
      port map ( I0 => ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND0 , I1 => N336 , 
      O => ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND1 ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_5_FGBLOCK_LUTRAM_GLUT_AND1 , 
      I1 => ALU_A_IN_5_FGBLOCK_1N7 , O => ALU_A_IN_5_G ) ;
    ALU_A_IN_5_HLUT_AND0_1587 : X_AND2 
      port map ( I0 => ALU_A_IN_5_HLUT_AND0_0_INV , I1 => ALU_A_IN_5_H0 , 
      O => ALU_A_IN_5_HLUT_AND0 ) ;
    ALU_A_IN_5_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_5_F , I1 => ALU_A_IN_5_HLUT_AND0 , 
      O => ALU_A_IN_5_H ) ;
    ALU_A_IN_4_H0_1610 : X_BUF 
      port map ( I => ALU_A_IN_4_G , O => ALU_A_IN_4_H0 ) ;
    ALU_A_IN_4_H1_1611 : X_BUF 
      port map ( I => ALU_A_IN_4_3_INV , O => ALU_A_IN_4_H1 ) ;
    ALU_A_IN_4_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_A_IN_4_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N337 ) ;
    ALU_A_IN_4_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_A_IN_4_H , O => ALU_A_IN(4) ) ;
    ALU_A_IN_4_FGBLOCK_G2MUX : X_BUF 
      port map ( I => N345 , O => ALU_A_IN_4_FGBLOCK_1N8 ) ;
    ALU_A_IN_4_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_N503 , O => ALU_A_IN_4_FGBLOCK_1N18 ) ;
    ALU_A_IN_4_FGBLOCK_G3MUX : X_BUF 
      port map ( I => N337 , O => ALU_A_IN_4_FGBLOCK_1N7 ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0_1598 : X_AND2 
      port map ( I0 => ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => ALU_A_IN_4_FGBLOCK_1N18 , O => ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0 
      ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR3 
      port map ( I0 => ALU_N551 , I1 => ALU_U228_O_2_0 , 
      I2 => ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0 , O => ALU_A_IN_4_F ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND0_1601 : X_AND2 
      port map ( I0 => ALU_A_IN_4_FGBLOCK_1N8 , I1 => ALU_N497 , 
      O => ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND1_1602 : X_AND2 
      port map ( I0 => ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => ALU_A_IN_4_FGBLOCK_1N7 , O => ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND1 
      ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_4_FGBLOCK_LUTRAM_GLUT_AND1 , I1 => ALU_N547 , 
      O => ALU_A_IN_4_G ) ;
    ALU_A_IN_4_HLUT_AND0_1608 : X_AND2 
      port map ( I0 => ALU_A_IN_4_HLUT_AND0_0_INV , I1 => ALU_A_IN_4_H0 , 
      O => ALU_A_IN_4_HLUT_AND0 ) ;
    ALU_A_IN_4_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_4_F , I1 => ALU_A_IN_4_HLUT_AND0 , 
      O => ALU_A_IN_4_H ) ;
    ALU_A_IN_3_H0_1630 : X_BUF 
      port map ( I => ALU_A_IN_3_G , O => ALU_A_IN_3_H0 ) ;
    ALU_A_IN_3_H1_1631 : X_BUF 
      port map ( I => ALU_A_IN_3_0_INV , O => ALU_A_IN_3_H1 ) ;
    ALU_A_IN_3_DFF_OUT_FFX : X_FF 
      port map ( I => ALU_A_IN_3_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N338 ) ;
    ALU_A_IN_3_DFF_OUT_XMUX : X_BUF 
      port map ( I => ALU_A_IN_3_H , O => ALU_A_IN(3) ) ;
    ALU_A_IN_3_FGBLOCK_G2MUX : X_BUF 
      port map ( I => N346 , O => ALU_A_IN_3_FGBLOCK_1N8 ) ;
    ALU_A_IN_3_FGBLOCK_G3MUX : X_BUF 
      port map ( I => ALU_N513 , O => ALU_A_IN_3_FGBLOCK_1N7 ) ;
    ALU_A_IN_3_FGBLOCK_LUTRAM_FLUT_OR0_1619 : X_OR2 
      port map ( I0 => ALU_U187_O_2_0 , I1 => ALU_U187_GATE1 , 
      O => ALU_A_IN_3_FGBLOCK_LUTRAM_FLUT_OR0 ) ;
    ALU_A_IN_3_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_3_FGBLOCK_LUTRAM_FLUT_OR0 , I1 => ALU_N520 , 
      O => ALU_A_IN_3_F ) ;
    ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND0_1622 : X_AND2 
      port map ( I0 => N338 , I1 => ALU_N497 , 
      O => ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND1_1623 : X_AND2 
      port map ( I0 => ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => ALU_A_IN_3_FGBLOCK_1N8 , O => ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND1 
      ) ;
    ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_3_FGBLOCK_LUTRAM_GLUT_AND1 , 
      I1 => ALU_A_IN_3_FGBLOCK_1N7 , O => ALU_A_IN_3_G ) ;
    ALU_A_IN_3_HLUT_AND0_1628 : X_AND2 
      port map ( I0 => ALU_A_IN_3_HLUT_AND0_0_INV , I1 => ALU_A_IN_3_H0 , 
      O => ALU_A_IN_3_HLUT_AND0 ) ;
    ALU_A_IN_3_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_3_F , I1 => ALU_A_IN_3_HLUT_AND0 , 
      O => ALU_A_IN_3_H ) ;
    ALU_A_IN_2_H0_1651 : X_BUF 
      port map ( I => ALU_A_IN_2_G , O => ALU_A_IN_2_H0 ) ;
    ALU_A_IN_2_H1_1652 : X_BUF 
      port map ( I => ALU_A_IN_2_3_INV , O => ALU_A_IN_2_H1 ) ;
    ALU_A_IN_2_DFF_OUT_FFX : X_FF 
      port map ( I => ALU_A_IN_2_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N339 ) ;
    ALU_A_IN_2_DFF_OUT_XMUX : X_BUF 
      port map ( I => ALU_A_IN_2_H , O => ALU_A_IN(2) ) ;
    ALU_A_IN_2_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_N497 , O => ALU_A_IN_2_FGBLOCK_1N8 ) ;
    ALU_A_IN_2_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_N560 , O => ALU_A_IN_2_FGBLOCK_1N18 ) ;
    ALU_A_IN_2_FGBLOCK_G3MUX : X_BUF 
      port map ( I => N347 , O => ALU_A_IN_2_FGBLOCK_1N7 ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0_1639 : X_AND2 
      port map ( I0 => ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => ALU_N503 , O => ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR3 
      port map ( I0 => ALU_A_IN_2_FGBLOCK_1N18 , I1 => ALU_U238_O_2_0 , 
      I2 => ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0 , O => ALU_A_IN_2_F ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND0_1642 : X_AND2 
      port map ( I0 => ALU_A_IN_2_FGBLOCK_1N7 , I1 => ALU_A_IN_2_FGBLOCK_1N8 , 
      O => ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND1_1643 : X_AND2 
      port map ( I0 => ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND0 , I1 => N339 , 
      O => ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND1 ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_2_FGBLOCK_LUTRAM_GLUT_AND1 , I1 => ALU_N556 , 
      O => ALU_A_IN_2_G ) ;
    ALU_A_IN_2_HLUT_AND0_1649 : X_AND2 
      port map ( I0 => ALU_A_IN_2_HLUT_AND0_0_INV , I1 => ALU_A_IN_2_H0 , 
      O => ALU_A_IN_2_HLUT_AND0 ) ;
    ALU_A_IN_2_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_2_F , I1 => ALU_A_IN_2_HLUT_AND0 , 
      O => ALU_A_IN_2_H ) ;
    ALU_A_IN_1_H0_1672 : X_BUF 
      port map ( I => ALU_A_IN_1_G , O => ALU_A_IN_1_H0 ) ;
    ALU_A_IN_1_H1_1673 : X_BUF 
      port map ( I => ALU_A_IN_1_1_INV , O => ALU_A_IN_1_H1 ) ;
    ALU_A_IN_1_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_A_IN_1_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N340 ) ;
    ALU_A_IN_1_DFF_OUT_XMUX : X_BUF 
      port map ( I => ALU_A_IN_1_H , O => ALU_A_IN(1) ) ;
    ALU_A_IN_1_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_N505 , O => ALU_A_IN_1_FGBLOCK_1N8 ) ;
    ALU_A_IN_1_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_N512 , O => ALU_A_IN_1_FGBLOCK_1N18 ) ;
    ALU_A_IN_1_FGBLOCK_G3MUX : X_BUF 
      port map ( I => N340 , O => ALU_A_IN_1_FGBLOCK_1N7 ) ;
    ALU_A_IN_1_FGBLOCK_LUTRAM_FLUT_OR0_1660 : X_OR2 
      port map ( I0 => ALU_U178_O_2_0 , I1 => ALU_U178_GATE1 , 
      O => ALU_A_IN_1_FGBLOCK_LUTRAM_FLUT_OR0 ) ;
    ALU_A_IN_1_FGBLOCK_LUTRAM_FLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_1_FGBLOCK_LUTRAM_FLUT_OR0 , 
      I1 => ALU_A_IN_1_FGBLOCK_1N18 , O => ALU_A_IN_1_F ) ;
    ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND0_1663 : X_AND2 
      port map ( I0 => ALU_A_IN_1_FGBLOCK_1N7 , I1 => ALU_N497 , 
      O => ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND1_1664 : X_AND2 
      port map ( I0 => ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND0 , I1 => N348 , 
      O => ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND1 ) ;
    ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_1_FGBLOCK_LUTRAM_GLUT_AND1 , 
      I1 => ALU_A_IN_1_FGBLOCK_1N8 , O => ALU_A_IN_1_G ) ;
    ALU_A_IN_1_HLUT_AND0_1670 : X_AND2 
      port map ( I0 => ALU_A_IN_1_HLUT_AND0_0_INV , I1 => ALU_A_IN_1_H0 , 
      O => ALU_A_IN_1_HLUT_AND0 ) ;
    ALU_A_IN_1_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_1_F , I1 => ALU_A_IN_1_HLUT_AND0 , 
      O => ALU_A_IN_1_H ) ;
    ALU_A_IN_0_H0_1693 : X_BUF 
      port map ( I => ALU_CTR_ALU(3) , O => ALU_A_IN_0_H0 ) ;
    ALU_A_IN_0_H1_1694 : X_BUF 
      port map ( I => JUMP_ADR(0) , O => ALU_A_IN_0_H1 ) ;
    ALU_A_IN_0_DFF_OUT_FFX : X_FF 
      port map ( I => ALU_A_IN_0_H , CLK => N125 , CE => ALU_N_2164 , 
      SET => GND , RST => GSR , O => N341 ) ;
    ALU_A_IN_0_DFF_OUT_YMUX : X_BUF 
      port map ( I => ALU_A_IN_0_G , O => ALU_N503 ) ;
    ALU_A_IN_0_DFF_OUT_XMUX : X_BUF 
      port map ( I => ALU_A_IN_0_H , O => ALU_A_IN(0) ) ;
    ALU_A_IN_0_FGBLOCK_G2MUX : X_BUF 
      port map ( I => ALU_CTR_ALU(7) , O => ALU_A_IN_0_FGBLOCK_1N8 ) ;
    ALU_A_IN_0_FGBLOCK_F4MUX : X_BUF 
      port map ( I => ALU_N573 , O => ALU_A_IN_0_FGBLOCK_1N18 ) ;
    ALU_A_IN_0_FGBLOCK_G3MUX : X_BUF 
      port map ( I => ALU_A_IN_0_11_INV , O => ALU_A_IN_0_FGBLOCK_1N7 ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0_1681 : X_AND2 
      port map ( I0 => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => ALU_N503 , O => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_OR1_1682 : X_OR2 
      port map ( I0 => ALU_U242_O_2_0 , 
      I1 => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0 , 
      O => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_OR1 ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_OR2 : X_OR2 
      port map ( I0 => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_OR1 , 
      I1 => ALU_A_IN_0_FGBLOCK_1N18 , O => ALU_A_IN_0_F ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0_1685 : X_AND2 
      port map ( I0 => ALU_A_IN_0_FGBLOCK_1N8 , 
      I1 => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0_1_INV , 
      O => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1 : X_AND3 
      port map ( I0 => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_1_INV , 
      I2 => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_2_INV , O => ALU_A_IN_0_G ) ;
    ALU_A_IN_0_HLUT_AND0_1691 : X_AND2 
      port map ( I0 => ALU_A_IN_0_H1 , I1 => ALU_A_IN_0_H0 , 
      O => ALU_A_IN_0_HLUT_AND0 ) ;
    ALU_A_IN_0_HLUT_OR1 : X_OR2 
      port map ( I0 => ALU_A_IN_0_F , I1 => ALU_A_IN_0_HLUT_AND0 , 
      O => ALU_A_IN_0_H ) ;
    IDU_N71_H0_1721 : X_BUF 
      port map ( I => IDU_N71_G , O => IDU_N71_H0 ) ;
    IDU_N71_DFF_OUT_FFY : X_FF 
      port map ( I => IDU_N71_H , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(8) ) ;
    IDU_N71_DFF_OUT_XMUX : X_BUF 
      port map ( I => IDU_N71_F , O => IDU_N71 ) ;
    IDU_N71_FGBLOCK_G2MUX : X_BUF 
      port map ( I => IDU_N68 , O => IDU_N71_FGBLOCK_1N8 ) ;
    IDU_N71_FGBLOCK_G3MUX : X_BUF 
      port map ( I => IDU_I(0) , O => IDU_N71_FGBLOCK_1N7 ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND0_1706 : X_AND2 
      port map ( I0 => IDU_N102 , I1 => IDU_N71_2_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_1707 : X_AND2 
      port map ( I0 => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_0_INV , 
      I1 => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1 ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND2_1708 : X_AND2 
      port map ( I0 => IDU_N102 , I1 => IDU_N71_2_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND2 ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3_1709 : X_AND2 
      port map ( I0 => IDU_N66 , I1 => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3_1_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3 ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_OR4 : X_OR2 
      port map ( I0 => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1 , 
      I1 => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3 , O => IDU_N71_F ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_AND0_1712 : X_AND2 
      port map ( I0 => IDU_N71_FGBLOCK_1N7 , I1 => IDU_N71_FGBLOCK_1N8 , 
      O => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1_1713 : X_AND2 
      port map ( I0 => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1_0_INV , 
      I1 => IDU_N71_FGBLOCK_1N8 , O => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1 ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_OR2_1714 : X_OR2 
      port map ( I0 => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1 , 
      O => IDU_N71_FGBLOCK_LUTRAM_GLUT_OR2 ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_AND3_1715 : X_AND2 
      port map ( I0 => IDU_N66 , I1 => IDU_N71_FGBLOCK_1N8 , 
      O => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND3 ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_OR4 : X_OR2 
      port map ( I0 => IDU_N71_FGBLOCK_LUTRAM_GLUT_OR2 , 
      I1 => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND3 , O => IDU_N71_G ) ;
    IDU_N71_HLUT_AND0 : X_AND2 
      port map ( I0 => IDU_N71_F , I1 => IDU_N71_H0 , 
      O => IDU_N71_HLUT_AND0_2_INV ) ;
    CTR_1_9_H1_1733 : X_BUF 
      port map ( I => IDU_N68 , O => CTR_1_9_H1 ) ;
    CTR_1_9_DFF_OUT_FFY : X_FF 
      port map ( I => CTR_1_9_H , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(6) ) ;
    CTR_1_9_DFF_OUT_YMUX : X_BUF 
      port map ( I => CTR_1_9_H , O => CTR_1(10) ) ;
    CTR_1_9_DFF_OUT_XMUX : X_BUF 
      port map ( I => CTR_1_9_F , O => CTR_1(9) ) ;
    CTR_1_9_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_N71_2_INV , O => CTR_1_9_FGBLOCK_1N18 ) ;
    CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND0_1728 : X_AND2 
      port map ( I0 => IDU_N102 , I1 => CTR_1_9_FGBLOCK_1N18 , 
      O => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1 : X_AND2 
      port map ( I0 => IDU_N67 , I1 => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
      O => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_2_INV ) ;
    CTR_1_9_HLUT_AND0 : X_AND2 
      port map ( I0 => CTR_1_9_HLUT_AND0_0_INV , I1 => CTR_1_9_H1 , 
      O => CTR_1_9_HLUT_AND0_2_INV ) ;
    IDU_U76_O_SEC_B_2_0 : X_OR2 
      port map ( I0 => CTR_1(4) , I1 => IDU_N105 , O => IDU_U76_O_2_0 ) ;
    IDU_U76_O_SEC_B : X_OR2 
      port map ( I0 => IDU_U76_O_2_0 , I1 => IDU_U76_GATE1 , O => SEC_B ) ;
    IDU_N96_H0_1755 : X_BUF 
      port map ( I => IDU_I(1) , O => IDU_N96_H0 ) ;
    IDU_N96_H1_1756 : X_BUF 
      port map ( I => IDU_I(4) , O => IDU_N96_H1 ) ;
    IDU_N96_DFF_OUT_FFY : X_FF 
      port map ( I => IDU_N96_G , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(9) ) ;
    IDU_N96_DFF_OUT_YMUX : X_BUF 
      port map ( I => IDU_N96_H , O => IDU_U76_GATE1 ) ;
    IDU_N96_DFF_OUT_XMUX : X_BUF 
      port map ( I => IDU_N96_F , O => IDU_N96 ) ;
    IDU_N96_FGBLOCK_G2MUX : X_BUF 
      port map ( I => IDU_I(1) , O => IDU_N96_FGBLOCK_1N8 ) ;
    IDU_N96_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_I(3) , O => IDU_N96_FGBLOCK_1N18 ) ;
    IDU_N96_FGBLOCK_G3MUX : X_BUF 
      port map ( I => ALU_CTR_ALU_9_4_INV , O => IDU_N96_FGBLOCK_1N7 ) ;
    IDU_N96_FGBLOCK_LUTRAM_FLUT_AND0_1744 : X_AND2 
      port map ( I0 => IDU_I(2) , I1 => IDU_N96_FGBLOCK_1N18 , 
      O => IDU_N96_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    IDU_N96_FGBLOCK_LUTRAM_FLUT_AND1 : X_AND3 
      port map ( I0 => IDU_N96_FGBLOCK_LUTRAM_FLUT_AND0 , I1 => IDU_I(6) , 
      I2 => IDU_N96_FGBLOCK_LUTRAM_FLUT_AND1_2_INV , O => IDU_N96_F ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0_1747 : X_AND3 
      port map ( I0 => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0_0_INV , 
      I1 => IDU_N96_FGBLOCK_1N8 , I2 => IDU_I(0) , 
      O => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1 : X_AND2 
      port map ( I0 => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_0_INV , 
      I1 => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_1_INV , 
      O => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_2_INV ) ;
    IDU_N96_HLUT_AND0_1753 : X_AND2 
      port map ( I0 => IDU_N96_H1 , I1 => IDU_N96_F , O => IDU_N96_HLUT_AND0 ) ;
    IDU_N96_HLUT_AND1 : X_AND2 
      port map ( I0 => IDU_N96_HLUT_AND0 , I1 => IDU_N96_HLUT_AND1_1_INV , 
      O => IDU_N96_H ) ;
    ALU_CTR_ALU_4_H1_1769 : X_BUF 
      port map ( I => ALU_CTR_ALU_9_12_INV , O => ALU_CTR_ALU_4_H1 ) ;
    ALU_CTR_ALU_4_DFF_OUT_FFX : X_FF 
      port map ( I => CTR_1(9) , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(5) ) ;
    ALU_CTR_ALU_4_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_CTR_ALU_4_H , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(4) ) ;
    ALU_CTR_ALU_4_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_N71 , O => ALU_CTR_ALU_4_FGBLOCK_1N18 ) ;
    ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0_1764 : X_AND3 
      port map ( I0 => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => IDU_I(1) , I2 => IDU_I(0) , 
      O => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND1 : X_AND2 
      port map ( I0 => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND1_0_INV , 
      I1 => ALU_CTR_ALU_4_FGBLOCK_1N18 , O => ALU_CTR_ALU_4_F ) ;
    ALU_CTR_ALU_4_HLUT_AND0 : X_AND2 
      port map ( I0 => ALU_CTR_ALU_4_F , I1 => ALU_CTR_ALU_4_HLUT_AND0_1_INV , 
      O => ALU_CTR_ALU_4_HLUT_AND0_2_INV ) ;
    ALU_CTR_ALU_2_DFF_OUT_FFX : X_FF 
      port map ( I => ALU_CTR_ALU_2_G , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(3) ) ;
    ALU_CTR_ALU_2_DFF_OUT_FFY : X_FF 
      port map ( I => ALU_CTR_ALU_2_F , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(2) ) ;
    ALU_CTR_ALU_2_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_I(4) , O => ALU_CTR_ALU_2_FGBLOCK_1N18 ) ;
    ALU_CTR_ALU_2_FGBLOCK_G3MUX : X_BUF 
      port map ( I => IDU_N96 , O => ALU_CTR_ALU_2_FGBLOCK_1N7 ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND0_1776 : X_AND2 
      port map ( I0 => IDU_I(1) , I1 => IDU_I(0) , 
      O => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1_1777 : X_AND2 
      port map ( I0 => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND0 , 
      I1 => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1_1_INV , 
      O => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1 ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND2 : X_AND2 
      port map ( I0 => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1 , I1 => IDU_N96 , 
      O => ALU_CTR_ALU_2_F ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0_1780 : X_AND2 
      port map ( I0 => IDU_N60 , 
      I1 => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0_1_INV , 
      O => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND1 : X_AND2 
      port map ( I0 => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => ALU_CTR_ALU_2_FGBLOCK_1N7 , O => ALU_CTR_ALU_2_G ) ;
    CTR_1_0_H0_1800 : X_BUF 
      port map ( I => CTR_1_0_G , O => CTR_1_0_H0 ) ;
    CTR_1_0_DFF_OUT_FFX : X_FF 
      port map ( I => CTR_1_0_H , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => CTR_2(2) ) ;
    CTR_1_0_DFF_OUT_FFY : X_FF 
      port map ( I => CTR_1_0_G , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => CTR_2(1) ) ;
    CTR_1_0_DFF_OUT_XMUX : X_BUF 
      port map ( I => CTR_1_0_F , O => CTR_1_0_4299 ) ;
    CTR_1_0_FGBLOCK_G2MUX : X_BUF 
      port map ( I => IDU_N96 , O => CTR_1_0_FGBLOCK_1N8 ) ;
    CTR_1_0_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_N96 , O => CTR_1_0_FGBLOCK_1N18 ) ;
    CTR_1_0_FGBLOCK_G3MUX : X_BUF 
      port map ( I => IDU_I(4) , O => CTR_1_0_FGBLOCK_1N7 ) ;
    CTR_1_0_FGBLOCK_LUTRAM_FLUT_AND0_1790 : X_AND2 
      port map ( I0 => IDU_I(4) , I1 => CTR_1_0_FGBLOCK_1N18 , 
      O => CTR_1_0_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    CTR_1_0_FGBLOCK_LUTRAM_FLUT_AND1 : X_AND2 
      port map ( I0 => CTR_1_0_FGBLOCK_LUTRAM_FLUT_AND0 , I1 => IDU_N60 , 
      O => CTR_1_0_F ) ;
    CTR_1_0_FGBLOCK_LUTRAM_GLUT_AND0_1793 : X_AND2 
      port map ( I0 => CTR_1_0_FGBLOCK_1N7 , I1 => CTR_1_0_FGBLOCK_1N8 , 
      O => CTR_1_0_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    CTR_1_0_FGBLOCK_LUTRAM_GLUT_AND1 : X_AND3 
      port map ( I0 => CTR_1_0_FGBLOCK_LUTRAM_GLUT_AND0 , I1 => IDU_I(1) , 
      I2 => IDU_I(0) , O => CTR_1_0_G ) ;
    CTR_1_0_HLUT_AND0 : X_AND2 
      port map ( I0 => CTR_1_0_HLUT_AND0_0_INV , I1 => CTR_1_0_HLUT_AND0_1_INV 
      , O => CTR_1_0_HLUT_AND0_2_INV ) ;
    IDU_N105_DFF_OUT_FFX : X_FF 
      port map ( I => CTR_1_0_4299 , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => CTR_2(0) ) ;
    IDU_N105_DFF_OUT_FFY : X_FF 
      port map ( I => IDU_N105_F , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => CTR_2(3) ) ;
    IDU_N105_DFF_OUT_YMUX : X_BUF 
      port map ( I => IDU_N105_G , O => IDU_N105 ) ;
    IDU_N105_FGBLOCK_G2MUX : X_BUF 
      port map ( I => IDU_I(4) , O => IDU_N105_FGBLOCK_1N8 ) ;
    IDU_N105_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_I(1) , O => IDU_N105_FGBLOCK_1N18 ) ;
    IDU_N105_FGBLOCK_G3MUX : X_BUF 
      port map ( I => IDU_N96 , O => IDU_N105_FGBLOCK_1N7 ) ;
    IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_1808 : X_AND2 
      port map ( I0 => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_0_INV , 
      I1 => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_1_INV , 
      O => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0 ) ;
    IDU_N105_FGBLOCK_LUTRAM_FLUT_AND1 : X_AND3 
      port map ( I0 => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0 , I1 => IDU_I(4) , 
      I2 => IDU_N96 , O => IDU_N105_F ) ;
    IDU_N105_FGBLOCK_LUTRAM_GLUT_AND0_1811 : X_AND2 
      port map ( I0 => IDU_N105_FGBLOCK_1N7 , I1 => IDU_I(0) , 
      O => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    IDU_N105_FGBLOCK_LUTRAM_GLUT_AND1_1812 : X_AND2 
      port map ( I0 => IDU_N62 , I1 => IDU_N105_FGBLOCK_1N8 , 
      O => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND1 ) ;
    IDU_N105_FGBLOCK_LUTRAM_GLUT_AND2_1813 : X_AND2 
      port map ( I0 => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND1 , I1 => IDU_I(0) , 
      O => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND2 ) ;
    IDU_N105_FGBLOCK_LUTRAM_GLUT_OR3 : X_OR2 
      port map ( I0 => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => IDU_N105_FGBLOCK_LUTRAM_GLUT_AND2 , O => IDU_N105_G ) ;
    CTR_1_4_H0_1835 : X_BUF 
      port map ( I => CTR_1_4_G , O => CTR_1_4_H0 ) ;
    CTR_1_4_H1_1836 : X_BUF 
      port map ( I => IDU_I(0) , O => CTR_1_4_H1 ) ;
    CTR_1_4_DFF_OUT_FFX : X_FF 
      port map ( I => CTR_1_4_H , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(1) ) ;
    CTR_1_4_DFF_OUT_FFY : X_FF 
      port map ( I => CTR_1_4_G , CLK => N125 , CE => EN , SET => GND , 
      RST => GSR , O => ALU_CTR_ALU(0) ) ;
    CTR_1_4_DFF_OUT_YMUX : X_BUF 
      port map ( I => CTR_1_4_G , O => CTR_1(4) ) ;
    CTR_1_4_FGBLOCK_G2MUX : X_BUF 
      port map ( I => IDU_I(1) , O => CTR_1_4_FGBLOCK_1N8 ) ;
    CTR_1_4_FGBLOCK_F4MUX : X_BUF 
      port map ( I => IDU_N62 , O => CTR_1_4_FGBLOCK_1N18 ) ;
    CTR_1_4_FGBLOCK_G3MUX : X_BUF 
      port map ( I => IDU_I(4) , O => CTR_1_4_FGBLOCK_1N7 ) ;
    CTR_1_4_FGBLOCK_LUTRAM_FLUT_AND0 : X_AND3 
      port map ( I0 => IDU_N60 , I1 => CTR_1_4_FGBLOCK_1N18 , I2 => IDU_I(4) , 
      O => CTR_1_4_F ) ;
    CTR_1_4_FGBLOCK_LUTRAM_GLUT_AND0_1827 : X_AND2 
      port map ( I0 => IDU_N62 , I1 => CTR_1_4_FGBLOCK_1N7 , 
      O => CTR_1_4_FGBLOCK_LUTRAM_GLUT_AND0 ) ;
    CTR_1_4_FGBLOCK_LUTRAM_GLUT_AND1 : X_AND2 
      port map ( I0 => CTR_1_4_FGBLOCK_LUTRAM_GLUT_AND0 , 
      I1 => CTR_1_4_FGBLOCK_1N8 , O => CTR_1_4_G ) ;
    CTR_1_4_HLUT_AND0_1833 : X_AND2 
      port map ( I0 => CTR_1_4_H0 , I1 => CTR_1_4_H1 , O => CTR_1_4_HLUT_AND0 
      ) ;
    CTR_1_4_HLUT_OR1 : X_OR2 
      port map ( I0 => CTR_1_4_HLUT_AND0 , I1 => CTR_1_4_F , O => CTR_1_4_H ) ;
    IFU_U61_2_INV_1844 : X_INV 
      port map ( I => IFU_U61_2_INV , O => IFU_N136 ) ;
    ALU_U167_2_INV_1845 : X_INV 
      port map ( I => ALU_U167_2_INV , O => ALU_N500 ) ;
    ALU_U178_GATE1_0_INV_1846 : X_INV 
      port map ( I => N340 , O => ALU_U178_GATE1_0_INV ) ;
    ALU_U187_GATE1_0_INV_1847 : X_INV 
      port map ( I => N338 , O => ALU_U187_GATE1_0_INV ) ;
    ALU_U196_GATE1_0_INV_1848 : X_INV 
      port map ( I => N335 , O => ALU_U196_GATE1_0_INV ) ;
    MAU_U94_GATE1_0_INV_1849 : X_INV 
      port map ( I => EN , O => MAU_U94_GATE1_0_INV ) ;
    MAU_U95_GATE1_0_INV_1850 : X_INV 
      port map ( I => EN , O => MAU_U95_GATE1_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_1_INV_1851 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C5 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_2_INV_1852 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_A_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_0_INV_1853 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_2_INV_1854 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_AND3_B_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND_1_INV_1855 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C0 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C1_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT_2_INV_1856 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXA_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND_1_INV_1857 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C3 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C2_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND_1_INV_1858 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_MUXC_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR_0_INV_1859 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_C6 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND_1_INV_1860 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_3_CY4_G4_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_1_INV_1861 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C5 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_2_INV_1862 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_A_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_0_INV_1863 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_2_INV_1864 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_AND3_B_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND_1_INV_1865 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C0 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C1_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT_2_INV_1866 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXA_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND_1_INV_1867 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C3 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C2_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND_1_INV_1868 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_MUXC_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR_0_INV_1869 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_C6 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND_1_INV_1870 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_2_CY4_G4_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_1_INV_1871 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C5 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_2_INV_1872 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_A_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_0_INV_1873 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_2_INV_1874 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_AND3_B_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND_1_INV_1875 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C0 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C1_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT_2_INV_1876 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXA_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND_1_INV_1877 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C3 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C2_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND_1_INV_1878 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_MUXC_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR_0_INV_1879 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_C6 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND_1_INV_1880 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_1_CY4_G4_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_1_INV_1881 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C5 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_2_INV_1882 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_A_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_0_INV_1883 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_2_INV_1884 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C4 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_AND3_B_2_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND_1_INV_1885 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C0 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C1_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT_2_INV_1886 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT_2_INV , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXA_OUT ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND_1_INV_1887 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C3 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C2_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND_1_INV_1888 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXB_OUT , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_MUXC_AND_1_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR_0_INV_1889 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_C6 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR_0_INV ) ;
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND_1_INV_1890 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_C6_OR , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_CY4_0_CY4_G4_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_1_INV_1891 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_2_INV_1892 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_A_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_0_INV_1893 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_2_INV_1894 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_AND3_B_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND_1_INV_1895 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C0 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C1_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT_2_INV_1896 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXA_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND_1_INV_1897 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C2_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND_1_INV_1898 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_MUXC_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR_0_INV_1899 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_C6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND_1_INV_1900 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_5_CY4_G4_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_1_INV_1901 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_2_INV_1902 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_A_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_0_INV_1903 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_2_INV_1904 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_AND3_B_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND_1_INV_1905 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C0 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C1_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT_2_INV_1906 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXA_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND_1_INV_1907 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C2_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND_1_INV_1908 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_MUXC_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR_0_INV_1909 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_C6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND_1_INV_1910 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_4_CY4_G4_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_1_INV_1911 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_2_INV_1912 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_A_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_0_INV_1913 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_2_INV_1914 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_AND3_B_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND_1_INV_1915 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C0 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C1_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT_2_INV_1916 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXA_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND_1_INV_1917 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C2_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND_1_INV_1918 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_MUXC_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR_0_INV_1919 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_C6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND_1_INV_1920 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_3_CY4_G4_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_1_INV_1921 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_2_INV_1922 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_A_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_0_INV_1923 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_2_INV_1924 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_AND3_B_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND_1_INV_1925 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C0 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C1_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT_2_INV_1926 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXA_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND_1_INV_1927 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C2_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND_1_INV_1928 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_MUXC_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR_0_INV_1929 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_C6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND_1_INV_1930 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_2_CY4_G4_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_1_INV_1931 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C5 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_2_INV_1932 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_A_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B_2_INV_1933 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C4 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_AND3_B_2_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND_1_INV_1934 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C0 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C1_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT_2_INV_1935 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT_2_INV , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXA_OUT ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND_1_INV_1936 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C3 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C2_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND_1_INV_1937 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXB_OUT , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_MUXC_AND_1_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR_0_INV_1938 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_C6 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND_1_INV_1939 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_C6_OR , 
      O => ALU_ADD_111_PLUS_U10_S0_1_CY4_0_CY4_G4_AND_1_INV ) ;
    IFU_U44_GATE1_IFU_U44_GATE1_1_INV_1940 : X_INV 
      port map ( I => JDEC , O => IFU_U44_GATE1_IFU_U44_GATE1_1_INV ) ;
    IFU_U45_GATE1_IFU_U45_GATE1_1_INV_1941 : X_INV 
      port map ( I => JDEC , O => IFU_U45_GATE1_IFU_U45_GATE1_1_INV ) ;
    IFU_U46_GATE1_IFU_U46_GATE1_1_INV_1942 : X_INV 
      port map ( I => JDEC , O => IFU_U46_GATE1_IFU_U46_GATE1_1_INV ) ;
    IFU_U47_GATE1_IFU_U47_GATE1_1_INV_1943 : X_INV 
      port map ( I => JDEC , O => IFU_U47_GATE1_IFU_U47_GATE1_1_INV ) ;
    IFU_U48_GATE1_IFU_U48_GATE1_1_INV_1944 : X_INV 
      port map ( I => JDEC , O => IFU_U48_GATE1_IFU_U48_GATE1_1_INV ) ;
    IFU_U49_GATE1_IFU_U49_GATE1_1_INV_1945 : X_INV 
      port map ( I => JDEC , O => IFU_U49_GATE1_IFU_U49_GATE1_1_INV ) ;
    IFU_U50_GATE1_IFU_U50_GATE1_1_INV_1946 : X_INV 
      port map ( I => JDEC , O => IFU_U50_GATE1_IFU_U50_GATE1_1_INV ) ;
    IFU_U51_GATE1_IFU_U51_GATE1_1_INV_1947 : X_INV 
      port map ( I => JDEC , O => IFU_U51_GATE1_IFU_U51_GATE1_1_INV ) ;
    ALU_U129_GATE1_ALU_U129_GATE1_1_INV_1948 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U129_GATE1_ALU_U129_GATE1_1_INV 
      ) ;
    ALU_U130_GATE1_ALU_U130_GATE1_1_INV_1949 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U130_GATE1_ALU_U130_GATE1_1_INV 
      ) ;
    ALU_U131_GATE1_ALU_U131_GATE1_1_INV_1950 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U131_GATE1_ALU_U131_GATE1_1_INV 
      ) ;
    ALU_U132_GATE1_ALU_U132_GATE1_1_INV_1951 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U132_GATE1_ALU_U132_GATE1_1_INV 
      ) ;
    ALU_U133_GATE1_ALU_U133_GATE1_1_INV_1952 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U133_GATE1_ALU_U133_GATE1_1_INV 
      ) ;
    ALU_U134_GATE1_ALU_U134_GATE1_1_INV_1953 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U134_GATE1_ALU_U134_GATE1_1_INV 
      ) ;
    ALU_U135_GATE1_ALU_U135_GATE1_1_INV_1954 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U135_GATE1_ALU_U135_GATE1_1_INV 
      ) ;
    ALU_U136_GATE1_ALU_U136_GATE1_1_INV_1955 : X_INV 
      port map ( I => ALU_CTR_ALU(2) , O => ALU_U136_GATE1_ALU_U136_GATE1_1_INV 
      ) ;
    ALU_U137_GATE1_ALU_U137_GATE1_1_INV_1956 : X_INV 
      port map ( I => ALU_CTR_ALU(5) , O => ALU_U137_GATE1_ALU_U137_GATE1_1_INV 
      ) ;
    ALU_U138_GATE1_ALU_U138_GATE1_1_INV_1957 : X_INV 
      port map ( I => ALU_CTR_ALU(6) , O => ALU_U138_GATE1_ALU_U138_GATE1_1_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_2_0_0_INV_1958 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR7_G_SUM_3_IFU_RETURN89_7_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_2_0_0_INV_1959 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR6_F_SUM_3_IFU_RETURN89_6_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_2_0_0_INV_1960 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR5_G_SUM_2_IFU_RETURN89_5_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_2_0_0_INV_1961 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR4_F_SUM_2_IFU_RETURN89_4_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_2_0_0_INV_1962 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR3_G_SUM_1_IFU_RETURN89_3_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_2_0_0_INV_1963 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR2_F_SUM_1_IFU_RETURN89_2_2_0_0_INV 
      ) ;
    
    IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_2_0_0_INV_1964 : X_INV 
      port map ( I => IFU_ADD_59_PLUS_PLUS_N19 , 
      O => IFU_ADD_59_PLUS_PLUS_U8_S0_1_XOR1_G_SUM_0_IFU_RETURN89_1_2_0_0_INV 
      ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_0_0_INV_1965 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR9_F_SUM_5_ALU_ADD_7_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_0_0_INV_1966 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR8_G_SUM_4_ALU_ADD_6_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_0_0_INV_1967 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR7_F_SUM_4_ALU_ADD_5_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_0_0_INV_1968 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR6_G_SUM_3_ALU_ADD_4_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_0_0_INV_1969 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR5_F_SUM_3_ALU_ADD_3_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_0_0_INV_1970 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR4_G_SUM_2_ALU_ADD_2_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_0_0_INV_1971 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR3_F_SUM_2_ALU_ADD_1_2_0_0_INV ) ;
    ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_2_0_0_INV_1972 : X_INV 
      port map ( I => ALU_ADD_111_PLUS_N27 , 
      O => ALU_ADD_111_PLUS_U10_S0_1_XOR10_G_SUM_5_ALU_ADD_8_2_0_0_INV ) ;
    IDU_U58_IDU_N66_2_INV_1973 : X_INV 
      port map ( I => IDU_U58_IDU_N66_2_INV , O => IDU_N66 ) ;
    IDU_U68_IDU_N67_2_INV_1974 : X_INV 
      port map ( I => IDU_U68_IDU_N67_2_INV , O => IDU_N67 ) ;
    IDU_U70_IDU_N68_2_INV_1975 : X_INV 
      port map ( I => IDU_U70_IDU_N68_2_INV , O => IDU_N68 ) ;
    ALU_U251_ALU_F_IN_1_2_INV_1976 : X_INV 
      port map ( I => ALU_U251_ALU_F_IN_1_2_INV , O => ALU_F_IN(1) ) ;
    U134_1I20_GTS_TRI_2_INV_1977 : X_INV 
      port map ( I => GTS , O => U134_1I20_GTS_TRI_2_INV ) ;
    U135_1I20_GTS_TRI_2_INV_1978 : X_INV 
      port map ( I => GTS , O => U135_1I20_GTS_TRI_2_INV ) ;
    U136_1I20_GTS_TRI_2_INV_1979 : X_INV 
      port map ( I => GTS , O => U136_1I20_GTS_TRI_2_INV ) ;
    U137_1I20_GTS_TRI_2_INV_1980 : X_INV 
      port map ( I => GTS , O => U137_1I20_GTS_TRI_2_INV ) ;
    U138_1I20_GTS_TRI_2_INV_1981 : X_INV 
      port map ( I => GTS , O => U138_1I20_GTS_TRI_2_INV ) ;
    U139_1I20_GTS_TRI_2_INV_1982 : X_INV 
      port map ( I => GTS , O => U139_1I20_GTS_TRI_2_INV ) ;
    U140_1I20_GTS_TRI_2_INV_1983 : X_INV 
      port map ( I => GTS , O => U140_1I20_GTS_TRI_2_INV ) ;
    U141_1I20_GTS_TRI_2_INV_1984 : X_INV 
      port map ( I => GTS , O => U141_1I20_GTS_TRI_2_INV ) ;
    U158_1I20_GTS_TRI_2_INV_1985 : X_INV 
      port map ( I => GTS , O => U158_1I20_GTS_TRI_2_INV ) ;
    U159_1I20_GTS_TRI_2_INV_1986 : X_INV 
      port map ( I => GTS , O => U159_1I20_GTS_TRI_2_INV ) ;
    U160_1I20_GTS_TRI_2_INV_1987 : X_INV 
      port map ( I => GTS , O => U160_1I20_GTS_TRI_2_INV ) ;
    U161_1I20_GTS_TRI_2_INV_1988 : X_INV 
      port map ( I => GTS , O => U161_1I20_GTS_TRI_2_INV ) ;
    U162_1I20_GTS_TRI_2_INV_1989 : X_INV 
      port map ( I => GTS , O => U162_1I20_GTS_TRI_2_INV ) ;
    U163_1I20_GTS_TRI_2_INV_1990 : X_INV 
      port map ( I => GTS , O => U163_1I20_GTS_TRI_2_INV ) ;
    U164_1I20_GTS_TRI_2_INV_1991 : X_INV 
      port map ( I => GTS , O => U164_1I20_GTS_TRI_2_INV ) ;
    U165_1I20_GTS_TRI_2_INV_1992 : X_INV 
      port map ( I => GTS , O => U165_1I20_GTS_TRI_2_INV ) ;
    U166_1I20_GTS_TRI_2_INV_1993 : X_INV 
      port map ( I => GTS , O => U166_1I20_GTS_TRI_2_INV ) ;
    U167_1I20_GTS_TRI_2_INV_1994 : X_INV 
      port map ( I => GTS , O => U167_1I20_GTS_TRI_2_INV ) ;
    U168_1I20_GTS_TRI_2_INV_1995 : X_INV 
      port map ( I => GTS , O => U168_1I20_GTS_TRI_2_INV ) ;
    U169_1I20_GTS_TRI_2_INV_1996 : X_INV 
      port map ( I => GTS , O => U169_1I20_GTS_TRI_2_INV ) ;
    U170_1I20_GTS_TRI_2_INV_1997 : X_INV 
      port map ( I => GTS , O => U170_1I20_GTS_TRI_2_INV ) ;
    U171_1I20_GTS_TRI_2_INV_1998 : X_INV 
      port map ( I => GTS , O => U171_1I20_GTS_TRI_2_INV ) ;
    U172_1I20_GTS_TRI_2_INV_1999 : X_INV 
      port map ( I => GTS , O => U172_1I20_GTS_TRI_2_INV ) ;
    U173_1I20_GTS_TRI_2_INV_2000 : X_INV 
      port map ( I => GTS , O => U173_1I20_GTS_TRI_2_INV ) ;
    U174_1I20_GTS_TRI_2_INV_2001 : X_INV 
      port map ( I => GTS , O => U174_1I20_GTS_TRI_2_INV ) ;
    U175_1I20_GTS_TRI_2_INV_2002 : X_INV 
      port map ( I => GTS , O => U175_1I20_GTS_TRI_2_INV ) ;
    U176_1I20_GTS_TRI_2_INV_2003 : X_INV 
      port map ( I => GTS , O => U176_1I20_GTS_TRI_2_INV ) ;
    U177_1I20_GTS_TRI_2_INV_2004 : X_INV 
      port map ( I => GTS , O => U177_1I20_GTS_TRI_2_INV ) ;
    U178_1I20_GTS_TRI_2_INV_2005 : X_INV 
      port map ( I => GTS , O => U178_1I20_GTS_TRI_2_INV ) ;
    U179_1I20_GTS_TRI_2_INV_2006 : X_INV 
      port map ( I => GTS , O => U179_1I20_GTS_TRI_2_INV ) ;
    U180_1I20_GTS_TRI_2_INV_2007 : X_INV 
      port map ( I => GTS , O => U180_1I20_GTS_TRI_2_INV ) ;
    U181_1I20_GTS_TRI_2_INV_2008 : X_INV 
      port map ( I => GTS , O => U181_1I20_GTS_TRI_2_INV ) ;
    U182_1I20_GTS_TRI_2_INV_2009 : X_INV 
      port map ( I => GTS , O => U182_1I20_GTS_TRI_2_INV ) ;
    U183_1I20_GTS_TRI_2_INV_2010 : X_INV 
      port map ( I => GTS , O => U183_1I20_GTS_TRI_2_INV ) ;
    U184_1I20_GTS_TRI_2_INV_2011 : X_INV 
      port map ( I => GTS , O => U184_1I20_GTS_TRI_2_INV ) ;
    U185_1I20_GTS_TRI_2_INV_2012 : X_INV 
      port map ( I => GTS , O => U185_1I20_GTS_TRI_2_INV ) ;
    U186_1I20_GTS_TRI_2_INV_2013 : X_INV 
      port map ( I => GTS , O => U186_1I20_GTS_TRI_2_INV ) ;
    U187_1I20_GTS_TRI_2_INV_2014 : X_INV 
      port map ( I => GTS , O => U187_1I20_GTS_TRI_2_INV ) ;
    U188_1I20_GTS_TRI_2_INV_2015 : X_INV 
      port map ( I => GTS , O => U188_1I20_GTS_TRI_2_INV ) ;
    U189_1I20_GTS_TRI_2_INV_2016 : X_INV 
      port map ( I => GTS , O => U189_1I20_GTS_TRI_2_INV ) ;
    U190_1I20_GTS_TRI_2_INV_2017 : X_INV 
      port map ( I => GTS , O => U190_1I20_GTS_TRI_2_INV ) ;
    U191_1I20_GTS_TRI_2_INV_2018 : X_INV 
      port map ( I => GTS , O => U191_1I20_GTS_TRI_2_INV ) ;
    U192_1I20_GTS_TRI_2_INV_2019 : X_INV 
      port map ( I => GTS , O => U192_1I20_GTS_TRI_2_INV ) ;
    U193_1I20_GTS_TRI_2_INV_2020 : X_INV 
      port map ( I => GTS , O => U193_1I20_GTS_TRI_2_INV ) ;
    
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3_0_INV_2021 : X_INV 
      port map ( 
      I => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR1 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND3_0_INV ) ;
    
    ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5_0_INV_2022 : X_INV 
      port map ( 
      I => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_XOR3 , 
      O => ALU_ADD_111_PLUS_U10_ALU_ADD_0_FGBLOCK_LUTRAM_CARRYBLK_AND5_0_INV ) ;
    ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0_0_INV_2023 : X_INV 
      port map ( I => ALU_N491_FGBLOCK_1N7 , 
      O => ALU_N491_FGBLOCK_LUTRAM_GLUT_AND0_0_INV ) ;
    ALU_N491_HLUT_AND0_0_INV_2024 : X_INV 
      port map ( I => ALU_N491_F , O => ALU_N491_HLUT_AND0_0_INV ) ;
    ALU_A_IN_6_HLUT_AND0_0_INV_2025 : X_INV 
      port map ( I => ALU_A_IN_6_H1 , O => ALU_A_IN_6_HLUT_AND0_0_INV ) ;
    ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2026 : X_INV 
      port map ( I => N336 , O => ALU_A_IN_5_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    ALU_A_IN_5_HLUT_AND0_0_INV_2027 : X_INV 
      port map ( I => ALU_A_IN_5_H1 , O => ALU_A_IN_5_HLUT_AND0_0_INV ) ;
    ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2028 : X_INV 
      port map ( I => N337 , O => ALU_A_IN_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    ALU_A_IN_4_HLUT_AND0_0_INV_2029 : X_INV 
      port map ( I => ALU_A_IN_4_H1 , O => ALU_A_IN_4_HLUT_AND0_0_INV ) ;
    ALU_A_IN_3_HLUT_AND0_0_INV_2030 : X_INV 
      port map ( I => ALU_A_IN_3_H1 , O => ALU_A_IN_3_HLUT_AND0_0_INV ) ;
    ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2031 : X_INV 
      port map ( I => N339 , O => ALU_A_IN_2_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    ALU_A_IN_2_HLUT_AND0_0_INV_2032 : X_INV 
      port map ( I => ALU_A_IN_2_H1 , O => ALU_A_IN_2_HLUT_AND0_0_INV ) ;
    ALU_A_IN_1_HLUT_AND0_0_INV_2033 : X_INV 
      port map ( I => ALU_A_IN_1_H1 , O => ALU_A_IN_1_HLUT_AND0_0_INV ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2034 : X_INV 
      port map ( I => N341 , O => ALU_A_IN_0_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0_1_INV_2035 : X_INV 
      port map ( I => ALU_A_IN_0_9_INV , 
      O => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND0_1_INV ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_1_INV_2036 : X_INV 
      port map ( I => ALU_A_IN_0_FGBLOCK_1N7 , 
      O => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_1_INV ) ;
    ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_2_INV_2037 : X_INV 
      port map ( I => ALU_A_IN_0_12_INV , 
      O => ALU_A_IN_0_FGBLOCK_LUTRAM_GLUT_AND1_2_INV ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_0_INV_2038 : X_INV 
      port map ( I => IDU_N71_2_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_0_INV ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_1_INV_2039 : X_INV 
      port map ( I => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND0 , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND1_1_INV ) ;
    IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3_1_INV_2040 : X_INV 
      port map ( I => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND2 , 
      O => IDU_N71_FGBLOCK_LUTRAM_FLUT_AND3_1_INV ) ;
    IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1_0_INV_2041 : X_INV 
      port map ( I => IDU_N71_4_INV , 
      O => IDU_N71_FGBLOCK_LUTRAM_GLUT_AND1_0_INV ) ;
    IDU_N71_HLUT_AND0_2_INV_2042 : X_INV 
      port map ( I => IDU_N71_HLUT_AND0_2_INV , O => IDU_N71_H ) ;
    CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_1_INV_2043 : X_INV 
      port map ( I => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND0 , 
      O => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_1_INV ) ;
    CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_2_INV_2044 : X_INV 
      port map ( I => CTR_1_9_FGBLOCK_LUTRAM_FLUT_AND1_2_INV , O => CTR_1_9_F 
      ) ;
    CTR_1_9_HLUT_AND0_0_INV_2045 : X_INV 
      port map ( I => CTR_1_9_F , O => CTR_1_9_HLUT_AND0_0_INV ) ;
    CTR_1_9_HLUT_AND0_2_INV_2046 : X_INV 
      port map ( I => CTR_1_9_HLUT_AND0_2_INV , O => CTR_1_9_H ) ;
    IDU_N96_FGBLOCK_LUTRAM_FLUT_AND1_2_INV_2047 : X_INV 
      port map ( I => ALU_CTR_ALU_9_1_INV , 
      O => IDU_N96_FGBLOCK_LUTRAM_FLUT_AND1_2_INV ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0_0_INV_2048 : X_INV 
      port map ( I => ALU_CTR_ALU_9_5_INV , 
      O => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0_0_INV ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_0_INV_2049 : X_INV 
      port map ( I => IDU_N96_FGBLOCK_1N7 , 
      O => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_0_INV ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_1_INV_2050 : X_INV 
      port map ( I => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND0 , 
      O => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_1_INV ) ;
    IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_2_INV_2051 : X_INV 
      port map ( I => IDU_N96_FGBLOCK_LUTRAM_GLUT_AND1_2_INV , O => IDU_N96_G 
      ) ;
    IDU_N96_HLUT_AND1_1_INV_2052 : X_INV 
      port map ( I => IDU_N96_H0 , O => IDU_N96_HLUT_AND1_1_INV ) ;
    ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2053 : X_INV 
      port map ( I => ALU_CTR_ALU_9_5_INV , 
      O => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND1_0_INV_2054 : X_INV 
      port map ( I => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND0 , 
      O => ALU_CTR_ALU_4_FGBLOCK_LUTRAM_FLUT_AND1_0_INV ) ;
    ALU_CTR_ALU_4_HLUT_AND0_1_INV_2055 : X_INV 
      port map ( I => ALU_CTR_ALU_4_H1 , O => ALU_CTR_ALU_4_HLUT_AND0_1_INV ) ;
    ALU_CTR_ALU_4_HLUT_AND0_2_INV_2056 : X_INV 
      port map ( I => ALU_CTR_ALU_4_HLUT_AND0_2_INV , O => ALU_CTR_ALU_4_H ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1_1_INV_2057 : X_INV 
      port map ( I => ALU_CTR_ALU_2_FGBLOCK_1N18 , 
      O => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_FLUT_AND1_1_INV ) ;
    ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0_1_INV_2058 : X_INV 
      port map ( I => IDU_I(4) , 
      O => ALU_CTR_ALU_2_FGBLOCK_LUTRAM_GLUT_AND0_1_INV ) ;
    CTR_1_0_HLUT_AND0_0_INV_2059 : X_INV 
      port map ( I => CTR_1_0_F , O => CTR_1_0_HLUT_AND0_0_INV ) ;
    CTR_1_0_HLUT_AND0_1_INV_2060 : X_INV 
      port map ( I => CTR_1_0_H0 , O => CTR_1_0_HLUT_AND0_1_INV ) ;
    CTR_1_0_HLUT_AND0_2_INV_2061 : X_INV 
      port map ( I => CTR_1_0_HLUT_AND0_2_INV , O => CTR_1_0_H ) ;
    IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_0_INV_2062 : X_INV 
      port map ( I => IDU_N105_FGBLOCK_1N18 , 
      O => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_0_INV ) ;
    IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_1_INV_2063 : X_INV 
      port map ( I => IDU_I(0) , O => IDU_N105_FGBLOCK_LUTRAM_FLUT_AND0_1_INV 
      ) ;
    GND_2064 : X_ZERO 
      port map ( O => GND ) ;
    VCC_2065 : X_ONE 
      port map ( O => VCC ) ;
end STRUCTURE ;

