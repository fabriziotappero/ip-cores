-------------------------------------------------------------------------------
--
-- The Program Status Word (PSW).
-- Implements the PSW with its special bits.
--
-- $Id: psw-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_psw_rtl_c0 of t48_psw is

  for rtl
  end for;

end t48_psw_rtl_c0;
