-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             -- Internal ROM Memory --              #
-- #        Pre-installed bootloader available          #
-- # ************************************************** #
-- # Last modified: 24.05.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.STORM_core_package.all;

entity BOOT_ROM_FILE is
	generic	(
				MEM_SIZE      : natural := 1024;  -- memory cells
				LOG2_MEM_SIZE : natural := 10;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE; -- use output gate
				INIT_IMAGE_ID : string  := "-"    -- init image
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end BOOT_ROM_FILE;

architecture Behavioral of BOOT_ROM_FILE is

	--- Internal signals ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- ROM Type ---
	type BOOT_ROM_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);


-- ############################################################################
-- # STORM SoC Basic Configuration Bootloader                                 #
-- # 8*1024 byte ROM, 32*1024 byte RAM                                        #
-- ############################################################################
	constant STORM_SOC_BASIC_BL_32_8 : BOOT_ROM_TYPE :=
	(
		000000 => x"EA000006",
		000001 => x"EAFFFFFE",
		000002 => x"EAFFFFFE",
		000003 => x"EAFFFFFE",
		000004 => x"EAFFFFFE",
		000005 => x"E1A00000",
		000006 => x"EAFFFFFE",
		000007 => x"EAFFFFFE",
		000008 => x"E59F0034",
		000009 => x"E10F1000",
		000010 => x"E3C1107F",
		000011 => x"E38110DF",
		000012 => x"E129F001",
		000013 => x"E1A0D000",
		000014 => x"E3A00000",
		000015 => x"E1A01000",
		000016 => x"E1A02000",
		000017 => x"E1A0B000",
		000018 => x"E1A07000",
		000019 => x"E59FA00C",
		000020 => x"E1A0E00F",
		000021 => x"E1A0F00A",
		000022 => x"EAFFFFFE",
		000023 => x"00008000",
		000024 => x"FFF00700",
		000025 => x"E3E03A0F",
		000026 => x"E5131FFB",
		000027 => x"E20020FF",
		000028 => x"E3A00001",
		000029 => x"E0010210",
		000030 => x"E1A0F00E",
		000031 => x"E3E03A0F",
		000032 => x"E5130FFB",
		000033 => x"E1A0F00E",
		000034 => x"E3E01A0F",
		000035 => x"E5113FFF",
		000036 => x"E20000FF",
		000037 => x"E3A02001",
		000038 => x"E1833012",
		000039 => x"E5013FFF",
		000040 => x"E1A0F00E",
		000041 => x"E20000FF",
		000042 => x"E3A02001",
		000043 => x"E1A02012",
		000044 => x"E3E01A0F",
		000045 => x"E5113FFF",
		000046 => x"E1E02002",
		000047 => x"E0033002",
		000048 => x"E5013FFF",
		000049 => x"E1A0F00E",
		000050 => x"E3E01A0F",
		000051 => x"E5113FFF",
		000052 => x"E20000FF",
		000053 => x"E3A02001",
		000054 => x"E0233012",
		000055 => x"E5013FFF",
		000056 => x"E1A0F00E",
		000057 => x"E3E03A0F",
		000058 => x"E5030FFF",
		000059 => x"E1A0F00E",
		000060 => x"E20000FF",
		000061 => x"E3500007",
		000062 => x"E92D4010",
		000063 => x"E3A0C000",
		000064 => x"E3E0E0FF",
		000065 => x"E20110FF",
		000066 => x"8A000011",
		000067 => x"E2403004",
		000068 => x"E20330FF",
		000069 => x"E3500003",
		000070 => x"E1A0E183",
		000071 => x"E3E04A0F",
		000072 => x"E1A0C180",
		000073 => x"9A000007",
		000074 => x"E3A030FF",
		000075 => x"E1A03E13",
		000076 => x"E5142F8B",
		000077 => x"E1E03003",
		000078 => x"E0022003",
		000079 => x"E1822E11",
		000080 => x"E5042F8B",
		000081 => x"E8BD8010",
		000082 => x"E3A030FF",
		000083 => x"E1A03C13",
		000084 => x"E1E0E003",
		000085 => x"E3E02A0F",
		000086 => x"E5123F8F",
		000087 => x"E003300E",
		000088 => x"E1833C11",
		000089 => x"E5023F8F",
		000090 => x"E8BD8010",
		000091 => x"E20000FF",
		000092 => x"E3500007",
		000093 => x"E3A02000",
		000094 => x"8A00000A",
		000095 => x"E2403004",
		000096 => x"E3500003",
		000097 => x"E20320FF",
		000098 => x"9A000005",
		000099 => x"E3E03A0F",
		000100 => x"E5130F8B",
		000101 => x"E1A02182",
		000102 => x"E1A00230",
		000103 => x"E20000FF",
		000104 => x"E1A0F00E",
		000105 => x"E1A02180",
		000106 => x"E3E03A0F",
		000107 => x"E5130F8F",
		000108 => x"E1A00230",
		000109 => x"E20000FF",
		000110 => x"E1A0F00E",
		000111 => x"E3E02A0F",
		000112 => x"E5123FE3",
		000113 => x"E3130002",
		000114 => x"E3E00000",
		000115 => x"15120FE7",
		000116 => x"E1A0F00E",
		000117 => x"E3E02A0F",
		000118 => x"E5123FE3",
		000119 => x"E3130001",
		000120 => x"0AFFFFFC",
		000121 => x"E20030FF",
		000122 => x"E5023FE7",
		000123 => x"E1A0F00E",
		000124 => x"E20000FF",
		000125 => x"E3500001",
		000126 => x"E3812B01",
		000127 => x"03E03A0F",
		000128 => x"E3811B09",
		000129 => x"13E03A0F",
		000130 => x"05031FCF",
		000131 => x"15032FCF",
		000132 => x"E1A0F00E",
		000133 => x"E3E03A0F",
		000134 => x"E5030FCB",
		000135 => x"E1A0F00E",
		000136 => x"E3E02A0F",
		000137 => x"E5123FCF",
		000138 => x"E3130C01",
		000139 => x"1AFFFFFC",
		000140 => x"E5020FBF",
		000141 => x"E5123FCF",
		000142 => x"E3833C01",
		000143 => x"E5023FCF",
		000144 => x"E3E02A0F",
		000145 => x"E5123FCF",
		000146 => x"E3130C01",
		000147 => x"1AFFFFFC",
		000148 => x"E5120FBF",
		000149 => x"E1A0F00E",
		000150 => x"E3E01A0F",
		000151 => x"E5113FC7",
		000152 => x"E20000FF",
		000153 => x"E3A02001",
		000154 => x"E1833012",
		000155 => x"E5013FC7",
		000156 => x"E1A0F00E",
		000157 => x"E20000FF",
		000158 => x"E3A02001",
		000159 => x"E1A02012",
		000160 => x"E3E01A0F",
		000161 => x"E5113FC7",
		000162 => x"E1E02002",
		000163 => x"E0033002",
		000164 => x"E5013FC7",
		000165 => x"E1A0F00E",
		000166 => x"E3E02A0F",
		000167 => x"E5123F97",
		000168 => x"E1A01420",
		000169 => x"E3C33080",
		000170 => x"E5023F97",
		000171 => x"E5020F9F",
		000172 => x"E5021F9B",
		000173 => x"E5123F97",
		000174 => x"E3833080",
		000175 => x"E5023F97",
		000176 => x"E1A0F00E",
		000177 => x"E92D4030",
		000178 => x"E3A0C090",
		000179 => x"E20140FE",
		000180 => x"E3E0EA0F",
		000181 => x"E5DD500F",
		000182 => x"E20000FF",
		000183 => x"E50E4F93",
		000184 => x"E20110FF",
		000185 => x"E50ECFAF",
		000186 => x"E1A04002",
		000187 => x"E203C0FF",
		000188 => x"E51E3FAF",
		000189 => x"E3130002",
		000190 => x"1AFFFFFC",
		000191 => x"E51E3FAF",
		000192 => x"E3130080",
		000193 => x"13E00000",
		000194 => x"18BD8030",
		000195 => x"E35C0000",
		000196 => x"0A000012",
		000197 => x"E24C3001",
		000198 => x"E203C0FF",
		000199 => x"E35C0001",
		000200 => x"01A02424",
		000201 => x"03E03A0F",
		000202 => x"13E03A0F",
		000203 => x"05032F93",
		000204 => x"15034F93",
		000205 => x"E3E02A0F",
		000206 => x"E3A03010",
		000207 => x"E5023FAF",
		000208 => x"E5123FAF",
		000209 => x"E3130002",
		000210 => x"1AFFFFFC",
		000211 => x"E5123FAF",
		000212 => x"E3130080",
		000213 => x"0AFFFFEC",
		000214 => x"E3E00001",
		000215 => x"E8BD8030",
		000216 => x"E3500077",
		000217 => x"1A00000C",
		000218 => x"E3E03A0F",
		000219 => x"E3A02050",
		000220 => x"E5035F93",
		000221 => x"E5032FAF",
		000222 => x"E1A02003",
		000223 => x"E5123FAF",
		000224 => x"E3130002",
		000225 => x"1AFFFFFC",
		000226 => x"E5123FAF",
		000227 => x"E2130080",
		000228 => x"08BD8030",
		000229 => x"E3E00002",
		000230 => x"E8BD8030",
		000231 => x"E3500072",
		000232 => x"13E00003",
		000233 => x"18BD8030",
		000234 => x"E3813001",
		000235 => x"E3E02A0F",
		000236 => x"E3A01090",
		000237 => x"E5023F93",
		000238 => x"E5021FAF",
		000239 => x"E5123FAF",
		000240 => x"E3130002",
		000241 => x"1AFFFFFC",
		000242 => x"E5123FAF",
		000243 => x"E3130080",
		000244 => x"1AFFFFEF",
		000245 => x"E3A03068",
		000246 => x"E5023FAF",
		000247 => x"E3E00A0F",
		000248 => x"E5103FAF",
		000249 => x"E3130002",
		000250 => x"1AFFFFFC",
		000251 => x"E5100F93",
		000252 => x"E8BD8030",
		000253 => x"E20000FF",
		000254 => x"E350000D",
		000255 => x"979FF100",
		000256 => x"EA000015",
		000257 => x"FFF0043C",
		000258 => x"FFF00484",
		000259 => x"FFF0047C",
		000260 => x"FFF0045C",
		000261 => x"FFF0045C",
		000262 => x"FFF0045C",
		000263 => x"FFF00474",
		000264 => x"FFF0045C",
		000265 => x"FFF0046C",
		000266 => x"FFF00464",
		000267 => x"FFF0045C",
		000268 => x"FFF00454",
		000269 => x"FFF0044C",
		000270 => x"FFF00444",
		000271 => x"EE100F10",
		000272 => x"E1A0F00E",
		000273 => x"EE1D0F1D",
		000274 => x"E1A0F00E",
		000275 => x"EE1C0F1C",
		000276 => x"E1A0F00E",
		000277 => x"EE1B0F1B",
		000278 => x"E1A0F00E",
		000279 => x"E3A00000",
		000280 => x"E1A0F00E",
		000281 => x"EE190F19",
		000282 => x"E1A0F00E",
		000283 => x"EE180F18",
		000284 => x"E1A0F00E",
		000285 => x"EE160F16",
		000286 => x"E1A0F00E",
		000287 => x"EE120F12",
		000288 => x"E1A0F00E",
		000289 => x"EE110F11",
		000290 => x"E1A0F00E",
		000291 => x"E20110FF",
		000292 => x"E2411006",
		000293 => x"E3510007",
		000294 => x"979FF101",
		000295 => x"EA000008",
		000296 => x"FFF004C8",
		000297 => x"FFF004C4",
		000298 => x"FFF004C4",
		000299 => x"FFF004C4",
		000300 => x"FFF004C4",
		000301 => x"FFF004D0",
		000302 => x"FFF004D8",
		000303 => x"FFF004C0",
		000304 => x"EE0D0F1D",
		000305 => x"E1A0F00E",
		000306 => x"EE060F16",
		000307 => x"E1A0F00E",
		000308 => x"EE0B0F1B",
		000309 => x"E1A0F00E",
		000310 => x"EE0C0F1C",
		000311 => x"E1A0F00E",
		000312 => x"E10F0000",
		000313 => x"E1A0F00E",
		000314 => x"E129F000",
		000315 => x"E1A0F00E",
		000316 => x"E52DE004",
		000317 => x"EBFFFFF9",
		000318 => x"E3C00080",
		000319 => x"E49DE004",
		000320 => x"EAFFFFF8",
		000321 => x"E52DE004",
		000322 => x"EBFFFFF4",
		000323 => x"E3800080",
		000324 => x"E49DE004",
		000325 => x"EAFFFFF3",
		000326 => x"E92D4010",
		000327 => x"E1A04000",
		000328 => x"E5D00000",
		000329 => x"E3500000",
		000330 => x"1A000003",
		000331 => x"EA000005",
		000332 => x"E5F40001",
		000333 => x"E3500000",
		000334 => x"0A000002",
		000335 => x"EBFFFF24",
		000336 => x"E3500000",
		000337 => x"CAFFFFF9",
		000338 => x"E1A00004",
		000339 => x"E8BD8010",
		000340 => x"E92D4070",
		000341 => x"E2514000",
		000342 => x"E1A05000",
		000343 => x"E20260FF",
		000344 => x"D8BD8070",
		000345 => x"EBFFFF14",
		000346 => x"E3700001",
		000347 => x"E20030FF",
		000348 => x"0A000005",
		000349 => x"E3560001",
		000350 => x"E5C53000",
		000351 => x"E1A00003",
		000352 => x"E2855001",
		000353 => x"0A000003",
		000354 => x"E2444001",
		000355 => x"E3540000",
		000356 => x"CAFFFFF3",
		000357 => x"E8BD8070",
		000358 => x"EBFFFF0D",
		000359 => x"EAFFFFF9",
		000360 => x"E92D4030",
		000361 => x"E2514000",
		000362 => x"E1A05000",
		000363 => x"D8BD8030",
		000364 => x"E4D50001",
		000365 => x"EBFFFF06",
		000366 => x"E2544001",
		000367 => x"1AFFFFFB",
		000368 => x"E8BD8030",
		000369 => x"E92D4010",
		000370 => x"E20240FF",
		000371 => x"E3540008",
		000372 => x"83A04008",
		000373 => x"8A000001",
		000374 => x"E3540000",
		000375 => x"03A04001",
		000376 => x"E1A02001",
		000377 => x"E1A0E004",
		000378 => x"E1A0310E",
		000379 => x"E35E0001",
		000380 => x"E2433004",
		000381 => x"E1A0C000",
		000382 => x"81A0C330",
		000383 => x"E24E3001",
		000384 => x"E20CC00F",
		000385 => x"E203E0FF",
		000386 => x"E35C0009",
		000387 => x"E28C3030",
		000388 => x"828C3037",
		000389 => x"E35E0000",
		000390 => x"E4C23001",
		000391 => x"1AFFFFF1",
		000392 => x"E2443001",
		000393 => x"E20330FF",
		000394 => x"E0813003",
		000395 => x"E5C3E001",
		000396 => x"E8BD8010",
		000397 => x"E20110FF",
		000398 => x"E3510008",
		000399 => x"E92D4010",
		000400 => x"E1A04000",
		000401 => x"8A000016",
		000402 => x"E3510000",
		000403 => x"0A000014",
		000404 => x"E3A00000",
		000405 => x"EA000006",
		000406 => x"E2413001",
		000407 => x"E20310FF",
		000408 => x"E202200F",
		000409 => x"E1A03101",
		000410 => x"E3510000",
		000411 => x"E1800312",
		000412 => x"08BD8010",
		000413 => x"E4D43001",
		000414 => x"E2432030",
		000415 => x"E3520009",
		000416 => x"E243C041",
		000417 => x"9AFFFFF3",
		000418 => x"E35C0005",
		000419 => x"E243E061",
		000420 => x"E2432037",
		000421 => x"9AFFFFEF",
		000422 => x"E35E0005",
		000423 => x"E2432057",
		000424 => x"9AFFFFEC",
		000425 => x"E3A00000",
		000426 => x"E8BD8010",
		000427 => x"E1A03000",
		000428 => x"E5D00001",
		000429 => x"E283C001",
		000430 => x"E5D32000",
		000431 => x"E5DC1002",
		000432 => x"E1A00800",
		000433 => x"E1800C02",
		000434 => x"E5DC3001",
		000435 => x"E1800001",
		000436 => x"E1800403",
		000437 => x"E1A0F00E",
		000438 => x"E0603280",
		000439 => x"E0800103",
		000440 => x"E0800100",
		000441 => x"E1A00200",
		000442 => x"E3500000",
		000443 => x"D1A0F00E",
		000444 => x"E1A00000",
		000445 => x"E2500001",
		000446 => x"1AFFFFFC",
		000447 => x"E1A0F00E",
		000448 => x"E92D45F0",
		000449 => x"E3A00000",
		000450 => x"E24DD00C",
		000451 => x"EBFFFE74",
		000452 => x"E3A0100D",
		000453 => x"E3A000C3",
		000454 => x"EBFFFF5B",
		000455 => x"E3A00063",
		000456 => x"EBFFFEDC",
		000457 => x"E3A00006",
		000458 => x"EBFFFF31",
		000459 => x"E3A01006",
		000460 => x"E3800008",
		000461 => x"EBFFFF54",
		000462 => x"E3A0000D",
		000463 => x"EBFFFF2C",
		000464 => x"E1A008A0",
		000465 => x"E1E00000",
		000466 => x"E200000F",
		000467 => x"E3500001",
		000468 => x"03A04030",
		000469 => x"028DA007",
		000470 => x"0A00001A",
		000471 => x"E3500002",
		000472 => x"0A000070",
		000473 => x"E59F07E8",
		000474 => x"EBFFFF6A",
		000475 => x"E59F07E4",
		000476 => x"EBFFFF68",
		000477 => x"E59F07E0",
		000478 => x"EBFFFF66",
		000479 => x"E59F07DC",
		000480 => x"EBFFFF64",
		000481 => x"E59F07D8",
		000482 => x"EBFFFF62",
		000483 => x"E59F07D4",
		000484 => x"EBFFFF60",
		000485 => x"E59F07D0",
		000486 => x"EBFFFF5E",
		000487 => x"E59F07CC",
		000488 => x"EBFFFF5C",
		000489 => x"E59F07C8",
		000490 => x"EBFFFF5A",
		000491 => x"E59F07C4",
		000492 => x"EBFFFF58",
		000493 => x"E59F07C0",
		000494 => x"EBFFFF56",
		000495 => x"E28DA007",
		000496 => x"EBFFFE7D",
		000497 => x"E1A04000",
		000498 => x"E3A0000D",
		000499 => x"EBFFFF08",
		000500 => x"E3100801",
		000501 => x"03A06001",
		000502 => x"03A050A0",
		000503 => x"1A000035",
		000504 => x"E3A04000",
		000505 => x"E59F0794",
		000506 => x"EBFFFF4A",
		000507 => x"E1A01005",
		000508 => x"E1A02004",
		000509 => x"E3A03002",
		000510 => x"E3A00072",
		000511 => x"E58D4000",
		000512 => x"EBFFFEAF",
		000513 => x"E1A01005",
		000514 => x"E5CD0007",
		000515 => x"E3A02001",
		000516 => x"E3A03002",
		000517 => x"E3A00072",
		000518 => x"E58D4000",
		000519 => x"EBFFFEA8",
		000520 => x"E3A02002",
		000521 => x"E1A03002",
		000522 => x"E5CD0008",
		000523 => x"E1A01005",
		000524 => x"E3A00072",
		000525 => x"E58D4000",
		000526 => x"EBFFFEA1",
		000527 => x"E3A03002",
		000528 => x"E5CD0009",
		000529 => x"E1A01005",
		000530 => x"E3A00072",
		000531 => x"E3A02003",
		000532 => x"E58D4000",
		000533 => x"EBFFFE9A",
		000534 => x"E5DD3007",
		000535 => x"E20000FF",
		000536 => x"E3530053",
		000537 => x"E5CD000A",
		000538 => x"1A000002",
		000539 => x"E5DD3008",
		000540 => x"E353004D",
		000541 => x"0A000062",
		000542 => x"E59F0704",
		000543 => x"EBFFFF25",
		000544 => x"E3560000",
		000545 => x"0AFFFFCD",
		000546 => x"E59F06F8",
		000547 => x"EBFFFF21",
		000548 => x"E3A0100D",
		000549 => x"E3A00000",
		000550 => x"EBFFFEFB",
		000551 => x"E3A00006",
		000552 => x"EBFFFED3",
		000553 => x"E3A01006",
		000554 => x"E3C00008",
		000555 => x"EBFFFEF6",
		000556 => x"E3A0F000",
		000557 => x"EAFFFFFE",
		000558 => x"E3540034",
		000559 => x"0A000028",
		000560 => x"CA00001B",
		000561 => x"E3540031",
		000562 => x"0A000035",
		000563 => x"DA000096",
		000564 => x"E3540032",
		000565 => x"0A0000A0",
		000566 => x"E3540033",
		000567 => x"1A000096",
		000568 => x"E1A00004",
		000569 => x"EBFFFE3A",
		000570 => x"E59F069C",
		000571 => x"EBFFFF09",
		000572 => x"E1A0000A",
		000573 => x"E3A01002",
		000574 => x"E3A02001",
		000575 => x"EBFFFF13",
		000576 => x"E3A01002",
		000577 => x"E1A0000A",
		000578 => x"EBFFFF49",
		000579 => x"E21010FF",
		000580 => x"11A05001",
		000581 => x"13A06000",
		000582 => x"1AFFFFB0",
		000583 => x"E59F066C",
		000584 => x"EBFFFEFC",
		000585 => x"EAFFFFA5",
		000586 => x"E3A04033",
		000587 => x"E28DA007",
		000588 => x"EAFFFFA4",
		000589 => x"E3540066",
		000590 => x"0A00002A",
		000591 => x"DA0000A4",
		000592 => x"E3540068",
		000593 => x"0A000106",
		000594 => x"E3540072",
		000595 => x"1A00007A",
		000596 => x"E1A00004",
		000597 => x"EBFFFE1E",
		000598 => x"E3A006FF",
		000599 => x"E280F20F",
		000600 => x"EAFFFFFE",
		000601 => x"E1A00004",
		000602 => x"EBFFFE19",
		000603 => x"E59F0618",
		000604 => x"EBFFFEE8",
		000605 => x"E1A0000A",
		000606 => x"E3A01002",
		000607 => x"E3A02001",
		000608 => x"EBFFFEF2",
		000609 => x"E1A0000A",
		000610 => x"E3A01002",
		000611 => x"EBFFFF28",
		000612 => x"E21080FF",
		000613 => x"1A00009B",
		000614 => x"E59F05F4",
		000615 => x"EBFFFEDD",
		000616 => x"EAFFFF86",
		000617 => x"E1A00004",
		000618 => x"EBFFFE09",
		000619 => x"E59F05E4",
		000620 => x"EBFFFED8",
		000621 => x"E1A0000A",
		000622 => x"E3A01004",
		000623 => x"E3A02000",
		000624 => x"EBFFFEE2",
		000625 => x"E5DD3007",
		000626 => x"E3530053",
		000627 => x"1A000002",
		000628 => x"E5DD3008",
		000629 => x"E353004D",
		000630 => x"0A00010C",
		000631 => x"E59F05B8",
		000632 => x"EBFFFECC",
		000633 => x"EAFFFF75",
		000634 => x"E1A00004",
		000635 => x"EBFFFDF8",
		000636 => x"E59F05A8",
		000637 => x"EBFFFEC7",
		000638 => x"E59F05A4",
		000639 => x"EBFFFEC5",
		000640 => x"EAFFFF6E",
		000641 => x"E5DD3009",
		000642 => x"E3530042",
		000643 => x"1AFFFF99",
		000644 => x"E3500052",
		000645 => x"1AFFFF97",
		000646 => x"E1A01005",
		000647 => x"E3A02004",
		000648 => x"E2433040",
		000649 => x"E2800020",
		000650 => x"E58D4000",
		000651 => x"EBFFFE24",
		000652 => x"E1A01005",
		000653 => x"E5CD0007",
		000654 => x"E3A02005",
		000655 => x"E3A03002",
		000656 => x"E3A00072",
		000657 => x"E58D4000",
		000658 => x"EBFFFE1D",
		000659 => x"E1A01005",
		000660 => x"E5CD0008",
		000661 => x"E3A02006",
		000662 => x"E3A03002",
		000663 => x"E3A00072",
		000664 => x"E58D4000",
		000665 => x"EBFFFE16",
		000666 => x"E1A01005",
		000667 => x"E5CD0009",
		000668 => x"E3A02007",
		000669 => x"E3A03002",
		000670 => x"E3A00072",
		000671 => x"E58D4000",
		000672 => x"EBFFFE0F",
		000673 => x"E5CD000A",
		000674 => x"E1A0000A",
		000675 => x"EBFFFF06",
		000676 => x"E2907004",
		000677 => x"0A000021",
		000678 => x"E1A06004",
		000679 => x"E2842008",
		000680 => x"E1A01005",
		000681 => x"E3A03002",
		000682 => x"E3A00072",
		000683 => x"E58D6000",
		000684 => x"EBFFFE03",
		000685 => x"E2842009",
		000686 => x"E5CD0007",
		000687 => x"E1A01005",
		000688 => x"E3A03002",
		000689 => x"E3A00072",
		000690 => x"E58D6000",
		000691 => x"EBFFFDFC",
		000692 => x"E284200A",
		000693 => x"E5CD0008",
		000694 => x"E1A01005",
		000695 => x"E3A03002",
		000696 => x"E3A00072",
		000697 => x"E58D6000",
		000698 => x"EBFFFDF5",
		000699 => x"E284200B",
		000700 => x"E5CD0009",
		000701 => x"E1A01005",
		000702 => x"E3A03002",
		000703 => x"E3A00072",
		000704 => x"E58D6000",
		000705 => x"EBFFFDEE",
		000706 => x"E5CD000A",
		000707 => x"E1A0000A",
		000708 => x"EBFFFEE5",
		000709 => x"E4840004",
		000710 => x"E1540007",
		000711 => x"1AFFFFDE",
		000712 => x"E59F0480",
		000713 => x"EBFFFE7B",
		000714 => x"EAFFFF56",
		000715 => x"E3740001",
		000716 => x"0AFFFF22",
		000717 => x"E3540030",
		000718 => x"0A000004",
		000719 => x"E20400FF",
		000720 => x"EBFFFDA3",
		000721 => x"E59F0460",
		000722 => x"EBFFFE72",
		000723 => x"EAFFFF1B",
		000724 => x"E1A00004",
		000725 => x"EBFFFD9E",
		000726 => x"EAFFFF4A",
		000727 => x"E1A00004",
		000728 => x"EBFFFD9B",
		000729 => x"E59F0444",
		000730 => x"EBFFFE6A",
		000731 => x"EBFFFD92",
		000732 => x"E3700001",
		000733 => x"0AFFFFFC",
		000734 => x"EBFFFD8F",
		000735 => x"E3700001",
		000736 => x"1AFFFFFC",
		000737 => x"E3A05000",
		000738 => x"EA000001",
		000739 => x"E3550902",
		000740 => x"0A00000C",
		000741 => x"E5954000",
		000742 => x"E1A00C24",
		000743 => x"EBFFFD8C",
		000744 => x"E1A00824",
		000745 => x"EBFFFD8A",
		000746 => x"E1A00424",
		000747 => x"EBFFFD88",
		000748 => x"E1A00004",
		000749 => x"EBFFFD86",
		000750 => x"EBFFFD7F",
		000751 => x"E3700001",
		000752 => x"E2855004",
		000753 => x"0AFFFFF0",
		000754 => x"E59F03E4",
		000755 => x"EBFFFE51",
		000756 => x"EAFFFEFA",
		000757 => x"E3540035",
		000758 => x"0A0000A9",
		000759 => x"E3540061",
		000760 => x"1AFFFFD5",
		000761 => x"E1A00004",
		000762 => x"EBFFFD79",
		000763 => x"E59F03C4",
		000764 => x"EBFFFE48",
		000765 => x"E59F03C0",
		000766 => x"EBFFFE46",
		000767 => x"E59F03BC",
		000768 => x"EBFFFE44",
		000769 => x"EAFFFEED",
		000770 => x"E59F03B4",
		000771 => x"EBFFFE41",
		000772 => x"E1A0000A",
		000773 => x"E3A01004",
		000774 => x"E3A02000",
		000775 => x"EBFFFE4B",
		000776 => x"E5DD3007",
		000777 => x"E3530053",
		000778 => x"1A000002",
		000779 => x"E5DD2008",
		000780 => x"E352004D",
		000781 => x"0A000004",
		000782 => x"E59F0388",
		000783 => x"EBFFFE35",
		000784 => x"E59F0384",
		000785 => x"EBFFFE33",
		000786 => x"EAFFFEDC",
		000787 => x"E5DD1009",
		000788 => x"E3510042",
		000789 => x"1AFFFFF7",
		000790 => x"E5DD000A",
		000791 => x"E3500052",
		000792 => x"1AFFFFF4",
		000793 => x"E3A04000",
		000794 => x"E5C43000",
		000795 => x"E1A00000",
		000796 => x"E5C42001",
		000797 => x"E1A00000",
		000798 => x"E5C41002",
		000799 => x"E1A00000",
		000800 => x"E5C40003",
		000801 => x"E1A00000",
		000802 => x"E241103E",
		000803 => x"E1A0000A",
		000804 => x"E1A02004",
		000805 => x"EBFFFE2D",
		000806 => x"E5DD3007",
		000807 => x"E5C43004",
		000808 => x"E5DD2008",
		000809 => x"E5C42005",
		000810 => x"E5DD3009",
		000811 => x"E5C43006",
		000812 => x"E5DD200A",
		000813 => x"E1A0000A",
		000814 => x"E5C42007",
		000815 => x"EBFFFE7A",
		000816 => x"E3A03CFF",
		000817 => x"E28330FC",
		000818 => x"E1500003",
		000819 => x"E1A05000",
		000820 => x"8A000095",
		000821 => x"E3700004",
		000822 => x"12844008",
		000823 => x"1280600B",
		000824 => x"0A000006",
		000825 => x"EBFFFD34",
		000826 => x"E3700001",
		000827 => x"0AFFFFFC",
		000828 => x"E1560004",
		000829 => x"E5C40000",
		000830 => x"E2844001",
		000831 => x"1AFFFFF8",
		000832 => x"E59F02C8",
		000833 => x"EBFFFE03",
		000834 => x"E59F02C4",
		000835 => x"EBFFFE01",
		000836 => x"E375000C",
		000837 => x"0A00000F",
		000838 => x"E3A04000",
		000839 => x"E285700C",
		000840 => x"E1A06004",
		000841 => x"E5D45000",
		000842 => x"E3A00077",
		000843 => x"E1A01008",
		000844 => x"E1A02006",
		000845 => x"E3A03002",
		000846 => x"E58D5000",
		000847 => x"EBFFFD60",
		000848 => x"E3500000",
		000849 => x"1AFFFFF7",
		000850 => x"E2844001",
		000851 => x"E1540007",
		000852 => x"E1A06004",
		000853 => x"1AFFFFF2",
		000854 => x"E59F0278",
		000855 => x"EBFFFDED",
		000856 => x"EAFFFFB6",
		000857 => x"E1A00004",
		000858 => x"EBFFFD19",
		000859 => x"E59F0268",
		000860 => x"EBFFFDE8",
		000861 => x"E59F0264",
		000862 => x"EBFFFDE6",
		000863 => x"E59F0260",
		000864 => x"EBFFFDE4",
		000865 => x"E59F025C",
		000866 => x"EBFFFDE2",
		000867 => x"E59F0258",
		000868 => x"EBFFFDE0",
		000869 => x"E59F0254",
		000870 => x"EBFFFDDE",
		000871 => x"E59F0250",
		000872 => x"EBFFFDDC",
		000873 => x"E59F024C",
		000874 => x"EBFFFDDA",
		000875 => x"E59F0248",
		000876 => x"EBFFFDD8",
		000877 => x"E59F0244",
		000878 => x"EBFFFDD6",
		000879 => x"E59F0240",
		000880 => x"EBFFFDD4",
		000881 => x"E59F023C",
		000882 => x"EBFFFDD2",
		000883 => x"E59F0238",
		000884 => x"EBFFFDD0",
		000885 => x"E59F0234",
		000886 => x"EBFFFDCE",
		000887 => x"E59F0230",
		000888 => x"EBFFFDCC",
		000889 => x"E59F022C",
		000890 => x"EBFFFDCA",
		000891 => x"E59F0228",
		000892 => x"EBFFFDC8",
		000893 => x"E59F0224",
		000894 => x"EBFFFDC6",
		000895 => x"E59F0220",
		000896 => x"EBFFFDC4",
		000897 => x"E59F021C",
		000898 => x"EBFFFDC2",
		000899 => x"EAFFFE6B",
		000900 => x"E5DD3009",
		000901 => x"E3530042",
		000902 => x"1AFFFEEF",
		000903 => x"E5DD300A",
		000904 => x"E3530052",
		000905 => x"1AFFFEEC",
		000906 => x"E3A01004",
		000907 => x"E3A02000",
		000908 => x"E1A0000A",
		000909 => x"EBFFFDC5",
		000910 => x"E1A0000A",
		000911 => x"EBFFFE1A",
		000912 => x"E3A03C7F",
		000913 => x"E28330F8",
		000914 => x"E1500003",
		000915 => x"8A000036",
		000916 => x"E2905004",
		000917 => x"0AFFFE8B",
		000918 => x"E3A04000",
		000919 => x"E3A01004",
		000920 => x"E3A02000",
		000921 => x"E1A0000A",
		000922 => x"EBFFFDB8",
		000923 => x"E1A0000A",
		000924 => x"EBFFFE0D",
		000925 => x"E4840004",
		000926 => x"E1540005",
		000927 => x"1AFFFFF6",
		000928 => x"EAFFFE80",
		000929 => x"E1A00004",
		000930 => x"EBFFFCD1",
		000931 => x"E59F0198",
		000932 => x"EBFFFDA0",
		000933 => x"E1A0000A",
		000934 => x"E3A01002",
		000935 => x"E3A02001",
		000936 => x"EBFFFDAA",
		000937 => x"E1A0000A",
		000938 => x"E3A01002",
		000939 => x"EBFFFDE0",
		000940 => x"E21060FF",
		000941 => x"0AFFFE98",
		000942 => x"E59F0170",
		000943 => x"EBFFFD95",
		000944 => x"E59F016C",
		000945 => x"EBFFFD93",
		000946 => x"EBFFFCBB",
		000947 => x"E3700001",
		000948 => x"0AFFFFFC",
		000949 => x"EBFFFCB8",
		000950 => x"E3700001",
		000951 => x"1AFFFFFC",
		000952 => x"E3A05000",
		000953 => x"EA000001",
		000954 => x"E3540000",
		000955 => x"AA000011",
		000956 => x"E3A0C000",
		000957 => x"E1A02005",
		000958 => x"E1A01006",
		000959 => x"E3A03002",
		000960 => x"E3A00072",
		000961 => x"E58DC000",
		000962 => x"EBFFFCED",
		000963 => x"E1A04000",
		000964 => x"EBFFFCA9",
		000965 => x"E3700001",
		000966 => x"E1A00004",
		000967 => x"0AFFFFF1",
		000968 => x"E59F0110",
		000969 => x"EBFFFD7B",
		000970 => x"EAFFFF26",
		000971 => x"E59F0108",
		000972 => x"EBFFFD78",
		000973 => x"EAFFFE21",
		000974 => x"EBFFFCA5",
		000975 => x"E3A03801",
		000976 => x"E2855001",
		000977 => x"E2433001",
		000978 => x"E1550003",
		000979 => x"1AFFFFE7",
		000980 => x"EAFFFF1C",
		000981 => x"FFF01040",
		000982 => x"FFF0108C",
		000983 => x"FFF010D4",
		000984 => x"FFF0111C",
		000985 => x"FFF01164",
		000986 => x"FFF011AC",
		000987 => x"FFF011F4",
		000988 => x"FFF01260",
		000989 => x"FFF01298",
		000990 => x"FFF012FC",
		000991 => x"FFF01360",
		000992 => x"FFF01538",
		000993 => x"FFF0159C",
		000994 => x"FFF01CA0",
		000995 => x"FFF014DC",
		000996 => x"FFF01518",
		000997 => x"FFF015C8",
		000998 => x"FFF013B0",
		000999 => x"FFF01448",
		001000 => x"FFF01C24",
		001001 => x"FFF01C54",
		001002 => x"FFF01588",
		001003 => x"FFF01C7C",
		001004 => x"FFF01470",
		001005 => x"FFF014B8",
		001006 => x"FFF01778",
		001007 => x"FFF017AC",
		001008 => x"FFF01818",
		001009 => x"FFF015E8",
		001010 => x"FFF01690",
		001011 => x"FFF01C70",
		001012 => x"FFF01648",
		001013 => x"FFF01660",
		001014 => x"FFF01680",
		001015 => x"FFF0185C",
		001016 => x"FFF01878",
		001017 => x"FFF01898",
		001018 => x"FFF018D8",
		001019 => x"FFF0190C",
		001020 => x"FFF01948",
		001021 => x"FFF01984",
		001022 => x"FFF019A8",
		001023 => x"FFF019E4",
		001024 => x"FFF01A00",
		001025 => x"FFF01A18",
		001026 => x"FFF01A60",
		001027 => x"FFF01AA0",
		001028 => x"FFF01AD8",
		001029 => x"FFF01AFC",
		001030 => x"FFF01B40",
		001031 => x"FFF01B80",
		001032 => x"FFF01BAC",
		001033 => x"FFF01BD8",
		001034 => x"FFF01BFC",
		001035 => x"FFF016B4",
		001036 => x"FFF016F0",
		001037 => x"FFF01730",
		001038 => x"FFF01CC4",
		001039 => x"FFF01424",
		001040 => x"0D0A0D0A",
		001041 => x"0D0A2B2D",
		001042 => x"2D2D2D2D",
		001043 => x"2D2D2D2D",
		001044 => x"2D2D2D2D",
		001045 => x"2D2D2D2D",
		001046 => x"2D2D2D2D",
		001047 => x"2D2D2D2D",
		001048 => x"2D2D2D2D",
		001049 => x"2D2D2D2D",
		001050 => x"2D2D2D2D",
		001051 => x"2D2D2D2D",
		001052 => x"2D2D2D2D",
		001053 => x"2D2D2D2D",
		001054 => x"2D2D2D2D",
		001055 => x"2D2D2D2D",
		001056 => x"2D2D2D2D",
		001057 => x"2D2D2D2B",
		001058 => x"0D0A0000",
		001059 => x"7C202020",
		001060 => x"203C3C3C",
		001061 => x"2053544F",
		001062 => x"524D2043",
		001063 => x"6F726520",
		001064 => x"50726F63",
		001065 => x"6573736F",
		001066 => x"72205379",
		001067 => x"7374656D",
		001068 => x"202D2042",
		001069 => x"79205374",
		001070 => x"65706861",
		001071 => x"6E204E6F",
		001072 => x"6C74696E",
		001073 => x"67203E3E",
		001074 => x"3E202020",
		001075 => x"207C0D0A",
		001076 => x"00000000",
		001077 => x"2B2D2D2D",
		001078 => x"2D2D2D2D",
		001079 => x"2D2D2D2D",
		001080 => x"2D2D2D2D",
		001081 => x"2D2D2D2D",
		001082 => x"2D2D2D2D",
		001083 => x"2D2D2D2D",
		001084 => x"2D2D2D2D",
		001085 => x"2D2D2D2D",
		001086 => x"2D2D2D2D",
		001087 => x"2D2D2D2D",
		001088 => x"2D2D2D2D",
		001089 => x"2D2D2D2D",
		001090 => x"2D2D2D2D",
		001091 => x"2D2D2D2D",
		001092 => x"2D2D2D2D",
		001093 => x"2D2B0D0A",
		001094 => x"00000000",
		001095 => x"7C202020",
		001096 => x"20202020",
		001097 => x"2020426F",
		001098 => x"6F746C6F",
		001099 => x"61646572",
		001100 => x"20666F72",
		001101 => x"2053544F",
		001102 => x"524D2053",
		001103 => x"6F432020",
		001104 => x"20566572",
		001105 => x"73696F6E",
		001106 => x"3A203230",
		001107 => x"31323035",
		001108 => x"32342D43",
		001109 => x"20202020",
		001110 => x"20202020",
		001111 => x"207C0D0A",
		001112 => x"00000000",
		001113 => x"7C202020",
		001114 => x"20202020",
		001115 => x"20202020",
		001116 => x"20202020",
		001117 => x"436F6E74",
		001118 => x"6163743A",
		001119 => x"2073746E",
		001120 => x"6F6C7469",
		001121 => x"6E674067",
		001122 => x"6F6F676C",
		001123 => x"656D6169",
		001124 => x"6C2E636F",
		001125 => x"6D202020",
		001126 => x"20202020",
		001127 => x"20202020",
		001128 => x"20202020",
		001129 => x"207C0D0A",
		001130 => x"00000000",
		001131 => x"2B2D2D2D",
		001132 => x"2D2D2D2D",
		001133 => x"2D2D2D2D",
		001134 => x"2D2D2D2D",
		001135 => x"2D2D2D2D",
		001136 => x"2D2D2D2D",
		001137 => x"2D2D2D2D",
		001138 => x"2D2D2D2D",
		001139 => x"2D2D2D2D",
		001140 => x"2D2D2D2D",
		001141 => x"2D2D2D2D",
		001142 => x"2D2D2D2D",
		001143 => x"2D2D2D2D",
		001144 => x"2D2D2D2D",
		001145 => x"2D2D2D2D",
		001146 => x"2D2D2D2D",
		001147 => x"2D2B0D0A",
		001148 => x"0D0A0000",
		001149 => x"203C2057",
		001150 => x"656C636F",
		001151 => x"6D652074",
		001152 => x"6F207468",
		001153 => x"65205354",
		001154 => x"4F524D20",
		001155 => x"536F4320",
		001156 => x"626F6F74",
		001157 => x"6C6F6164",
		001158 => x"65722063",
		001159 => x"6F6E736F",
		001160 => x"6C652120",
		001161 => x"3E0D0A20",
		001162 => x"3C205365",
		001163 => x"6C656374",
		001164 => x"20616E20",
		001165 => x"6F706572",
		001166 => x"6174696F",
		001167 => x"6E206672",
		001168 => x"6F6D2074",
		001169 => x"6865206D",
		001170 => x"656E7520",
		001171 => x"62656C6F",
		001172 => x"77206F72",
		001173 => x"20707265",
		001174 => x"7373203E",
		001175 => x"0D0A0000",
		001176 => x"203C2074",
		001177 => x"68652062",
		001178 => x"6F6F7420",
		001179 => x"6B657920",
		001180 => x"666F7220",
		001181 => x"696D6D65",
		001182 => x"64696174",
		001183 => x"65206170",
		001184 => x"706C6963",
		001185 => x"6174696F",
		001186 => x"6E207374",
		001187 => x"6172742E",
		001188 => x"203E0D0A",
		001189 => x"0D0A0000",
		001190 => x"2030202D",
		001191 => x"20626F6F",
		001192 => x"74206672",
		001193 => x"6F6D2063",
		001194 => x"6F726520",
		001195 => x"52414D20",
		001196 => x"28737461",
		001197 => x"72742061",
		001198 => x"70706C69",
		001199 => x"63617469",
		001200 => x"6F6E290D",
		001201 => x"0A203120",
		001202 => x"2D207072",
		001203 => x"6F677261",
		001204 => x"6D20636F",
		001205 => x"72652052",
		001206 => x"414D2076",
		001207 => x"69612055",
		001208 => x"4152545F",
		001209 => x"300D0A20",
		001210 => x"32202D20",
		001211 => x"636F7265",
		001212 => x"2052414D",
		001213 => x"2064756D",
		001214 => x"700D0A00",
		001215 => x"2033202D",
		001216 => x"20626F6F",
		001217 => x"74206672",
		001218 => x"6F6D2049",
		001219 => x"32432045",
		001220 => x"4550524F",
		001221 => x"4D0D0A20",
		001222 => x"34202D20",
		001223 => x"70726F67",
		001224 => x"72616D20",
		001225 => x"49324320",
		001226 => x"45455052",
		001227 => x"4F4D2076",
		001228 => x"69612055",
		001229 => x"4152545F",
		001230 => x"300D0A20",
		001231 => x"35202D20",
		001232 => x"73686F77",
		001233 => x"20636F6E",
		001234 => x"74656E74",
		001235 => x"206F6620",
		001236 => x"49324320",
		001237 => x"45455052",
		001238 => x"4F4D0D0A",
		001239 => x"00000000",
		001240 => x"2061202D",
		001241 => x"20617574",
		001242 => x"6F6D6174",
		001243 => x"69632062",
		001244 => x"6F6F7420",
		001245 => x"636F6E66",
		001246 => x"69677572",
		001247 => x"6174696F",
		001248 => x"6E0D0A20",
		001249 => x"68202D20",
		001250 => x"68656C70",
		001251 => x"0D0A2072",
		001252 => x"202D2072",
		001253 => x"65737461",
		001254 => x"72742073",
		001255 => x"79737465",
		001256 => x"6D0D0A0D",
		001257 => x"0A53656C",
		001258 => x"6563743A",
		001259 => x"20000000",
		001260 => x"0D0A0D0A",
		001261 => x"4170706C",
		001262 => x"69636174",
		001263 => x"696F6E20",
		001264 => x"77696C6C",
		001265 => x"20737461",
		001266 => x"72742061",
		001267 => x"75746F6D",
		001268 => x"61746963",
		001269 => x"616C6C79",
		001270 => x"20616674",
		001271 => x"65722064",
		001272 => x"6F776E6C",
		001273 => x"6F61642E",
		001274 => x"0D0A2D3E",
		001275 => x"20576169",
		001276 => x"74696E67",
		001277 => x"20666F72",
		001278 => x"20277374",
		001279 => x"6F726D5F",
		001280 => x"70726F67",
		001281 => x"72616D2E",
		001282 => x"62696E27",
		001283 => x"20696E20",
		001284 => x"62797465",
		001285 => x"2D737472",
		001286 => x"65616D20",
		001287 => x"6D6F6465",
		001288 => x"2E2E2E00",
		001289 => x"20455252",
		001290 => x"4F522120",
		001291 => x"50726F67",
		001292 => x"72616D20",
		001293 => x"66696C65",
		001294 => x"20746F6F",
		001295 => x"20626967",
		001296 => x"210D0A0D",
		001297 => x"0A000000",
		001298 => x"20496E76",
		001299 => x"616C6964",
		001300 => x"2070726F",
		001301 => x"6772616D",
		001302 => x"6D696E67",
		001303 => x"2066696C",
		001304 => x"65210D0A",
		001305 => x"0D0A5365",
		001306 => x"6C656374",
		001307 => x"3A200000",
		001308 => x"0D0A0D0A",
		001309 => x"41626F72",
		001310 => x"74206475",
		001311 => x"6D70696E",
		001312 => x"67206279",
		001313 => x"20707265",
		001314 => x"7373696E",
		001315 => x"6720616E",
		001316 => x"79206B65",
		001317 => x"792E0D0A",
		001318 => x"50726573",
		001319 => x"7320616E",
		001320 => x"79206B65",
		001321 => x"7920746F",
		001322 => x"20636F6E",
		001323 => x"74696E75",
		001324 => x"652E0D0A",
		001325 => x"0D0A0000",
		001326 => x"0D0A0D0A",
		001327 => x"44756D70",
		001328 => x"696E6720",
		001329 => x"636F6D70",
		001330 => x"6C657465",
		001331 => x"642E0D0A",
		001332 => x"0D0A5365",
		001333 => x"6C656374",
		001334 => x"3A200000",
		001335 => x"0D0A0D0A",
		001336 => x"456E7465",
		001337 => x"72206465",
		001338 => x"76696365",
		001339 => x"20616464",
		001340 => x"72657373",
		001341 => x"20283278",
		001342 => x"20686578",
		001343 => x"5F636861",
		001344 => x"72732C20",
		001345 => x"73657420",
		001346 => x"4C534220",
		001347 => x"746F2027",
		001348 => x"3027293A",
		001349 => x"20000000",
		001350 => x"20496E76",
		001351 => x"616C6964",
		001352 => x"20616464",
		001353 => x"72657373",
		001354 => x"210D0A0D",
		001355 => x"0A53656C",
		001356 => x"6563743A",
		001357 => x"20000000",
		001358 => x"0D0A4170",
		001359 => x"706C6963",
		001360 => x"6174696F",
		001361 => x"6E207769",
		001362 => x"6C6C2073",
		001363 => x"74617274",
		001364 => x"20617574",
		001365 => x"6F6D6174",
		001366 => x"6963616C",
		001367 => x"6C792061",
		001368 => x"66746572",
		001369 => x"2075706C",
		001370 => x"6F61642E",
		001371 => x"0D0A2D3E",
		001372 => x"204C6F61",
		001373 => x"64696E67",
		001374 => x"20626F6F",
		001375 => x"7420696D",
		001376 => x"6167652E",
		001377 => x"2E2E0000",
		001378 => x"2055706C",
		001379 => x"6F616420",
		001380 => x"636F6D70",
		001381 => x"6C657465",
		001382 => x"0D0A0000",
		001383 => x"20496E76",
		001384 => x"616C6964",
		001385 => x"20626F6F",
		001386 => x"74206465",
		001387 => x"76696365",
		001388 => x"206F7220",
		001389 => x"66696C65",
		001390 => x"210D0A0D",
		001391 => x"0A53656C",
		001392 => x"6563743A",
		001393 => x"20000000",
		001394 => x"0D0A496E",
		001395 => x"76616C69",
		001396 => x"64206164",
		001397 => x"64726573",
		001398 => x"73210D0A",
		001399 => x"0D0A5365",
		001400 => x"6C656374",
		001401 => x"3A200000",
		001402 => x"0D0A4461",
		001403 => x"74612077",
		001404 => x"696C6C20",
		001405 => x"6F766572",
		001406 => x"77726974",
		001407 => x"65205241",
		001408 => x"4D20636F",
		001409 => x"6E74656E",
		001410 => x"74210D0A",
		001411 => x"2D3E2057",
		001412 => x"61697469",
		001413 => x"6E672066",
		001414 => x"6F722027",
		001415 => x"73746F72",
		001416 => x"6D5F7072",
		001417 => x"6F677261",
		001418 => x"6D2E6269",
		001419 => x"6E272069",
		001420 => x"6E206279",
		001421 => x"74652D73",
		001422 => x"74726561",
		001423 => x"6D206D6F",
		001424 => x"64652E2E",
		001425 => x"2E000000",
		001426 => x"20446F77",
		001427 => x"6E6C6F61",
		001428 => x"6420636F",
		001429 => x"6D706C65",
		001430 => x"7465640D",
		001431 => x"0A000000",
		001432 => x"57726974",
		001433 => x"696E6720",
		001434 => x"62756666",
		001435 => x"65722074",
		001436 => x"6F206932",
		001437 => x"63204545",
		001438 => x"50524F4D",
		001439 => x"2E2E2E00",
		001440 => x"20436F6D",
		001441 => x"706C6574",
		001442 => x"65640D0A",
		001443 => x"0D0A0000",
		001444 => x"20496E76",
		001445 => x"616C6964",
		001446 => x"20626F6F",
		001447 => x"74206465",
		001448 => x"76696365",
		001449 => x"206F7220",
		001450 => x"66696C65",
		001451 => x"210D0A0D",
		001452 => x"0A000000",
		001453 => x"0D0A0D0A",
		001454 => x"456E7465",
		001455 => x"72206465",
		001456 => x"76696365",
		001457 => x"20616464",
		001458 => x"72657373",
		001459 => x"20283220",
		001460 => x"6865782D",
		001461 => x"63686172",
		001462 => x"732C2073",
		001463 => x"6574204C",
		001464 => x"53422074",
		001465 => x"6F202730",
		001466 => x"27293A20",
		001467 => x"00000000",
		001468 => x"0D0A0D0A",
		001469 => x"41626F72",
		001470 => x"74206475",
		001471 => x"6D70696E",
		001472 => x"67206279",
		001473 => x"20707265",
		001474 => x"7373696E",
		001475 => x"6720616E",
		001476 => x"79206B65",
		001477 => x"792E2049",
		001478 => x"66206E6F",
		001479 => x"20646174",
		001480 => x"61206973",
		001481 => x"2073686F",
		001482 => x"776E2C0D",
		001483 => x"0A000000",
		001484 => x"74686520",
		001485 => x"73656C65",
		001486 => x"63746564",
		001487 => x"20646576",
		001488 => x"69636520",
		001489 => x"6973206E",
		001490 => x"6F742072",
		001491 => x"6573706F",
		001492 => x"6E64696E",
		001493 => x"672E2050",
		001494 => x"72657373",
		001495 => x"20616E79",
		001496 => x"206B6579",
		001497 => x"20746F20",
		001498 => x"636F6E74",
		001499 => x"696E7565",
		001500 => x"2E0D0A0D",
		001501 => x"0A000000",
		001502 => x"0D0A0D0A",
		001503 => x"4175746F",
		001504 => x"6D617469",
		001505 => x"6320626F",
		001506 => x"6F742063",
		001507 => x"6F6E6669",
		001508 => x"67757261",
		001509 => x"74696F6E",
		001510 => x"20666F72",
		001511 => x"20706F77",
		001512 => x"65722D75",
		001513 => x"703A0D0A",
		001514 => x"00000000",
		001515 => x"5B333231",
		001516 => x"305D2063",
		001517 => x"6F6E6669",
		001518 => x"67757261",
		001519 => x"74696F6E",
		001520 => x"20444950",
		001521 => x"20737769",
		001522 => x"7463680D",
		001523 => x"0A203030",
		001524 => x"3030202D",
		001525 => x"20537461",
		001526 => x"72742062",
		001527 => x"6F6F746C",
		001528 => x"6F616465",
		001529 => x"7220636F",
		001530 => x"6E736F6C",
		001531 => x"650D0A20",
		001532 => x"30303031",
		001533 => x"202D2041",
		001534 => x"75746F6D",
		001535 => x"61746963",
		001536 => x"20626F6F",
		001537 => x"74206672",
		001538 => x"6F6D2063",
		001539 => x"6F726520",
		001540 => x"52414D0D",
		001541 => x"0A000000",
		001542 => x"20303031",
		001543 => x"30202D20",
		001544 => x"4175746F",
		001545 => x"6D617469",
		001546 => x"6320626F",
		001547 => x"6F742066",
		001548 => x"726F6D20",
		001549 => x"49324320",
		001550 => x"45455052",
		001551 => x"4F4D2028",
		001552 => x"41646472",
		001553 => x"65737320",
		001554 => x"30784130",
		001555 => x"290D0A0D",
		001556 => x"0A53656C",
		001557 => x"6563743A",
		001558 => x"20000000",
		001559 => x"0D0A0D0A",
		001560 => x"53544F52",
		001561 => x"4D20536F",
		001562 => x"4320626F",
		001563 => x"6F746C6F",
		001564 => x"61646572",
		001565 => x"0D0A0000",
		001566 => x"2730273A",
		001567 => x"20457865",
		001568 => x"63757465",
		001569 => x"2070726F",
		001570 => x"6772616D",
		001571 => x"20696E20",
		001572 => x"52414D2E",
		001573 => x"0D0A0000",
		001574 => x"2731273A",
		001575 => x"20577269",
		001576 => x"74652027",
		001577 => x"73746F72",
		001578 => x"6D5F7072",
		001579 => x"6F677261",
		001580 => x"6D2E6269",
		001581 => x"6E272074",
		001582 => x"6F207468",
		001583 => x"6520636F",
		001584 => x"72652773",
		001585 => x"2052414D",
		001586 => x"20766961",
		001587 => x"20554152",
		001588 => x"542E0D0A",
		001589 => x"00000000",
		001590 => x"2732273A",
		001591 => x"20507269",
		001592 => x"6E742063",
		001593 => x"75727265",
		001594 => x"6E742063",
		001595 => x"6F6E7465",
		001596 => x"6E74206F",
		001597 => x"6620636F",
		001598 => x"6D706C65",
		001599 => x"74652063",
		001600 => x"6F726520",
		001601 => x"52414D2E",
		001602 => x"0D0A0000",
		001603 => x"2733273A",
		001604 => x"204C6F61",
		001605 => x"6420626F",
		001606 => x"6F742069",
		001607 => x"6D616765",
		001608 => x"2066726F",
		001609 => x"6D204545",
		001610 => x"50524F4D",
		001611 => x"20616E64",
		001612 => x"20737461",
		001613 => x"72742061",
		001614 => x"70706C69",
		001615 => x"63617469",
		001616 => x"6F6E2E0D",
		001617 => x"0A000000",
		001618 => x"2734273A",
		001619 => x"20577269",
		001620 => x"74652027",
		001621 => x"73746F72",
		001622 => x"6D5F7072",
		001623 => x"6F677261",
		001624 => x"6D2E6269",
		001625 => x"6E272074",
		001626 => x"6F204932",
		001627 => x"43204545",
		001628 => x"50524F4D",
		001629 => x"20766961",
		001630 => x"20554152",
		001631 => x"542E0D0A",
		001632 => x"00000000",
		001633 => x"2735273A",
		001634 => x"20507269",
		001635 => x"6E742063",
		001636 => x"6F6E7465",
		001637 => x"6E74206F",
		001638 => x"66204932",
		001639 => x"43204545",
		001640 => x"50524F4D",
		001641 => x"2E0D0A00",
		001642 => x"2761273A",
		001643 => x"2053686F",
		001644 => x"77204449",
		001645 => x"50207377",
		001646 => x"69746368",
		001647 => x"20636F6E",
		001648 => x"66696775",
		001649 => x"72617469",
		001650 => x"6F6E7320",
		001651 => x"666F7220",
		001652 => x"6175746F",
		001653 => x"6D617469",
		001654 => x"6320626F",
		001655 => x"6F742E0D",
		001656 => x"0A000000",
		001657 => x"2768273A",
		001658 => x"2053686F",
		001659 => x"77207468",
		001660 => x"69732073",
		001661 => x"63726565",
		001662 => x"6E2E0D0A",
		001663 => x"00000000",
		001664 => x"2772273A",
		001665 => x"20526573",
		001666 => x"65742073",
		001667 => x"79737465",
		001668 => x"6D2E0D0A",
		001669 => x"0D0A0000",
		001670 => x"426F6F74",
		001671 => x"20454550",
		001672 => x"524F4D3A",
		001673 => x"20323478",
		001674 => x"786E6E6E",
		001675 => x"20286C69",
		001676 => x"6B652032",
		001677 => x"34414136",
		001678 => x"34292C20",
		001679 => x"37206269",
		001680 => x"74206164",
		001681 => x"64726573",
		001682 => x"73202B20",
		001683 => x"646F6E74",
		001684 => x"2D636172",
		001685 => x"65206269",
		001686 => x"742C0D0A",
		001687 => x"00000000",
		001688 => x"636F6E6E",
		001689 => x"65637465",
		001690 => x"6420746F",
		001691 => x"20493243",
		001692 => x"5F434F4E",
		001693 => x"54524F4C",
		001694 => x"4C45525F",
		001695 => x"302C206F",
		001696 => x"70657261",
		001697 => x"74696E67",
		001698 => x"20667265",
		001699 => x"7175656E",
		001700 => x"63792069",
		001701 => x"73203130",
		001702 => x"306B487A",
		001703 => x"2C0D0A00",
		001704 => x"6D617869",
		001705 => x"6D756D20",
		001706 => x"45455052",
		001707 => x"4F4D2073",
		001708 => x"697A6520",
		001709 => x"3D203635",
		001710 => x"35333620",
		001711 => x"62797465",
		001712 => x"203D3E20",
		001713 => x"31362062",
		001714 => x"69742061",
		001715 => x"64647265",
		001716 => x"73736573",
		001717 => x"2C0D0A00",
		001718 => x"66697865",
		001719 => x"6420626F",
		001720 => x"6F742064",
		001721 => x"65766963",
		001722 => x"65206164",
		001723 => x"64726573",
		001724 => x"733A2030",
		001725 => x"7841300D",
		001726 => x"0A0D0A00",
		001727 => x"5465726D",
		001728 => x"696E616C",
		001729 => x"20736574",
		001730 => x"75703A20",
		001731 => x"39363030",
		001732 => x"20626175",
		001733 => x"642C2038",
		001734 => x"20646174",
		001735 => x"61206269",
		001736 => x"74732C20",
		001737 => x"6E6F2070",
		001738 => x"61726974",
		001739 => x"792C2031",
		001740 => x"2073746F",
		001741 => x"70206269",
		001742 => x"740D0A0D",
		001743 => x"0A000000",
		001744 => x"466F7220",
		001745 => x"6D6F7265",
		001746 => x"20696E66",
		001747 => x"6F726D61",
		001748 => x"74696F6E",
		001749 => x"20736565",
		001750 => x"20746865",
		001751 => x"2053544F",
		001752 => x"524D2043",
		001753 => x"6F726520",
		001754 => x"2F205354",
		001755 => x"4F524D20",
		001756 => x"536F4320",
		001757 => x"64617461",
		001758 => x"73686565",
		001759 => x"740D0A00",
		001760 => x"68747470",
		001761 => x"3A2F2F6F",
		001762 => x"70656E63",
		001763 => x"6F726573",
		001764 => x"2E6F7267",
		001765 => x"2F70726F",
		001766 => x"6A656374",
		001767 => x"2C73746F",
		001768 => x"726D5F63",
		001769 => x"6F72650D",
		001770 => x"0A000000",
		001771 => x"68747470",
		001772 => x"3A2F2F6F",
		001773 => x"70656E63",
		001774 => x"6F726573",
		001775 => x"2E6F7267",
		001776 => x"2F70726F",
		001777 => x"6A656374",
		001778 => x"2C73746F",
		001779 => x"726D5F73",
		001780 => x"6F630D0A",
		001781 => x"00000000",
		001782 => x"436F6E74",
		001783 => x"6163743A",
		001784 => x"2073746E",
		001785 => x"6F6C7469",
		001786 => x"6E674067",
		001787 => x"6F6F676C",
		001788 => x"656D6169",
		001789 => x"6C2E636F",
		001790 => x"6D0D0A00",
		001791 => x"28632920",
		001792 => x"32303132",
		001793 => x"20627920",
		001794 => x"53746570",
		001795 => x"68616E20",
		001796 => x"4E6F6C74",
		001797 => x"696E670D",
		001798 => x"0A0D0A53",
		001799 => x"656C6563",
		001800 => x"743A2000",
		001801 => x"0D0A0D0A",
		001802 => x"5765276C",
		001803 => x"6C207365",
		001804 => x"6E642079",
		001805 => x"6F752062",
		001806 => x"61636B20",
		001807 => x"2D20746F",
		001808 => x"20746865",
		001809 => x"20667574",
		001810 => x"75726521",
		001811 => x"2E0D0A0D",
		001812 => x"0A000000",
		001813 => x"202D2044",
		001814 => x"6F63746F",
		001815 => x"7220456D",
		001816 => x"6D657420",
		001817 => x"4C2E2042",
		001818 => x"726F776E",
		001819 => x"0D0A0D0A",
		001820 => x"53656C65",
		001821 => x"63743A20",
		001822 => x"00000000",
		001823 => x"20496E76",
		001824 => x"616C6964",
		001825 => x"206F7065",
		001826 => x"72617469",
		001827 => x"6F6E210D",
		001828 => x"0A547279",
		001829 => x"20616761",
		001830 => x"696E3A20",
		001831 => x"00000000",
		001832 => x"0D0A0D0A",
		001833 => x"2D3E2053",
		001834 => x"74617274",
		001835 => x"696E6720",
		001836 => x"6170706C",
		001837 => x"69636174",
		001838 => x"696F6E2E",
		001839 => x"2E2E0D0A",
		001840 => x"0D0A0000",
		001841 => x"0D0A0D0A",
		001842 => x"41626F72",
		001843 => x"74656421",
		001844 => x"00000000",
		others => x"F0013007"
	);

	--- Init Memory Function ---
	function load_image(IMAGE_ID : string) return BOOT_ROM_TYPE is
		variable TEMP_MEM : BOOT_ROM_TYPE;
	begin
		if (IMAGE_ID = "STORM_SOC_BASIC_BL_32_8") then
			TEMP_MEM := STORM_SOC_BASIC_BL_32_8;
		else
			TEMP_MEM := (others => x"F0013007"); -- no image
		end if;
		return TEMP_MEM;
	end load_image;

	--- ROM Signal ---
	signal BOOT_ROM : BOOT_ROM_TYPE := load_image(INIT_IMAGE_ID);

begin

	-- ROM WB Access ---------------------------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		ROM_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read ---
				if (WB_STB_I = '1') then
					WB_DATA_INT <= BOOT_ROM(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I; -- data is valid one cycle later
				end if;
			end if;
		end process ROM_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else x"00000000";

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;