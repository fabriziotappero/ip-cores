
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package tinycpu is

        type regdatatype is array(15 downto 0) of std_logic_vector(7 downto 0);
        type regwritetype is array(15 downto 0) of std_logic;

end tinycpu;

package body tinycpu is

 
end tinycpu;
