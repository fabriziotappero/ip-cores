-------------------------------------------------------------------------------
--
-- The Port 2 unit.
-- Implements the Port 2 logic.
--
-- $Id: p2-c.vhd 295 2009-04-01 19:32:48Z arniml $
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t48_p2_rtl_c0 of t48_p2 is

  for rtl
  end for;

end t48_p2_rtl_c0;
