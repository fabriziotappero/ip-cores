function Action debug(Bool b, Action a);
  action

  if (b) a;

  endaction
endfunction 