-------------------------------------------------------------------------------
--
-- SNESpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: snespad_ctrl-c.vhd 41 2009-04-01 19:58:04Z arniml $
--
-------------------------------------------------------------------------------

configuration snespad_ctrl_rtl_c0 of snespad_ctrl is

  for rtl
  end for;

end snespad_ctrl_rtl_c0;
