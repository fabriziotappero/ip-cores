000000 => x"cafe",
000001 => x"00bd",
000002 => x"a78d",
000003 => x"524e",
000004 => x"445f",
000005 => x"4e55",
000006 => x"4d42",
000007 => x"4552",
000008 => x"bc0b",
000009 => x"bc04",
000010 => x"bc03",
000011 => x"bc02",
000012 => x"bc01",
000013 => x"be30",
000014 => x"c10e",
000015 => x"c901",
000016 => x"be21",
000017 => x"be2c",
000018 => x"bc00",
000019 => x"c12a",
000020 => x"c901",
000021 => x"be19",
000022 => x"c142",
000023 => x"c901",
000024 => x"be19",
000025 => x"be33",
000026 => x"ec4d",
000027 => x"be22",
000028 => x"c15e",
000029 => x"c901",
000030 => x"be13",
000031 => x"be2d",
000032 => x"d24f",
000033 => x"ec4e",
000034 => x"be1b",
000035 => x"c0b0",
000036 => x"be1e",
000037 => x"c0f8",
000038 => x"be1c",
000039 => x"ee05",
000040 => x"be49",
000041 => x"be14",
000042 => x"ec20",
000043 => x"dc0f",
000044 => x"b9ea",
000045 => x"bdf6",
000046 => x"c5ff",
000047 => x"0270",
000048 => x"bc03",
000049 => x"29b3",
000050 => x"0270",
000051 => x"78a9",
000052 => x"3c90",
000053 => x"c880",
000054 => x"3419",
000055 => x"8003",
000056 => x"be0a",
000057 => x"bdfa",
000058 => x"03c0",
000059 => x"343b",
000060 => x"f707",
000061 => x"0170",
000062 => x"c08d",
000063 => x"be03",
000064 => x"c08a",
000065 => x"03a0",
000066 => x"ec22",
000067 => x"dc05",
000068 => x"b9fe",
000069 => x"ed18",
000070 => x"3470",
000071 => x"ec20",
000072 => x"dc8f",
000073 => x"b9fe",
000074 => x"c800",
000075 => x"3470",
000076 => x"0170",
000077 => x"c200",
000078 => x"c184",
000079 => x"bff8",
000080 => x"c0c7",
000081 => x"1809",
000082 => x"9003",
000083 => x"c0a0",
000084 => x"1001",
000085 => x"c0b0",
000086 => x"1809",
000087 => x"91f8",
000088 => x"c0c6",
000089 => x"1818",
000090 => x"91f5",
000091 => x"c0b9",
000092 => x"1818",
000093 => x"a404",
000094 => x"c0c1",
000095 => x"1809",
000096 => x"a1ef",
000097 => x"0080",
000098 => x"bfe0",
000099 => x"c030",
000100 => x"1090",
000101 => x"c009",
000102 => x"1809",
000103 => x"a402",
000104 => x"0497",
000105 => x"3e42",
000106 => x"3e42",
000107 => x"3e42",
000108 => x"3e42",
000109 => x"2641",
000110 => x"05b9",
000111 => x"85e0",
000112 => x"3420",
000113 => x"0370",
000114 => x"3d42",
000115 => x"3d22",
000116 => x"3d22",
000117 => x"3d22",
000118 => x"be0f",
000119 => x"bfcb",
000120 => x"3d40",
000121 => x"be0c",
000122 => x"bfc8",
000123 => x"3d45",
000124 => x"3d25",
000125 => x"3d25",
000126 => x"3d25",
000127 => x"be06",
000128 => x"bfc2",
000129 => x"0140",
000130 => x"be03",
000131 => x"bfbf",
000132 => x"3460",
000133 => x"c08f",
000134 => x"2121",
000135 => x"c089",
000136 => x"181a",
000137 => x"8803",
000138 => x"c0b0",
000139 => x"bc02",
000140 => x"c0b7",
000141 => x"0892",
000142 => x"3470",
000143 => x"4578",
000144 => x"6365",
000145 => x"7074",
000146 => x"696f",
000147 => x"6e2f",
000148 => x"696e",
000149 => x"7465",
000150 => x"7272",
000151 => x"7570",
000152 => x"7420",
000153 => x"6572",
000154 => x"726f",
000155 => x"7221",
000156 => x"0000",
000157 => x"5261",
000158 => x"6e64",
000159 => x"6f6d",
000160 => x"204e",
000161 => x"756d",
000162 => x"6265",
000163 => x"7220",
000164 => x"4765",
000165 => x"6e65",
000166 => x"7261",
000167 => x"746f",
000168 => x"7200",
000169 => x"456e",
000170 => x"7465",
000171 => x"7220",
000172 => x"4c46",
000173 => x"5352",
000174 => x"2073",
000175 => x"6565",
000176 => x"6420",
000177 => x"2834",
000178 => x"6865",
000179 => x"7829",
000180 => x"3a20",
000181 => x"3078",
000182 => x"0000",
000183 => x"456e",
000184 => x"7465",
000185 => x"7220",
000186 => x"4c46",
000187 => x"5352",
000188 => x"2074",
000189 => x"6170",
000190 => x"7320",
000191 => x"2834",
000192 => x"6865",
000193 => x"7829",
000194 => x"3a20",
000195 => x"3078",
000196 => x"0000",
others => x"0000"