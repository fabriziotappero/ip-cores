library verilog;
use verilog.vl_types.all;
entity scalerTestbench is
    generic(
        BUFFER_SIZE     : integer := 4
    );
end scalerTestbench;
