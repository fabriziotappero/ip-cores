-------------------------------------------------------------------------------
--
-- The clock generation unit.
-- PHI1 clock and input/output clock enables are generated here.
--
-- $Id: t400_clkgen-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_clkgen_rtl_c0 of t400_clkgen is

  for rtl
  end for;

end t400_clkgen_rtl_c0;
