    wait;                               --
  end process;
end;
