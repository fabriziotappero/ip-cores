//This file was created by a tool wrietten with C.
module sim_rom (
    address,
    clock,
    q);
    input    [10:0]  address;
    input      clock;
    output    [11:0]  q;
    
reg [10:0]    address_latched;
// Instantiate the memory array itself.
reg [11:0]    mem[0:2048-1];
initial begin 
mem[0000] = 12'b101001100101;
mem[0001] = 12'b101000000011;
mem[0002] = 12'b101000011010;
mem[0003] = 12'b001000001110;
mem[0004] = 12'b000001101001;
mem[0005] = 12'b000010001101;
mem[0006] = 12'b011000000011;
mem[0007] = 12'b101000001011;
mem[0008] = 12'b001000001101;
mem[0009] = 12'b000000101000;
mem[0010] = 12'b101000010111;
mem[0011] = 12'b000001101000;
mem[0012] = 12'b110000001000;
mem[0013] = 12'b000000101111;
mem[0014] = 12'b001101101101;
mem[0015] = 12'b001101101000;
mem[0016] = 12'b001000001110;
mem[0017] = 12'b000010001000;
mem[0018] = 12'b011000000011;
mem[0019] = 12'b000000101000;
mem[0020] = 12'b001101101001;
mem[0021] = 12'b001011101111;
mem[0022] = 12'b101000001110;
mem[0023] = 12'b010010100011;
mem[0024] = 12'b010011000011;
mem[0025] = 12'b101001101110;
mem[0026] = 12'b001000001101;
mem[0027] = 12'b000000101000;
mem[0028] = 12'b001000101000;
mem[0029] = 12'b011001000011;
mem[0030] = 12'b101001000100;
mem[0031] = 12'b110000000001;
mem[0032] = 12'b000010001000;
mem[0033] = 12'b011001000011;
mem[0034] = 12'b101001000111;
mem[0035] = 12'b110000000010;
mem[0036] = 12'b000010001000;
mem[0037] = 12'b011001000011;
mem[0038] = 12'b101001001010;
mem[0039] = 12'b110000000011;
mem[0040] = 12'b000010001000;
mem[0041] = 12'b011001000011;
mem[0042] = 12'b101001001101;
mem[0043] = 12'b110000000100;
mem[0044] = 12'b000010001000;
mem[0045] = 12'b011001000011;
mem[0046] = 12'b101001010000;
mem[0047] = 12'b110000000101;
mem[0048] = 12'b000010001000;
mem[0049] = 12'b011001000011;
mem[0050] = 12'b101001010011;
mem[0051] = 12'b110000000110;
mem[0052] = 12'b000010001000;
mem[0053] = 12'b011001000011;
mem[0054] = 12'b101001010110;
mem[0055] = 12'b110000000111;
mem[0056] = 12'b000010001000;
mem[0057] = 12'b011001000011;
mem[0058] = 12'b101001011001;
mem[0059] = 12'b110000001000;
mem[0060] = 12'b000010001000;
mem[0061] = 12'b011001000011;
mem[0062] = 12'b101001011100;
mem[0063] = 12'b110000001001;
mem[0064] = 12'b000010001000;
mem[0065] = 12'b011001000011;
mem[0066] = 12'b101001011111;
mem[0067] = 12'b101001100010;
mem[0068] = 12'b110000110000;
mem[0069] = 12'b000000111111;
mem[0070] = 12'b101001100010;
mem[0071] = 12'b110000110001;
mem[0072] = 12'b000000111111;
mem[0073] = 12'b101001100010;
mem[0074] = 12'b110000110010;
mem[0075] = 12'b000000111111;
mem[0076] = 12'b101001100010;
mem[0077] = 12'b110000110011;
mem[0078] = 12'b000000111111;
mem[0079] = 12'b101001100010;
mem[0080] = 12'b110000110100;
mem[0081] = 12'b000000111111;
mem[0082] = 12'b101001100010;
mem[0083] = 12'b110000110101;
mem[0084] = 12'b000000111111;
mem[0085] = 12'b101001100010;
mem[0086] = 12'b110000110110;
mem[0087] = 12'b000000111111;
mem[0088] = 12'b101001100010;
mem[0089] = 12'b110000110111;
mem[0090] = 12'b000000111111;
mem[0091] = 12'b101001100010;
mem[0092] = 12'b110000111000;
mem[0093] = 12'b000000111111;
mem[0094] = 12'b101001100010;
mem[0095] = 12'b110000111001;
mem[0096] = 12'b000000111111;
mem[0097] = 12'b101001100010;
mem[0098] = 12'b010010100011;
mem[0099] = 12'b010011000011;
mem[0100] = 12'b101001110011;
mem[0101] = 12'b000001100100;
mem[0102] = 12'b000001101011;
mem[0103] = 12'b000001101100;
mem[0104] = 12'b001010101011;
mem[0105] = 12'b001000001011;
mem[0106] = 12'b000000101101;
mem[0107] = 12'b110000001010;
mem[0108] = 12'b000000101110;
mem[0109] = 12'b101000000001;
mem[0110] = 12'b001000001000;
mem[0111] = 12'b000000101011;
mem[0112] = 12'b001000001011;
mem[0113] = 12'b000000101101;
mem[0114] = 12'b101000000010;
mem[0115] = 12'b101001101000;
mem[0116] = 12'b000000000011;
mem[2047] = 12'b101000000000;
end
// Latch address
always @(posedge clock)
   address_latched <= address;
   
// READ
assign q = mem[address_latched];

endmodule

/*
0000: GOTO 101
0001: GOTO 3
0002: GOTO 26
0003: MOVFW 0x0e
0004: CLRF 0x09
0005: SUBWFW 0x0d
0006: BTFSC STATUS  [0]
0007: GOTO 11
0008: MOVFW 0x0d
0009: MOVWF 0x08
0010: GOTO 23
0011: CLRF 0x08
0012: MOVLW 8
0013: MOVWF 0x0f
0014: RLFF 0x0d
0015: RLFF 0x08
0016: MOVFW 0x0e
0017: SUBWFW 0x08
0018: BTFSC STATUS  [0]
0019: MOVWF 0x08
0020: RLFF 0x09
0021: DECFSZF 0x0f  [7]
0022: GOTO 14
0023: BCF STATUS  [5]
0024: BCF STATUS  [6]
0025: GOTO 110
0026: MOVFW 0x0d
0027: MOVWF 0x08
0028: MOVFF 0x08
0029: BTFSC STATUS  [2]
0030: GOTO 68
0031: MOVLW 1
0032: SUBWFW 0x08
0033: BTFSC STATUS  [2]
0034: GOTO 71
0035: MOVLW 2
0036: SUBWFW 0x08
0037: BTFSC STATUS  [2]
0038: GOTO 74
0039: MOVLW 3
0040: SUBWFW 0x08
0041: BTFSC STATUS  [2]
0042: GOTO 77
0043: MOVLW 4
0044: SUBWFW 0x08
0045: BTFSC STATUS  [2]
0046: GOTO 80
0047: MOVLW 5
0048: SUBWFW 0x08
0049: BTFSC STATUS  [2]
0050: GOTO 83
0051: MOVLW 6
0052: SUBWFW 0x08
0053: BTFSC STATUS  [2]
0054: GOTO 86
0055: MOVLW 7
0056: SUBWFW 0x08
0057: BTFSC STATUS  [2]
0058: GOTO 89
0059: MOVLW 8
0060: SUBWFW 0x08
0061: BTFSC STATUS  [2]
0062: GOTO 92
0063: MOVLW 9
0064: SUBWFW 0x08
0065: BTFSC STATUS  [2]
0066: GOTO 95
0067: GOTO 98
0068: MOVLW 48
0069: MOVWF 0x1f
0070: GOTO 98
0071: MOVLW 49
0072: MOVWF 0x1f
0073: GOTO 98
0074: MOVLW 50
0075: MOVWF 0x1f
0076: GOTO 98
0077: MOVLW 51
0078: MOVWF 0x1f
0079: GOTO 98
0080: MOVLW 52
0081: MOVWF 0x1f
0082: GOTO 98
0083: MOVLW 53
0084: MOVWF 0x1f
0085: GOTO 98
0086: MOVLW 54
0087: MOVWF 0x1f
0088: GOTO 98
0089: MOVLW 55
0090: MOVWF 0x1f
0091: GOTO 98
0092: MOVLW 56
0093: MOVWF 0x1f
0094: GOTO 98
0095: MOVLW 57
0096: MOVWF 0x1f
0097: GOTO 98
0098: BCF STATUS  [5]
0099: BCF STATUS  [6]
0100: GOTO 115
0101: CLRF FSR
0102: CLRF 0x0b
0103: CLRF 0x0c
0104: INCFF 0x0b
0105: MOVFW 0x0b
0106: MOVWF 0x0d
0107: MOVLW 10
0108: MOVWF 0x0e
0109: GOTO 1
0110: MOVFW 0x08
0111: MOVWF 0x0b
0112: MOVFW 0x0b
0113: MOVWF 0x0d
0114: GOTO 2
0115: GOTO 104
0116: NOP
2047: GOTO 0
*/
/*
covered instructions:

GOTO
MOVFW
CLRF
SUBWFW
BTFSC
MOVWF
MOVLW
RLFF
DECFSZF
BCF
MOVFF
INCFF
NOP
*/
