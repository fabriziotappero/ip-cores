entity csl_ctrl is
end entity;

architecture ctrl of  csl_ctrl is
begin
        -- 0in set_clock iClk -default
        -- 0in default_reset iRstSync -active_high -sync
end ctrl;

