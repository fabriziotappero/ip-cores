`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:01:47 02/03/2009 
// Design Name: Move map generator
// Module Name:    moves_map 
// Project Name: The FPGA Othello
// Target Devices: Spartan 3E, @50MHz
// Tool versions: 
// Description: 
//     1cc, combinational.
// Dependencies: 
//    n/a
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//         Marius TIVADAR.
//////////////////////////////////////////////////////////////////////////////////
module moves_map(clk, RST, B_, R_, player, M_);
input [63:0] B_;
input [63:0] R_;
input player;
input clk;
input RST;
output [63:0] M_;


wire [63:0] B;
wire [63:0] R;
reg [7:0] M [7:0][7:0];

reg [63:0] RES_Q;
reg [63:0] RES_D;

parameter ZEROP   = 3'd0;
parameter DOWN45P = 3'd1;
parameter DOWN    = 3'd2;
parameter DOWN45M = 3'd3;
parameter ZEROM   = 3'd4;
parameter UP45M   = 3'd5;
parameter UP      = 3'd6;
parameter UP45P   = 3'd7;

always @(posedge clk) begin
	if ( RST ) begin
		RES_Q <= 64'b0;
	end
	else begin
		RES_Q <= RES_D;
	end
end

/* continuous assignment, inputs are function of player */
assign R = (player) ? B_ : R_;
assign B = (player) ? R_ : B_;

always @( R or B ) begin


// Expresii generate pentru patrate A
    M[0][0][ZEROP] = (!R[0*8 + 0] && !B[0*8 + 0]) && 

                 (
                 (R[1*8 + 1] && B[2*8 + 2]) ||
                 (R[1*8 + 1] && R[2*8 + 2] && B[3*8 + 3]) ||
                 (R[1*8 + 1] && R[2*8 + 2] && R[3*8 + 3] && B[4*8 + 4]) ||
                 (R[1*8 + 1] && R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && B[5*8 + 5]) ||
                 (R[1*8 + 1] && R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && B[6*8 + 6]) ||
                 (R[1*8 + 1] && R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && R[6*8 + 6] && B[7*8 + 7]) 
                 );
    M[0][0][DOWN45P] = 1'b0;
    M[0][0][DOWN] = 1'b0;
    M[0][0][DOWN45M] = 1'b0;
    M[0][0][ZEROM] = (!R[0*8 + 0] && !B[0*8 + 0]) && 

                 (
                 (R[0*8 + 1] && B[0*8 + 2]) ||
                 (R[0*8 + 1] && R[0*8 + 2] && B[0*8 + 3]) ||
                 (R[0*8 + 1] && R[0*8 + 2] && R[0*8 + 3] && B[0*8 + 4]) ||
                 (R[0*8 + 1] && R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && B[0*8 + 5]) ||
                 (R[0*8 + 1] && R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && B[0*8 + 6]) ||
                 (R[0*8 + 1] && R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][0][UP45M] = (!R[0*8 + 0] && !B[0*8 + 0]) && 

                 (
                 (R[1*8 + 0] && B[2*8 + 0]) ||
                 (R[1*8 + 0] && R[2*8 + 0] && B[3*8 + 0]) ||
                 (R[1*8 + 0] && R[2*8 + 0] && R[3*8 + 0] && B[4*8 + 0]) ||
                 (R[1*8 + 0] && R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && B[5*8 + 0]) ||
                 (R[1*8 + 0] && R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && B[6*8 + 0]) ||
                 (R[1*8 + 0] && R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[0][0][UP] = 1'b0;
    M[0][0][UP45P] = 1'b0;
    M[0][7][ZEROP] = 1'b0;
    M[0][7][DOWN45P] = (!R[0*8 + 7] && !B[0*8 + 7]) && 

                 (
                 (R[1*8 + 6] && B[2*8 + 5]) ||
                 (R[1*8 + 6] && R[2*8 + 5] && B[3*8 + 4]) ||
                 (R[1*8 + 6] && R[2*8 + 5] && R[3*8 + 4] && B[4*8 + 3]) ||
                 (R[1*8 + 6] && R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && B[5*8 + 2]) ||
                 (R[1*8 + 6] && R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && B[6*8 + 1]) ||
                 (R[1*8 + 6] && R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && R[6*8 + 1] && B[7*8 + 0]) 
                 );
    M[0][7][DOWN] = 1'b0;
    M[0][7][DOWN45M] = 1'b0;
    M[0][7][ZEROM] = 1'b0;
    M[0][7][UP45M] = (!R[0*8 + 7] && !B[0*8 + 7]) && 

                 (
                 (R[1*8 + 7] && B[2*8 + 7]) ||
                 (R[1*8 + 7] && R[2*8 + 7] && B[3*8 + 7]) ||
                 (R[1*8 + 7] && R[2*8 + 7] && R[3*8 + 7] && B[4*8 + 7]) ||
                 (R[1*8 + 7] && R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && B[5*8 + 7]) ||
                 (R[1*8 + 7] && R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && B[6*8 + 7]) ||
                 (R[1*8 + 7] && R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[0][7][UP] = 1'b0;
    M[0][7][UP45P] = (!R[0*8 + 7] && !B[0*8 + 7]) && 

                 (
                 (R[0*8 + 6] && B[0*8 + 5]) ||
                 (R[0*8 + 6] && R[0*8 + 5] && B[0*8 + 4]) ||
                 (R[0*8 + 6] && R[0*8 + 5] && R[0*8 + 4] && B[0*8 + 3]) ||
                 (R[0*8 + 6] && R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && B[0*8 + 2]) ||
                 (R[0*8 + 6] && R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && B[0*8 + 1]) ||
                 (R[0*8 + 6] && R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[7][7][ZEROP] = 1'b0;
    M[7][7][DOWN45P] = 1'b0;
    M[7][7][DOWN] = (!R[7*8 + 7] && !B[7*8 + 7]) && 

                 (
                 (R[6*8 + 6] && B[5*8 + 5]) ||
                 (R[6*8 + 6] && R[5*8 + 5] && B[4*8 + 4]) ||
                 (R[6*8 + 6] && R[5*8 + 5] && R[4*8 + 4] && B[3*8 + 3]) ||
                 (R[6*8 + 6] && R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && B[2*8 + 2]) ||
                 (R[6*8 + 6] && R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && B[1*8 + 1]) ||
                 (R[6*8 + 6] && R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && R[1*8 + 1] && B[0*8 + 0]) 
                 );
    M[7][7][DOWN45M] = 1'b0;
    M[7][7][ZEROM] = 1'b0;
    M[7][7][UP45M] = 1'b0;
    M[7][7][UP] = (!R[7*8 + 7] && !B[7*8 + 7]) && 

                 (
                 (R[6*8 + 7] && B[5*8 + 7]) ||
                 (R[6*8 + 7] && R[5*8 + 7] && B[4*8 + 7]) ||
                 (R[6*8 + 7] && R[5*8 + 7] && R[4*8 + 7] && B[3*8 + 7]) ||
                 (R[6*8 + 7] && R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && B[2*8 + 7]) ||
                 (R[6*8 + 7] && R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && B[1*8 + 7]) ||
                 (R[6*8 + 7] && R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[7][7][UP45P] = (!R[7*8 + 7] && !B[7*8 + 7]) && 

                 (
                 (R[7*8 + 6] && B[7*8 + 5]) ||
                 (R[7*8 + 6] && R[7*8 + 5] && B[7*8 + 4]) ||
                 (R[7*8 + 6] && R[7*8 + 5] && R[7*8 + 4] && B[7*8 + 3]) ||
                 (R[7*8 + 6] && R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && B[7*8 + 2]) ||
                 (R[7*8 + 6] && R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && B[7*8 + 1]) ||
                 (R[7*8 + 6] && R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[7][0][ZEROP] = 1'b0;
    M[7][0][DOWN45P] = 1'b0;
    M[7][0][DOWN] = 1'b0;
    M[7][0][DOWN45M] = (!R[7*8 + 0] && !B[7*8 + 0]) && 

                 (
                 (R[6*8 + 1] && B[5*8 + 2]) ||
                 (R[6*8 + 1] && R[5*8 + 2] && B[4*8 + 3]) ||
                 (R[6*8 + 1] && R[5*8 + 2] && R[4*8 + 3] && B[3*8 + 4]) ||
                 (R[6*8 + 1] && R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && B[2*8 + 5]) ||
                 (R[6*8 + 1] && R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && B[1*8 + 6]) ||
                 (R[6*8 + 1] && R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && R[1*8 + 6] && B[0*8 + 7]) 
                 );
    M[7][0][ZEROM] = (!R[7*8 + 0] && !B[7*8 + 0]) && 

                 (
                 (R[7*8 + 1] && B[7*8 + 2]) ||
                 (R[7*8 + 1] && R[7*8 + 2] && B[7*8 + 3]) ||
                 (R[7*8 + 1] && R[7*8 + 2] && R[7*8 + 3] && B[7*8 + 4]) ||
                 (R[7*8 + 1] && R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && B[7*8 + 5]) ||
                 (R[7*8 + 1] && R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && B[7*8 + 6]) ||
                 (R[7*8 + 1] && R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][0][UP45M] = 1'b0;
    M[7][0][UP] = (!R[7*8 + 0] && !B[7*8 + 0]) && 

                 (
                 (R[6*8 + 0] && B[5*8 + 0]) ||
                 (R[6*8 + 0] && R[5*8 + 0] && B[4*8 + 0]) ||
                 (R[6*8 + 0] && R[5*8 + 0] && R[4*8 + 0] && B[3*8 + 0]) ||
                 (R[6*8 + 0] && R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && B[2*8 + 0]) ||
                 (R[6*8 + 0] && R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && B[1*8 + 0]) ||
                 (R[6*8 + 0] && R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[7][0][UP45P] = 1'b0;


// Expresii generate pentru patrate B
    M[0][1][ZEROP] = (!R[0*8 + 1] && !B[0*8 + 1]) && 

                 (
                 (R[1*8 + 2] && B[2*8 + 3]) ||
                 (R[1*8 + 2] && R[2*8 + 3] && B[3*8 + 4]) ||
                 (R[1*8 + 2] && R[2*8 + 3] && R[3*8 + 4] && B[4*8 + 5]) ||
                 (R[1*8 + 2] && R[2*8 + 3] && R[3*8 + 4] && R[4*8 + 5] && B[5*8 + 6]) ||
                 (R[1*8 + 2] && R[2*8 + 3] && R[3*8 + 4] && R[4*8 + 5] && R[5*8 + 6] && B[6*8 + 7]) 
                 );
    M[0][1][DOWN45P] = 1'b0;
    M[0][1][DOWN] = 1'b0;
    M[0][1][DOWN45M] = 1'b0;
    M[0][1][ZEROM] = (!R[0*8 + 1] && !B[0*8 + 1]) && 

                 (
                 (R[0*8 + 2] && B[0*8 + 3]) ||
                 (R[0*8 + 2] && R[0*8 + 3] && B[0*8 + 4]) ||
                 (R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && B[0*8 + 5]) ||
                 (R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && B[0*8 + 6]) ||
                 (R[0*8 + 2] && R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][1][UP45M] = (!R[0*8 + 1] && !B[0*8 + 1]) && 

                 (
                 (R[1*8 + 1] && B[2*8 + 1]) ||
                 (R[1*8 + 1] && R[2*8 + 1] && B[3*8 + 1]) ||
                 (R[1*8 + 1] && R[2*8 + 1] && R[3*8 + 1] && B[4*8 + 1]) ||
                 (R[1*8 + 1] && R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && B[5*8 + 1]) ||
                 (R[1*8 + 1] && R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && B[6*8 + 1]) ||
                 (R[1*8 + 1] && R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[0][1][UP] = 1'b0;
    M[0][1][UP45P] = 1'b0;
    M[0][6][ZEROP] = 1'b0;
    M[0][6][DOWN45P] = (!R[0*8 + 6] && !B[0*8 + 6]) && 

                 (
                 (R[1*8 + 5] && B[2*8 + 4]) ||
                 (R[1*8 + 5] && R[2*8 + 4] && B[3*8 + 3]) ||
                 (R[1*8 + 5] && R[2*8 + 4] && R[3*8 + 3] && B[4*8 + 2]) ||
                 (R[1*8 + 5] && R[2*8 + 4] && R[3*8 + 3] && R[4*8 + 2] && B[5*8 + 1]) ||
                 (R[1*8 + 5] && R[2*8 + 4] && R[3*8 + 3] && R[4*8 + 2] && R[5*8 + 1] && B[6*8 + 0]) 
                 );
    M[0][6][DOWN] = 1'b0;
    M[0][6][DOWN45M] = 1'b0;
    M[0][6][ZEROM] = 1'b0;
    M[0][6][UP45M] = (!R[0*8 + 6] && !B[0*8 + 6]) && 

                 (
                 (R[1*8 + 6] && B[2*8 + 6]) ||
                 (R[1*8 + 6] && R[2*8 + 6] && B[3*8 + 6]) ||
                 (R[1*8 + 6] && R[2*8 + 6] && R[3*8 + 6] && B[4*8 + 6]) ||
                 (R[1*8 + 6] && R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && B[5*8 + 6]) ||
                 (R[1*8 + 6] && R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && B[6*8 + 6]) ||
                 (R[1*8 + 6] && R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[0][6][UP] = 1'b0;
    M[0][6][UP45P] = (!R[0*8 + 6] && !B[0*8 + 6]) && 

                 (
                 (R[0*8 + 5] && B[0*8 + 4]) ||
                 (R[0*8 + 5] && R[0*8 + 4] && B[0*8 + 3]) ||
                 (R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && B[0*8 + 2]) ||
                 (R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && B[0*8 + 1]) ||
                 (R[0*8 + 5] && R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[1][7][ZEROP] = 1'b0;
    M[1][7][DOWN45P] = (!R[1*8 + 7] && !B[1*8 + 7]) && 

                 (
                 (R[2*8 + 6] && B[3*8 + 5]) ||
                 (R[2*8 + 6] && R[3*8 + 5] && B[4*8 + 4]) ||
                 (R[2*8 + 6] && R[3*8 + 5] && R[4*8 + 4] && B[5*8 + 3]) ||
                 (R[2*8 + 6] && R[3*8 + 5] && R[4*8 + 4] && R[5*8 + 3] && B[6*8 + 2]) ||
                 (R[2*8 + 6] && R[3*8 + 5] && R[4*8 + 4] && R[5*8 + 3] && R[6*8 + 2] && B[7*8 + 1]) 
                 );
    M[1][7][DOWN] = 1'b0;
    M[1][7][DOWN45M] = 1'b0;
    M[1][7][ZEROM] = 1'b0;
    M[1][7][UP45M] = (!R[1*8 + 7] && !B[1*8 + 7]) && 

                 (
                 (R[2*8 + 7] && B[3*8 + 7]) ||
                 (R[2*8 + 7] && R[3*8 + 7] && B[4*8 + 7]) ||
                 (R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && B[5*8 + 7]) ||
                 (R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && B[6*8 + 7]) ||
                 (R[2*8 + 7] && R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[1][7][UP] = 1'b0;
    M[1][7][UP45P] = (!R[1*8 + 7] && !B[1*8 + 7]) && 

                 (
                 (R[1*8 + 6] && B[1*8 + 5]) ||
                 (R[1*8 + 6] && R[1*8 + 5] && B[1*8 + 4]) ||
                 (R[1*8 + 6] && R[1*8 + 5] && R[1*8 + 4] && B[1*8 + 3]) ||
                 (R[1*8 + 6] && R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && B[1*8 + 2]) ||
                 (R[1*8 + 6] && R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && B[1*8 + 1]) ||
                 (R[1*8 + 6] && R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[6][7][ZEROP] = 1'b0;
    M[6][7][DOWN45P] = 1'b0;
    M[6][7][DOWN] = (!R[6*8 + 7] && !B[6*8 + 7]) && 

                 (
                 (R[5*8 + 6] && B[4*8 + 5]) ||
                 (R[5*8 + 6] && R[4*8 + 5] && B[3*8 + 4]) ||
                 (R[5*8 + 6] && R[4*8 + 5] && R[3*8 + 4] && B[2*8 + 3]) ||
                 (R[5*8 + 6] && R[4*8 + 5] && R[3*8 + 4] && R[2*8 + 3] && B[1*8 + 2]) ||
                 (R[5*8 + 6] && R[4*8 + 5] && R[3*8 + 4] && R[2*8 + 3] && R[1*8 + 2] && B[0*8 + 1]) 
                 );
    M[6][7][DOWN45M] = 1'b0;
    M[6][7][ZEROM] = 1'b0;
    M[6][7][UP45M] = 1'b0;
    M[6][7][UP] = (!R[6*8 + 7] && !B[6*8 + 7]) && 

                 (
                 (R[5*8 + 7] && B[4*8 + 7]) ||
                 (R[5*8 + 7] && R[4*8 + 7] && B[3*8 + 7]) ||
                 (R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && B[2*8 + 7]) ||
                 (R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && B[1*8 + 7]) ||
                 (R[5*8 + 7] && R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[6][7][UP45P] = (!R[6*8 + 7] && !B[6*8 + 7]) && 

                 (
                 (R[6*8 + 6] && B[6*8 + 5]) ||
                 (R[6*8 + 6] && R[6*8 + 5] && B[6*8 + 4]) ||
                 (R[6*8 + 6] && R[6*8 + 5] && R[6*8 + 4] && B[6*8 + 3]) ||
                 (R[6*8 + 6] && R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && B[6*8 + 2]) ||
                 (R[6*8 + 6] && R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && B[6*8 + 1]) ||
                 (R[6*8 + 6] && R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[7][6][ZEROP] = 1'b0;
    M[7][6][DOWN45P] = 1'b0;
    M[7][6][DOWN] = (!R[7*8 + 6] && !B[7*8 + 6]) && 

                 (
                 (R[6*8 + 5] && B[5*8 + 4]) ||
                 (R[6*8 + 5] && R[5*8 + 4] && B[4*8 + 3]) ||
                 (R[6*8 + 5] && R[5*8 + 4] && R[4*8 + 3] && B[3*8 + 2]) ||
                 (R[6*8 + 5] && R[5*8 + 4] && R[4*8 + 3] && R[3*8 + 2] && B[2*8 + 1]) ||
                 (R[6*8 + 5] && R[5*8 + 4] && R[4*8 + 3] && R[3*8 + 2] && R[2*8 + 1] && B[1*8 + 0]) 
                 );
    M[7][6][DOWN45M] = 1'b0;
    M[7][6][ZEROM] = 1'b0;
    M[7][6][UP45M] = 1'b0;
    M[7][6][UP] = (!R[7*8 + 6] && !B[7*8 + 6]) && 

                 (
                 (R[6*8 + 6] && B[5*8 + 6]) ||
                 (R[6*8 + 6] && R[5*8 + 6] && B[4*8 + 6]) ||
                 (R[6*8 + 6] && R[5*8 + 6] && R[4*8 + 6] && B[3*8 + 6]) ||
                 (R[6*8 + 6] && R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && B[2*8 + 6]) ||
                 (R[6*8 + 6] && R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && B[1*8 + 6]) ||
                 (R[6*8 + 6] && R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[7][6][UP45P] = (!R[7*8 + 6] && !B[7*8 + 6]) && 

                 (
                 (R[7*8 + 5] && B[7*8 + 4]) ||
                 (R[7*8 + 5] && R[7*8 + 4] && B[7*8 + 3]) ||
                 (R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && B[7*8 + 2]) ||
                 (R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && B[7*8 + 1]) ||
                 (R[7*8 + 5] && R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[7][1][ZEROP] = 1'b0;
    M[7][1][DOWN45P] = 1'b0;
    M[7][1][DOWN] = 1'b0;
    M[7][1][DOWN45M] = (!R[7*8 + 1] && !B[7*8 + 1]) && 

                 (
                 (R[6*8 + 2] && B[5*8 + 3]) ||
                 (R[6*8 + 2] && R[5*8 + 3] && B[4*8 + 4]) ||
                 (R[6*8 + 2] && R[5*8 + 3] && R[4*8 + 4] && B[3*8 + 5]) ||
                 (R[6*8 + 2] && R[5*8 + 3] && R[4*8 + 4] && R[3*8 + 5] && B[2*8 + 6]) ||
                 (R[6*8 + 2] && R[5*8 + 3] && R[4*8 + 4] && R[3*8 + 5] && R[2*8 + 6] && B[1*8 + 7]) 
                 );
    M[7][1][ZEROM] = (!R[7*8 + 1] && !B[7*8 + 1]) && 

                 (
                 (R[7*8 + 2] && B[7*8 + 3]) ||
                 (R[7*8 + 2] && R[7*8 + 3] && B[7*8 + 4]) ||
                 (R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && B[7*8 + 5]) ||
                 (R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && B[7*8 + 6]) ||
                 (R[7*8 + 2] && R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][1][UP45M] = 1'b0;
    M[7][1][UP] = (!R[7*8 + 1] && !B[7*8 + 1]) && 

                 (
                 (R[6*8 + 1] && B[5*8 + 1]) ||
                 (R[6*8 + 1] && R[5*8 + 1] && B[4*8 + 1]) ||
                 (R[6*8 + 1] && R[5*8 + 1] && R[4*8 + 1] && B[3*8 + 1]) ||
                 (R[6*8 + 1] && R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && B[2*8 + 1]) ||
                 (R[6*8 + 1] && R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && B[1*8 + 1]) ||
                 (R[6*8 + 1] && R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[7][1][UP45P] = 1'b0;
    M[6][0][ZEROP] = 1'b0;
    M[6][0][DOWN45P] = 1'b0;
    M[6][0][DOWN] = 1'b0;
    M[6][0][DOWN45M] = (!R[6*8 + 0] && !B[6*8 + 0]) && 

                 (
                 (R[5*8 + 1] && B[4*8 + 2]) ||
                 (R[5*8 + 1] && R[4*8 + 2] && B[3*8 + 3]) ||
                 (R[5*8 + 1] && R[4*8 + 2] && R[3*8 + 3] && B[2*8 + 4]) ||
                 (R[5*8 + 1] && R[4*8 + 2] && R[3*8 + 3] && R[2*8 + 4] && B[1*8 + 5]) ||
                 (R[5*8 + 1] && R[4*8 + 2] && R[3*8 + 3] && R[2*8 + 4] && R[1*8 + 5] && B[0*8 + 6]) 
                 );
    M[6][0][ZEROM] = (!R[6*8 + 0] && !B[6*8 + 0]) && 

                 (
                 (R[6*8 + 1] && B[6*8 + 2]) ||
                 (R[6*8 + 1] && R[6*8 + 2] && B[6*8 + 3]) ||
                 (R[6*8 + 1] && R[6*8 + 2] && R[6*8 + 3] && B[6*8 + 4]) ||
                 (R[6*8 + 1] && R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && B[6*8 + 5]) ||
                 (R[6*8 + 1] && R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && B[6*8 + 6]) ||
                 (R[6*8 + 1] && R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][0][UP45M] = 1'b0;
    M[6][0][UP] = (!R[6*8 + 0] && !B[6*8 + 0]) && 

                 (
                 (R[5*8 + 0] && B[4*8 + 0]) ||
                 (R[5*8 + 0] && R[4*8 + 0] && B[3*8 + 0]) ||
                 (R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && B[2*8 + 0]) ||
                 (R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && B[1*8 + 0]) ||
                 (R[5*8 + 0] && R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[6][0][UP45P] = 1'b0;
    M[1][0][ZEROP] = (!R[1*8 + 0] && !B[1*8 + 0]) && 

                 (
                 (R[2*8 + 1] && B[3*8 + 2]) ||
                 (R[2*8 + 1] && R[3*8 + 2] && B[4*8 + 3]) ||
                 (R[2*8 + 1] && R[3*8 + 2] && R[4*8 + 3] && B[5*8 + 4]) ||
                 (R[2*8 + 1] && R[3*8 + 2] && R[4*8 + 3] && R[5*8 + 4] && B[6*8 + 5]) ||
                 (R[2*8 + 1] && R[3*8 + 2] && R[4*8 + 3] && R[5*8 + 4] && R[6*8 + 5] && B[7*8 + 6]) 
                 );
    M[1][0][DOWN45P] = 1'b0;
    M[1][0][DOWN] = 1'b0;
    M[1][0][DOWN45M] = 1'b0;
    M[1][0][ZEROM] = (!R[1*8 + 0] && !B[1*8 + 0]) && 

                 (
                 (R[1*8 + 1] && B[1*8 + 2]) ||
                 (R[1*8 + 1] && R[1*8 + 2] && B[1*8 + 3]) ||
                 (R[1*8 + 1] && R[1*8 + 2] && R[1*8 + 3] && B[1*8 + 4]) ||
                 (R[1*8 + 1] && R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && B[1*8 + 5]) ||
                 (R[1*8 + 1] && R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && B[1*8 + 6]) ||
                 (R[1*8 + 1] && R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][0][UP45M] = (!R[1*8 + 0] && !B[1*8 + 0]) && 

                 (
                 (R[2*8 + 0] && B[3*8 + 0]) ||
                 (R[2*8 + 0] && R[3*8 + 0] && B[4*8 + 0]) ||
                 (R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && B[5*8 + 0]) ||
                 (R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && B[6*8 + 0]) ||
                 (R[2*8 + 0] && R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[1][0][UP] = 1'b0;
    M[1][0][UP45P] = 1'b0;


// Expresii generate pentru patrate C
    M[0][2][ZEROP] = (!R[0*8 + 2] && !B[0*8 + 2]) && 

                 (
                 (R[1*8 + 3] && B[2*8 + 4]) ||
                 (R[1*8 + 3] && R[2*8 + 4] && B[3*8 + 5]) ||
                 (R[1*8 + 3] && R[2*8 + 4] && R[3*8 + 5] && B[4*8 + 6]) ||
                 (R[1*8 + 3] && R[2*8 + 4] && R[3*8 + 5] && R[4*8 + 6] && B[5*8 + 7]) 
                 );
    M[0][2][DOWN45P] = (!R[0*8 + 2] && !B[0*8 + 2]) && 

                 (
                 (R[1*8 + 1] && B[2*8 + 0]) 
                 );
    M[0][2][DOWN] = 1'b0;
    M[0][2][DOWN45M] = 1'b0;
    M[0][2][ZEROM] = (!R[0*8 + 2] && !B[0*8 + 2]) && 

                 (
                 (R[0*8 + 3] && B[0*8 + 4]) ||
                 (R[0*8 + 3] && R[0*8 + 4] && B[0*8 + 5]) ||
                 (R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && B[0*8 + 6]) ||
                 (R[0*8 + 3] && R[0*8 + 4] && R[0*8 + 5] && R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][2][UP45M] = (!R[0*8 + 2] && !B[0*8 + 2]) && 

                 (
                 (R[1*8 + 2] && B[2*8 + 2]) ||
                 (R[1*8 + 2] && R[2*8 + 2] && B[3*8 + 2]) ||
                 (R[1*8 + 2] && R[2*8 + 2] && R[3*8 + 2] && B[4*8 + 2]) ||
                 (R[1*8 + 2] && R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && B[5*8 + 2]) ||
                 (R[1*8 + 2] && R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && B[6*8 + 2]) ||
                 (R[1*8 + 2] && R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[0][2][UP] = 1'b0;
    M[0][2][UP45P] = (!R[0*8 + 2] && !B[0*8 + 2]) && 

                 (
                 (R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[0][5][ZEROP] = (!R[0*8 + 5] && !B[0*8 + 5]) && 

                 (
                 (R[1*8 + 6] && B[2*8 + 7]) 
                 );
    M[0][5][DOWN45P] = (!R[0*8 + 5] && !B[0*8 + 5]) && 

                 (
                 (R[1*8 + 4] && B[2*8 + 3]) ||
                 (R[1*8 + 4] && R[2*8 + 3] && B[3*8 + 2]) ||
                 (R[1*8 + 4] && R[2*8 + 3] && R[3*8 + 2] && B[4*8 + 1]) ||
                 (R[1*8 + 4] && R[2*8 + 3] && R[3*8 + 2] && R[4*8 + 1] && B[5*8 + 0]) 
                 );
    M[0][5][DOWN] = 1'b0;
    M[0][5][DOWN45M] = 1'b0;
    M[0][5][ZEROM] = (!R[0*8 + 5] && !B[0*8 + 5]) && 

                 (
                 (R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][5][UP45M] = (!R[0*8 + 5] && !B[0*8 + 5]) && 

                 (
                 (R[1*8 + 5] && B[2*8 + 5]) ||
                 (R[1*8 + 5] && R[2*8 + 5] && B[3*8 + 5]) ||
                 (R[1*8 + 5] && R[2*8 + 5] && R[3*8 + 5] && B[4*8 + 5]) ||
                 (R[1*8 + 5] && R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && B[5*8 + 5]) ||
                 (R[1*8 + 5] && R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && B[6*8 + 5]) ||
                 (R[1*8 + 5] && R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[0][5][UP] = 1'b0;
    M[0][5][UP45P] = (!R[0*8 + 5] && !B[0*8 + 5]) && 

                 (
                 (R[0*8 + 4] && B[0*8 + 3]) ||
                 (R[0*8 + 4] && R[0*8 + 3] && B[0*8 + 2]) ||
                 (R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && B[0*8 + 1]) ||
                 (R[0*8 + 4] && R[0*8 + 3] && R[0*8 + 2] && R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[2][7][ZEROP] = 1'b0;
    M[2][7][DOWN45P] = (!R[2*8 + 7] && !B[2*8 + 7]) && 

                 (
                 (R[3*8 + 6] && B[4*8 + 5]) ||
                 (R[3*8 + 6] && R[4*8 + 5] && B[5*8 + 4]) ||
                 (R[3*8 + 6] && R[4*8 + 5] && R[5*8 + 4] && B[6*8 + 3]) ||
                 (R[3*8 + 6] && R[4*8 + 5] && R[5*8 + 4] && R[6*8 + 3] && B[7*8 + 2]) 
                 );
    M[2][7][DOWN] = (!R[2*8 + 7] && !B[2*8 + 7]) && 

                 (
                 (R[1*8 + 6] && B[0*8 + 5]) 
                 );
    M[2][7][DOWN45M] = 1'b0;
    M[2][7][ZEROM] = 1'b0;
    M[2][7][UP45M] = (!R[2*8 + 7] && !B[2*8 + 7]) && 

                 (
                 (R[3*8 + 7] && B[4*8 + 7]) ||
                 (R[3*8 + 7] && R[4*8 + 7] && B[5*8 + 7]) ||
                 (R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && B[6*8 + 7]) ||
                 (R[3*8 + 7] && R[4*8 + 7] && R[5*8 + 7] && R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[2][7][UP] = (!R[2*8 + 7] && !B[2*8 + 7]) && 

                 (
                 (R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[2][7][UP45P] = (!R[2*8 + 7] && !B[2*8 + 7]) && 

                 (
                 (R[2*8 + 6] && B[2*8 + 5]) ||
                 (R[2*8 + 6] && R[2*8 + 5] && B[2*8 + 4]) ||
                 (R[2*8 + 6] && R[2*8 + 5] && R[2*8 + 4] && B[2*8 + 3]) ||
                 (R[2*8 + 6] && R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && B[2*8 + 2]) ||
                 (R[2*8 + 6] && R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && B[2*8 + 1]) ||
                 (R[2*8 + 6] && R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[5][7][ZEROP] = 1'b0;
    M[5][7][DOWN45P] = (!R[5*8 + 7] && !B[5*8 + 7]) && 

                 (
                 (R[6*8 + 6] && B[7*8 + 5]) 
                 );
    M[5][7][DOWN] = (!R[5*8 + 7] && !B[5*8 + 7]) && 

                 (
                 (R[4*8 + 6] && B[3*8 + 5]) ||
                 (R[4*8 + 6] && R[3*8 + 5] && B[2*8 + 4]) ||
                 (R[4*8 + 6] && R[3*8 + 5] && R[2*8 + 4] && B[1*8 + 3]) ||
                 (R[4*8 + 6] && R[3*8 + 5] && R[2*8 + 4] && R[1*8 + 3] && B[0*8 + 2]) 
                 );
    M[5][7][DOWN45M] = 1'b0;
    M[5][7][ZEROM] = 1'b0;
    M[5][7][UP45M] = (!R[5*8 + 7] && !B[5*8 + 7]) && 

                 (
                 (R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[5][7][UP] = (!R[5*8 + 7] && !B[5*8 + 7]) && 

                 (
                 (R[4*8 + 7] && B[3*8 + 7]) ||
                 (R[4*8 + 7] && R[3*8 + 7] && B[2*8 + 7]) ||
                 (R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && B[1*8 + 7]) ||
                 (R[4*8 + 7] && R[3*8 + 7] && R[2*8 + 7] && R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[5][7][UP45P] = (!R[5*8 + 7] && !B[5*8 + 7]) && 

                 (
                 (R[5*8 + 6] && B[5*8 + 5]) ||
                 (R[5*8 + 6] && R[5*8 + 5] && B[5*8 + 4]) ||
                 (R[5*8 + 6] && R[5*8 + 5] && R[5*8 + 4] && B[5*8 + 3]) ||
                 (R[5*8 + 6] && R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && B[5*8 + 2]) ||
                 (R[5*8 + 6] && R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && B[5*8 + 1]) ||
                 (R[5*8 + 6] && R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && R[5*8 + 1] && B[5*8 + 0]) 
                 );
    M[7][5][ZEROP] = 1'b0;
    M[7][5][DOWN45P] = 1'b0;
    M[7][5][DOWN] = (!R[7*8 + 5] && !B[7*8 + 5]) && 

                 (
                 (R[6*8 + 4] && B[5*8 + 3]) ||
                 (R[6*8 + 4] && R[5*8 + 3] && B[4*8 + 2]) ||
                 (R[6*8 + 4] && R[5*8 + 3] && R[4*8 + 2] && B[3*8 + 1]) ||
                 (R[6*8 + 4] && R[5*8 + 3] && R[4*8 + 2] && R[3*8 + 1] && B[2*8 + 0]) 
                 );
    M[7][5][DOWN45M] = (!R[7*8 + 5] && !B[7*8 + 5]) && 

                 (
                 (R[6*8 + 6] && B[5*8 + 7]) 
                 );
    M[7][5][ZEROM] = (!R[7*8 + 5] && !B[7*8 + 5]) && 

                 (
                 (R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][5][UP45M] = 1'b0;
    M[7][5][UP] = (!R[7*8 + 5] && !B[7*8 + 5]) && 

                 (
                 (R[6*8 + 5] && B[5*8 + 5]) ||
                 (R[6*8 + 5] && R[5*8 + 5] && B[4*8 + 5]) ||
                 (R[6*8 + 5] && R[5*8 + 5] && R[4*8 + 5] && B[3*8 + 5]) ||
                 (R[6*8 + 5] && R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && B[2*8 + 5]) ||
                 (R[6*8 + 5] && R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && B[1*8 + 5]) ||
                 (R[6*8 + 5] && R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[7][5][UP45P] = (!R[7*8 + 5] && !B[7*8 + 5]) && 

                 (
                 (R[7*8 + 4] && B[7*8 + 3]) ||
                 (R[7*8 + 4] && R[7*8 + 3] && B[7*8 + 2]) ||
                 (R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && B[7*8 + 1]) ||
                 (R[7*8 + 4] && R[7*8 + 3] && R[7*8 + 2] && R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[7][2][ZEROP] = 1'b0;
    M[7][2][DOWN45P] = 1'b0;
    M[7][2][DOWN] = (!R[7*8 + 2] && !B[7*8 + 2]) && 

                 (
                 (R[6*8 + 1] && B[5*8 + 0]) 
                 );
    M[7][2][DOWN45M] = (!R[7*8 + 2] && !B[7*8 + 2]) && 

                 (
                 (R[6*8 + 3] && B[5*8 + 4]) ||
                 (R[6*8 + 3] && R[5*8 + 4] && B[4*8 + 5]) ||
                 (R[6*8 + 3] && R[5*8 + 4] && R[4*8 + 5] && B[3*8 + 6]) ||
                 (R[6*8 + 3] && R[5*8 + 4] && R[4*8 + 5] && R[3*8 + 6] && B[2*8 + 7]) 
                 );
    M[7][2][ZEROM] = (!R[7*8 + 2] && !B[7*8 + 2]) && 

                 (
                 (R[7*8 + 3] && B[7*8 + 4]) ||
                 (R[7*8 + 3] && R[7*8 + 4] && B[7*8 + 5]) ||
                 (R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && B[7*8 + 6]) ||
                 (R[7*8 + 3] && R[7*8 + 4] && R[7*8 + 5] && R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][2][UP45M] = 1'b0;
    M[7][2][UP] = (!R[7*8 + 2] && !B[7*8 + 2]) && 

                 (
                 (R[6*8 + 2] && B[5*8 + 2]) ||
                 (R[6*8 + 2] && R[5*8 + 2] && B[4*8 + 2]) ||
                 (R[6*8 + 2] && R[5*8 + 2] && R[4*8 + 2] && B[3*8 + 2]) ||
                 (R[6*8 + 2] && R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && B[2*8 + 2]) ||
                 (R[6*8 + 2] && R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && B[1*8 + 2]) ||
                 (R[6*8 + 2] && R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[7][2][UP45P] = (!R[7*8 + 2] && !B[7*8 + 2]) && 

                 (
                 (R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[5][0][ZEROP] = (!R[5*8 + 0] && !B[5*8 + 0]) && 

                 (
                 (R[6*8 + 1] && B[7*8 + 2]) 
                 );
    M[5][0][DOWN45P] = 1'b0;
    M[5][0][DOWN] = 1'b0;
    M[5][0][DOWN45M] = (!R[5*8 + 0] && !B[5*8 + 0]) && 

                 (
                 (R[4*8 + 1] && B[3*8 + 2]) ||
                 (R[4*8 + 1] && R[3*8 + 2] && B[2*8 + 3]) ||
                 (R[4*8 + 1] && R[3*8 + 2] && R[2*8 + 3] && B[1*8 + 4]) ||
                 (R[4*8 + 1] && R[3*8 + 2] && R[2*8 + 3] && R[1*8 + 4] && B[0*8 + 5]) 
                 );
    M[5][0][ZEROM] = (!R[5*8 + 0] && !B[5*8 + 0]) && 

                 (
                 (R[5*8 + 1] && B[5*8 + 2]) ||
                 (R[5*8 + 1] && R[5*8 + 2] && B[5*8 + 3]) ||
                 (R[5*8 + 1] && R[5*8 + 2] && R[5*8 + 3] && B[5*8 + 4]) ||
                 (R[5*8 + 1] && R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && B[5*8 + 5]) ||
                 (R[5*8 + 1] && R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && B[5*8 + 6]) ||
                 (R[5*8 + 1] && R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][0][UP45M] = (!R[5*8 + 0] && !B[5*8 + 0]) && 

                 (
                 (R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[5][0][UP] = (!R[5*8 + 0] && !B[5*8 + 0]) && 

                 (
                 (R[4*8 + 0] && B[3*8 + 0]) ||
                 (R[4*8 + 0] && R[3*8 + 0] && B[2*8 + 0]) ||
                 (R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && B[1*8 + 0]) ||
                 (R[4*8 + 0] && R[3*8 + 0] && R[2*8 + 0] && R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[5][0][UP45P] = 1'b0;
    M[2][0][ZEROP] = (!R[2*8 + 0] && !B[2*8 + 0]) && 

                 (
                 (R[3*8 + 1] && B[4*8 + 2]) ||
                 (R[3*8 + 1] && R[4*8 + 2] && B[5*8 + 3]) ||
                 (R[3*8 + 1] && R[4*8 + 2] && R[5*8 + 3] && B[6*8 + 4]) ||
                 (R[3*8 + 1] && R[4*8 + 2] && R[5*8 + 3] && R[6*8 + 4] && B[7*8 + 5]) 
                 );
    M[2][0][DOWN45P] = 1'b0;
    M[2][0][DOWN] = 1'b0;
    M[2][0][DOWN45M] = (!R[2*8 + 0] && !B[2*8 + 0]) && 

                 (
                 (R[1*8 + 1] && B[0*8 + 2]) 
                 );
    M[2][0][ZEROM] = (!R[2*8 + 0] && !B[2*8 + 0]) && 

                 (
                 (R[2*8 + 1] && B[2*8 + 2]) ||
                 (R[2*8 + 1] && R[2*8 + 2] && B[2*8 + 3]) ||
                 (R[2*8 + 1] && R[2*8 + 2] && R[2*8 + 3] && B[2*8 + 4]) ||
                 (R[2*8 + 1] && R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && B[2*8 + 5]) ||
                 (R[2*8 + 1] && R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && B[2*8 + 6]) ||
                 (R[2*8 + 1] && R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][0][UP45M] = (!R[2*8 + 0] && !B[2*8 + 0]) && 

                 (
                 (R[3*8 + 0] && B[4*8 + 0]) ||
                 (R[3*8 + 0] && R[4*8 + 0] && B[5*8 + 0]) ||
                 (R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && B[6*8 + 0]) ||
                 (R[3*8 + 0] && R[4*8 + 0] && R[5*8 + 0] && R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[2][0][UP] = (!R[2*8 + 0] && !B[2*8 + 0]) && 

                 (
                 (R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[2][0][UP45P] = 1'b0;


// Expresii generate pentru patrate D
    M[0][3][ZEROP] = (!R[0*8 + 3] && !B[0*8 + 3]) && 

                 (
                 (R[1*8 + 4] && B[2*8 + 5]) ||
                 (R[1*8 + 4] && R[2*8 + 5] && B[3*8 + 6]) ||
                 (R[1*8 + 4] && R[2*8 + 5] && R[3*8 + 6] && B[4*8 + 7]) 
                 );
    M[0][3][DOWN45P] = (!R[0*8 + 3] && !B[0*8 + 3]) && 

                 (
                 (R[1*8 + 2] && B[2*8 + 1]) ||
                 (R[1*8 + 2] && R[2*8 + 1] && B[3*8 + 0]) 
                 );
    M[0][3][DOWN] = 1'b0;
    M[0][3][DOWN45M] = 1'b0;
    M[0][3][ZEROM] = (!R[0*8 + 3] && !B[0*8 + 3]) && 

                 (
                 (R[0*8 + 4] && B[0*8 + 5]) ||
                 (R[0*8 + 4] && R[0*8 + 5] && B[0*8 + 6]) ||
                 (R[0*8 + 4] && R[0*8 + 5] && R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][3][UP45M] = (!R[0*8 + 3] && !B[0*8 + 3]) && 

                 (
                 (R[1*8 + 3] && B[2*8 + 3]) ||
                 (R[1*8 + 3] && R[2*8 + 3] && B[3*8 + 3]) ||
                 (R[1*8 + 3] && R[2*8 + 3] && R[3*8 + 3] && B[4*8 + 3]) ||
                 (R[1*8 + 3] && R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && B[5*8 + 3]) ||
                 (R[1*8 + 3] && R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && B[6*8 + 3]) ||
                 (R[1*8 + 3] && R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && R[6*8 + 3] && B[7*8 + 3]) 
                 );
    M[0][3][UP] = 1'b0;
    M[0][3][UP45P] = (!R[0*8 + 3] && !B[0*8 + 3]) && 

                 (
                 (R[0*8 + 2] && B[0*8 + 1]) ||
                 (R[0*8 + 2] && R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[0][4][ZEROP] = (!R[0*8 + 4] && !B[0*8 + 4]) && 

                 (
                 (R[1*8 + 5] && B[2*8 + 6]) ||
                 (R[1*8 + 5] && R[2*8 + 6] && B[3*8 + 7]) 
                 );
    M[0][4][DOWN45P] = (!R[0*8 + 4] && !B[0*8 + 4]) && 

                 (
                 (R[1*8 + 3] && B[2*8 + 2]) ||
                 (R[1*8 + 3] && R[2*8 + 2] && B[3*8 + 1]) ||
                 (R[1*8 + 3] && R[2*8 + 2] && R[3*8 + 1] && B[4*8 + 0]) 
                 );
    M[0][4][DOWN] = 1'b0;
    M[0][4][DOWN45M] = 1'b0;
    M[0][4][ZEROM] = (!R[0*8 + 4] && !B[0*8 + 4]) && 

                 (
                 (R[0*8 + 5] && B[0*8 + 6]) ||
                 (R[0*8 + 5] && R[0*8 + 6] && B[0*8 + 7]) 
                 );
    M[0][4][UP45M] = (!R[0*8 + 4] && !B[0*8 + 4]) && 

                 (
                 (R[1*8 + 4] && B[2*8 + 4]) ||
                 (R[1*8 + 4] && R[2*8 + 4] && B[3*8 + 4]) ||
                 (R[1*8 + 4] && R[2*8 + 4] && R[3*8 + 4] && B[4*8 + 4]) ||
                 (R[1*8 + 4] && R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && B[5*8 + 4]) ||
                 (R[1*8 + 4] && R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && B[6*8 + 4]) ||
                 (R[1*8 + 4] && R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && R[6*8 + 4] && B[7*8 + 4]) 
                 );
    M[0][4][UP] = 1'b0;
    M[0][4][UP45P] = (!R[0*8 + 4] && !B[0*8 + 4]) && 

                 (
                 (R[0*8 + 3] && B[0*8 + 2]) ||
                 (R[0*8 + 3] && R[0*8 + 2] && B[0*8 + 1]) ||
                 (R[0*8 + 3] && R[0*8 + 2] && R[0*8 + 1] && B[0*8 + 0]) 
                 );
    M[3][7][ZEROP] = 1'b0;
    M[3][7][DOWN45P] = (!R[3*8 + 7] && !B[3*8 + 7]) && 

                 (
                 (R[4*8 + 6] && B[5*8 + 5]) ||
                 (R[4*8 + 6] && R[5*8 + 5] && B[6*8 + 4]) ||
                 (R[4*8 + 6] && R[5*8 + 5] && R[6*8 + 4] && B[7*8 + 3]) 
                 );
    M[3][7][DOWN] = (!R[3*8 + 7] && !B[3*8 + 7]) && 

                 (
                 (R[2*8 + 6] && B[1*8 + 5]) ||
                 (R[2*8 + 6] && R[1*8 + 5] && B[0*8 + 4]) 
                 );
    M[3][7][DOWN45M] = 1'b0;
    M[3][7][ZEROM] = 1'b0;
    M[3][7][UP45M] = (!R[3*8 + 7] && !B[3*8 + 7]) && 

                 (
                 (R[4*8 + 7] && B[5*8 + 7]) ||
                 (R[4*8 + 7] && R[5*8 + 7] && B[6*8 + 7]) ||
                 (R[4*8 + 7] && R[5*8 + 7] && R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[3][7][UP] = (!R[3*8 + 7] && !B[3*8 + 7]) && 

                 (
                 (R[2*8 + 7] && B[1*8 + 7]) ||
                 (R[2*8 + 7] && R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[3][7][UP45P] = (!R[3*8 + 7] && !B[3*8 + 7]) && 

                 (
                 (R[3*8 + 6] && B[3*8 + 5]) ||
                 (R[3*8 + 6] && R[3*8 + 5] && B[3*8 + 4]) ||
                 (R[3*8 + 6] && R[3*8 + 5] && R[3*8 + 4] && B[3*8 + 3]) ||
                 (R[3*8 + 6] && R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && B[3*8 + 2]) ||
                 (R[3*8 + 6] && R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && B[3*8 + 1]) ||
                 (R[3*8 + 6] && R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && R[3*8 + 1] && B[3*8 + 0]) 
                 );
    M[4][7][ZEROP] = 1'b0;
    M[4][7][DOWN45P] = (!R[4*8 + 7] && !B[4*8 + 7]) && 

                 (
                 (R[5*8 + 6] && B[6*8 + 5]) ||
                 (R[5*8 + 6] && R[6*8 + 5] && B[7*8 + 4]) 
                 );
    M[4][7][DOWN] = (!R[4*8 + 7] && !B[4*8 + 7]) && 

                 (
                 (R[3*8 + 6] && B[2*8 + 5]) ||
                 (R[3*8 + 6] && R[2*8 + 5] && B[1*8 + 4]) ||
                 (R[3*8 + 6] && R[2*8 + 5] && R[1*8 + 4] && B[0*8 + 3]) 
                 );
    M[4][7][DOWN45M] = 1'b0;
    M[4][7][ZEROM] = 1'b0;
    M[4][7][UP45M] = (!R[4*8 + 7] && !B[4*8 + 7]) && 

                 (
                 (R[5*8 + 7] && B[6*8 + 7]) ||
                 (R[5*8 + 7] && R[6*8 + 7] && B[7*8 + 7]) 
                 );
    M[4][7][UP] = (!R[4*8 + 7] && !B[4*8 + 7]) && 

                 (
                 (R[3*8 + 7] && B[2*8 + 7]) ||
                 (R[3*8 + 7] && R[2*8 + 7] && B[1*8 + 7]) ||
                 (R[3*8 + 7] && R[2*8 + 7] && R[1*8 + 7] && B[0*8 + 7]) 
                 );
    M[4][7][UP45P] = (!R[4*8 + 7] && !B[4*8 + 7]) && 

                 (
                 (R[4*8 + 6] && B[4*8 + 5]) ||
                 (R[4*8 + 6] && R[4*8 + 5] && B[4*8 + 4]) ||
                 (R[4*8 + 6] && R[4*8 + 5] && R[4*8 + 4] && B[4*8 + 3]) ||
                 (R[4*8 + 6] && R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && B[4*8 + 2]) ||
                 (R[4*8 + 6] && R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && B[4*8 + 1]) ||
                 (R[4*8 + 6] && R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && R[4*8 + 1] && B[4*8 + 0]) 
                 );
    M[7][4][ZEROP] = 1'b0;
    M[7][4][DOWN45P] = 1'b0;
    M[7][4][DOWN] = (!R[7*8 + 4] && !B[7*8 + 4]) && 

                 (
                 (R[6*8 + 3] && B[5*8 + 2]) ||
                 (R[6*8 + 3] && R[5*8 + 2] && B[4*8 + 1]) ||
                 (R[6*8 + 3] && R[5*8 + 2] && R[4*8 + 1] && B[3*8 + 0]) 
                 );
    M[7][4][DOWN45M] = (!R[7*8 + 4] && !B[7*8 + 4]) && 

                 (
                 (R[6*8 + 5] && B[5*8 + 6]) ||
                 (R[6*8 + 5] && R[5*8 + 6] && B[4*8 + 7]) 
                 );
    M[7][4][ZEROM] = (!R[7*8 + 4] && !B[7*8 + 4]) && 

                 (
                 (R[7*8 + 5] && B[7*8 + 6]) ||
                 (R[7*8 + 5] && R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][4][UP45M] = 1'b0;
    M[7][4][UP] = (!R[7*8 + 4] && !B[7*8 + 4]) && 

                 (
                 (R[6*8 + 4] && B[5*8 + 4]) ||
                 (R[6*8 + 4] && R[5*8 + 4] && B[4*8 + 4]) ||
                 (R[6*8 + 4] && R[5*8 + 4] && R[4*8 + 4] && B[3*8 + 4]) ||
                 (R[6*8 + 4] && R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && B[2*8 + 4]) ||
                 (R[6*8 + 4] && R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && B[1*8 + 4]) ||
                 (R[6*8 + 4] && R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && R[1*8 + 4] && B[0*8 + 4]) 
                 );
    M[7][4][UP45P] = (!R[7*8 + 4] && !B[7*8 + 4]) && 

                 (
                 (R[7*8 + 3] && B[7*8 + 2]) ||
                 (R[7*8 + 3] && R[7*8 + 2] && B[7*8 + 1]) ||
                 (R[7*8 + 3] && R[7*8 + 2] && R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[7][3][ZEROP] = 1'b0;
    M[7][3][DOWN45P] = 1'b0;
    M[7][3][DOWN] = (!R[7*8 + 3] && !B[7*8 + 3]) && 

                 (
                 (R[6*8 + 2] && B[5*8 + 1]) ||
                 (R[6*8 + 2] && R[5*8 + 1] && B[4*8 + 0]) 
                 );
    M[7][3][DOWN45M] = (!R[7*8 + 3] && !B[7*8 + 3]) && 

                 (
                 (R[6*8 + 4] && B[5*8 + 5]) ||
                 (R[6*8 + 4] && R[5*8 + 5] && B[4*8 + 6]) ||
                 (R[6*8 + 4] && R[5*8 + 5] && R[4*8 + 6] && B[3*8 + 7]) 
                 );
    M[7][3][ZEROM] = (!R[7*8 + 3] && !B[7*8 + 3]) && 

                 (
                 (R[7*8 + 4] && B[7*8 + 5]) ||
                 (R[7*8 + 4] && R[7*8 + 5] && B[7*8 + 6]) ||
                 (R[7*8 + 4] && R[7*8 + 5] && R[7*8 + 6] && B[7*8 + 7]) 
                 );
    M[7][3][UP45M] = 1'b0;
    M[7][3][UP] = (!R[7*8 + 3] && !B[7*8 + 3]) && 

                 (
                 (R[6*8 + 3] && B[5*8 + 3]) ||
                 (R[6*8 + 3] && R[5*8 + 3] && B[4*8 + 3]) ||
                 (R[6*8 + 3] && R[5*8 + 3] && R[4*8 + 3] && B[3*8 + 3]) ||
                 (R[6*8 + 3] && R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && B[2*8 + 3]) ||
                 (R[6*8 + 3] && R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && B[1*8 + 3]) ||
                 (R[6*8 + 3] && R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && R[1*8 + 3] && B[0*8 + 3]) 
                 );
    M[7][3][UP45P] = (!R[7*8 + 3] && !B[7*8 + 3]) && 

                 (
                 (R[7*8 + 2] && B[7*8 + 1]) ||
                 (R[7*8 + 2] && R[7*8 + 1] && B[7*8 + 0]) 
                 );
    M[4][0][ZEROP] = (!R[4*8 + 0] && !B[4*8 + 0]) && 

                 (
                 (R[5*8 + 1] && B[6*8 + 2]) ||
                 (R[5*8 + 1] && R[6*8 + 2] && B[7*8 + 3]) 
                 );
    M[4][0][DOWN45P] = 1'b0;
    M[4][0][DOWN] = 1'b0;
    M[4][0][DOWN45M] = (!R[4*8 + 0] && !B[4*8 + 0]) && 

                 (
                 (R[3*8 + 1] && B[2*8 + 2]) ||
                 (R[3*8 + 1] && R[2*8 + 2] && B[1*8 + 3]) ||
                 (R[3*8 + 1] && R[2*8 + 2] && R[1*8 + 3] && B[0*8 + 4]) 
                 );
    M[4][0][ZEROM] = (!R[4*8 + 0] && !B[4*8 + 0]) && 

                 (
                 (R[4*8 + 1] && B[4*8 + 2]) ||
                 (R[4*8 + 1] && R[4*8 + 2] && B[4*8 + 3]) ||
                 (R[4*8 + 1] && R[4*8 + 2] && R[4*8 + 3] && B[4*8 + 4]) ||
                 (R[4*8 + 1] && R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && B[4*8 + 5]) ||
                 (R[4*8 + 1] && R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && B[4*8 + 6]) ||
                 (R[4*8 + 1] && R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && R[4*8 + 6] && B[4*8 + 7]) 
                 );
    M[4][0][UP45M] = (!R[4*8 + 0] && !B[4*8 + 0]) && 

                 (
                 (R[5*8 + 0] && B[6*8 + 0]) ||
                 (R[5*8 + 0] && R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[4][0][UP] = (!R[4*8 + 0] && !B[4*8 + 0]) && 

                 (
                 (R[3*8 + 0] && B[2*8 + 0]) ||
                 (R[3*8 + 0] && R[2*8 + 0] && B[1*8 + 0]) ||
                 (R[3*8 + 0] && R[2*8 + 0] && R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[4][0][UP45P] = 1'b0;
    M[3][0][ZEROP] = (!R[3*8 + 0] && !B[3*8 + 0]) && 

                 (
                 (R[4*8 + 1] && B[5*8 + 2]) ||
                 (R[4*8 + 1] && R[5*8 + 2] && B[6*8 + 3]) ||
                 (R[4*8 + 1] && R[5*8 + 2] && R[6*8 + 3] && B[7*8 + 4]) 
                 );
    M[3][0][DOWN45P] = 1'b0;
    M[3][0][DOWN] = 1'b0;
    M[3][0][DOWN45M] = (!R[3*8 + 0] && !B[3*8 + 0]) && 

                 (
                 (R[2*8 + 1] && B[1*8 + 2]) ||
                 (R[2*8 + 1] && R[1*8 + 2] && B[0*8 + 3]) 
                 );
    M[3][0][ZEROM] = (!R[3*8 + 0] && !B[3*8 + 0]) && 

                 (
                 (R[3*8 + 1] && B[3*8 + 2]) ||
                 (R[3*8 + 1] && R[3*8 + 2] && B[3*8 + 3]) ||
                 (R[3*8 + 1] && R[3*8 + 2] && R[3*8 + 3] && B[3*8 + 4]) ||
                 (R[3*8 + 1] && R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && B[3*8 + 5]) ||
                 (R[3*8 + 1] && R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && B[3*8 + 6]) ||
                 (R[3*8 + 1] && R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && R[3*8 + 6] && B[3*8 + 7]) 
                 );
    M[3][0][UP45M] = (!R[3*8 + 0] && !B[3*8 + 0]) && 

                 (
                 (R[4*8 + 0] && B[5*8 + 0]) ||
                 (R[4*8 + 0] && R[5*8 + 0] && B[6*8 + 0]) ||
                 (R[4*8 + 0] && R[5*8 + 0] && R[6*8 + 0] && B[7*8 + 0]) 
                 );
    M[3][0][UP] = (!R[3*8 + 0] && !B[3*8 + 0]) && 

                 (
                 (R[2*8 + 0] && B[1*8 + 0]) ||
                 (R[2*8 + 0] && R[1*8 + 0] && B[0*8 + 0]) 
                 );
    M[3][0][UP45P] = 1'b0;


// Expresii generate pentru patrate E
    M[1][1][ZEROP] = (!R[1*8 + 1] && !B[1*8 + 1]) && 

                 (
                 (R[2*8 + 2] && B[3*8 + 3]) ||
                 (R[2*8 + 2] && R[3*8 + 3] && B[4*8 + 4]) ||
                 (R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && B[5*8 + 5]) ||
                 (R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && B[6*8 + 6]) ||
                 (R[2*8 + 2] && R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && R[6*8 + 6] && B[7*8 + 7]) 
                 );
    M[1][1][DOWN45P] = 1'b0;
    M[1][1][DOWN] = 1'b0;
    M[1][1][DOWN45M] = 1'b0;
    M[1][1][ZEROM] = (!R[1*8 + 1] && !B[1*8 + 1]) && 

                 (
                 (R[1*8 + 2] && B[1*8 + 3]) ||
                 (R[1*8 + 2] && R[1*8 + 3] && B[1*8 + 4]) ||
                 (R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && B[1*8 + 5]) ||
                 (R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && B[1*8 + 6]) ||
                 (R[1*8 + 2] && R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][1][UP45M] = (!R[1*8 + 1] && !B[1*8 + 1]) && 

                 (
                 (R[2*8 + 1] && B[3*8 + 1]) ||
                 (R[2*8 + 1] && R[3*8 + 1] && B[4*8 + 1]) ||
                 (R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && B[5*8 + 1]) ||
                 (R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && B[6*8 + 1]) ||
                 (R[2*8 + 1] && R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[1][1][UP] = 1'b0;
    M[1][1][UP45P] = 1'b0;
    M[1][6][ZEROP] = 1'b0;
    M[1][6][DOWN45P] = (!R[1*8 + 6] && !B[1*8 + 6]) && 

                 (
                 (R[2*8 + 5] && B[3*8 + 4]) ||
                 (R[2*8 + 5] && R[3*8 + 4] && B[4*8 + 3]) ||
                 (R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && B[5*8 + 2]) ||
                 (R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && B[6*8 + 1]) ||
                 (R[2*8 + 5] && R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && R[6*8 + 1] && B[7*8 + 0]) 
                 );
    M[1][6][DOWN] = 1'b0;
    M[1][6][DOWN45M] = 1'b0;
    M[1][6][ZEROM] = 1'b0;
    M[1][6][UP45M] = (!R[1*8 + 6] && !B[1*8 + 6]) && 

                 (
                 (R[2*8 + 6] && B[3*8 + 6]) ||
                 (R[2*8 + 6] && R[3*8 + 6] && B[4*8 + 6]) ||
                 (R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && B[5*8 + 6]) ||
                 (R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && B[6*8 + 6]) ||
                 (R[2*8 + 6] && R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[1][6][UP] = 1'b0;
    M[1][6][UP45P] = (!R[1*8 + 6] && !B[1*8 + 6]) && 

                 (
                 (R[1*8 + 5] && B[1*8 + 4]) ||
                 (R[1*8 + 5] && R[1*8 + 4] && B[1*8 + 3]) ||
                 (R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && B[1*8 + 2]) ||
                 (R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && B[1*8 + 1]) ||
                 (R[1*8 + 5] && R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[6][6][ZEROP] = 1'b0;
    M[6][6][DOWN45P] = 1'b0;
    M[6][6][DOWN] = (!R[6*8 + 6] && !B[6*8 + 6]) && 

                 (
                 (R[5*8 + 5] && B[4*8 + 4]) ||
                 (R[5*8 + 5] && R[4*8 + 4] && B[3*8 + 3]) ||
                 (R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && B[2*8 + 2]) ||
                 (R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && B[1*8 + 1]) ||
                 (R[5*8 + 5] && R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && R[1*8 + 1] && B[0*8 + 0]) 
                 );
    M[6][6][DOWN45M] = 1'b0;
    M[6][6][ZEROM] = 1'b0;
    M[6][6][UP45M] = 1'b0;
    M[6][6][UP] = (!R[6*8 + 6] && !B[6*8 + 6]) && 

                 (
                 (R[5*8 + 6] && B[4*8 + 6]) ||
                 (R[5*8 + 6] && R[4*8 + 6] && B[3*8 + 6]) ||
                 (R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && B[2*8 + 6]) ||
                 (R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && B[1*8 + 6]) ||
                 (R[5*8 + 6] && R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[6][6][UP45P] = (!R[6*8 + 6] && !B[6*8 + 6]) && 

                 (
                 (R[6*8 + 5] && B[6*8 + 4]) ||
                 (R[6*8 + 5] && R[6*8 + 4] && B[6*8 + 3]) ||
                 (R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && B[6*8 + 2]) ||
                 (R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && B[6*8 + 1]) ||
                 (R[6*8 + 5] && R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[6][1][ZEROP] = 1'b0;
    M[6][1][DOWN45P] = 1'b0;
    M[6][1][DOWN] = 1'b0;
    M[6][1][DOWN45M] = (!R[6*8 + 1] && !B[6*8 + 1]) && 

                 (
                 (R[5*8 + 2] && B[4*8 + 3]) ||
                 (R[5*8 + 2] && R[4*8 + 3] && B[3*8 + 4]) ||
                 (R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && B[2*8 + 5]) ||
                 (R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && B[1*8 + 6]) ||
                 (R[5*8 + 2] && R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && R[1*8 + 6] && B[0*8 + 7]) 
                 );
    M[6][1][ZEROM] = (!R[6*8 + 1] && !B[6*8 + 1]) && 

                 (
                 (R[6*8 + 2] && B[6*8 + 3]) ||
                 (R[6*8 + 2] && R[6*8 + 3] && B[6*8 + 4]) ||
                 (R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && B[6*8 + 5]) ||
                 (R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && B[6*8 + 6]) ||
                 (R[6*8 + 2] && R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][1][UP45M] = 1'b0;
    M[6][1][UP] = (!R[6*8 + 1] && !B[6*8 + 1]) && 

                 (
                 (R[5*8 + 1] && B[4*8 + 1]) ||
                 (R[5*8 + 1] && R[4*8 + 1] && B[3*8 + 1]) ||
                 (R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && B[2*8 + 1]) ||
                 (R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && B[1*8 + 1]) ||
                 (R[5*8 + 1] && R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[6][1][UP45P] = 1'b0;


// Expresii generate pentru patrate F
    M[1][2][ZEROP] = (!R[1*8 + 2] && !B[1*8 + 2]) && 

                 (
                 (R[2*8 + 3] && B[3*8 + 4]) ||
                 (R[2*8 + 3] && R[3*8 + 4] && B[4*8 + 5]) ||
                 (R[2*8 + 3] && R[3*8 + 4] && R[4*8 + 5] && B[5*8 + 6]) ||
                 (R[2*8 + 3] && R[3*8 + 4] && R[4*8 + 5] && R[5*8 + 6] && B[6*8 + 7]) 
                 );
    M[1][2][DOWN45P] = (!R[1*8 + 2] && !B[1*8 + 2]) && 

                 (
                 (R[2*8 + 1] && B[3*8 + 0]) 
                 );
    M[1][2][DOWN] = 1'b0;
    M[1][2][DOWN45M] = 1'b0;
    M[1][2][ZEROM] = (!R[1*8 + 2] && !B[1*8 + 2]) && 

                 (
                 (R[1*8 + 3] && B[1*8 + 4]) ||
                 (R[1*8 + 3] && R[1*8 + 4] && B[1*8 + 5]) ||
                 (R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && B[1*8 + 6]) ||
                 (R[1*8 + 3] && R[1*8 + 4] && R[1*8 + 5] && R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][2][UP45M] = (!R[1*8 + 2] && !B[1*8 + 2]) && 

                 (
                 (R[2*8 + 2] && B[3*8 + 2]) ||
                 (R[2*8 + 2] && R[3*8 + 2] && B[4*8 + 2]) ||
                 (R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && B[5*8 + 2]) ||
                 (R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && B[6*8 + 2]) ||
                 (R[2*8 + 2] && R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[1][2][UP] = 1'b0;
    M[1][2][UP45P] = (!R[1*8 + 2] && !B[1*8 + 2]) && 

                 (
                 (R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[1][5][ZEROP] = (!R[1*8 + 5] && !B[1*8 + 5]) && 

                 (
                 (R[2*8 + 6] && B[3*8 + 7]) 
                 );
    M[1][5][DOWN45P] = (!R[1*8 + 5] && !B[1*8 + 5]) && 

                 (
                 (R[2*8 + 4] && B[3*8 + 3]) ||
                 (R[2*8 + 4] && R[3*8 + 3] && B[4*8 + 2]) ||
                 (R[2*8 + 4] && R[3*8 + 3] && R[4*8 + 2] && B[5*8 + 1]) ||
                 (R[2*8 + 4] && R[3*8 + 3] && R[4*8 + 2] && R[5*8 + 1] && B[6*8 + 0]) 
                 );
    M[1][5][DOWN] = 1'b0;
    M[1][5][DOWN45M] = 1'b0;
    M[1][5][ZEROM] = (!R[1*8 + 5] && !B[1*8 + 5]) && 

                 (
                 (R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][5][UP45M] = (!R[1*8 + 5] && !B[1*8 + 5]) && 

                 (
                 (R[2*8 + 5] && B[3*8 + 5]) ||
                 (R[2*8 + 5] && R[3*8 + 5] && B[4*8 + 5]) ||
                 (R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && B[5*8 + 5]) ||
                 (R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && B[6*8 + 5]) ||
                 (R[2*8 + 5] && R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[1][5][UP] = 1'b0;
    M[1][5][UP45P] = (!R[1*8 + 5] && !B[1*8 + 5]) && 

                 (
                 (R[1*8 + 4] && B[1*8 + 3]) ||
                 (R[1*8 + 4] && R[1*8 + 3] && B[1*8 + 2]) ||
                 (R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && B[1*8 + 1]) ||
                 (R[1*8 + 4] && R[1*8 + 3] && R[1*8 + 2] && R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[2][6][ZEROP] = 1'b0;
    M[2][6][DOWN45P] = (!R[2*8 + 6] && !B[2*8 + 6]) && 

                 (
                 (R[3*8 + 5] && B[4*8 + 4]) ||
                 (R[3*8 + 5] && R[4*8 + 4] && B[5*8 + 3]) ||
                 (R[3*8 + 5] && R[4*8 + 4] && R[5*8 + 3] && B[6*8 + 2]) ||
                 (R[3*8 + 5] && R[4*8 + 4] && R[5*8 + 3] && R[6*8 + 2] && B[7*8 + 1]) 
                 );
    M[2][6][DOWN] = (!R[2*8 + 6] && !B[2*8 + 6]) && 

                 (
                 (R[1*8 + 5] && B[0*8 + 4]) 
                 );
    M[2][6][DOWN45M] = 1'b0;
    M[2][6][ZEROM] = 1'b0;
    M[2][6][UP45M] = (!R[2*8 + 6] && !B[2*8 + 6]) && 

                 (
                 (R[3*8 + 6] && B[4*8 + 6]) ||
                 (R[3*8 + 6] && R[4*8 + 6] && B[5*8 + 6]) ||
                 (R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && B[6*8 + 6]) ||
                 (R[3*8 + 6] && R[4*8 + 6] && R[5*8 + 6] && R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[2][6][UP] = (!R[2*8 + 6] && !B[2*8 + 6]) && 

                 (
                 (R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[2][6][UP45P] = (!R[2*8 + 6] && !B[2*8 + 6]) && 

                 (
                 (R[2*8 + 5] && B[2*8 + 4]) ||
                 (R[2*8 + 5] && R[2*8 + 4] && B[2*8 + 3]) ||
                 (R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && B[2*8 + 2]) ||
                 (R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && B[2*8 + 1]) ||
                 (R[2*8 + 5] && R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[5][6][ZEROP] = 1'b0;
    M[5][6][DOWN45P] = (!R[5*8 + 6] && !B[5*8 + 6]) && 

                 (
                 (R[6*8 + 5] && B[7*8 + 4]) 
                 );
    M[5][6][DOWN] = (!R[5*8 + 6] && !B[5*8 + 6]) && 

                 (
                 (R[4*8 + 5] && B[3*8 + 4]) ||
                 (R[4*8 + 5] && R[3*8 + 4] && B[2*8 + 3]) ||
                 (R[4*8 + 5] && R[3*8 + 4] && R[2*8 + 3] && B[1*8 + 2]) ||
                 (R[4*8 + 5] && R[3*8 + 4] && R[2*8 + 3] && R[1*8 + 2] && B[0*8 + 1]) 
                 );
    M[5][6][DOWN45M] = 1'b0;
    M[5][6][ZEROM] = 1'b0;
    M[5][6][UP45M] = (!R[5*8 + 6] && !B[5*8 + 6]) && 

                 (
                 (R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[5][6][UP] = (!R[5*8 + 6] && !B[5*8 + 6]) && 

                 (
                 (R[4*8 + 6] && B[3*8 + 6]) ||
                 (R[4*8 + 6] && R[3*8 + 6] && B[2*8 + 6]) ||
                 (R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && B[1*8 + 6]) ||
                 (R[4*8 + 6] && R[3*8 + 6] && R[2*8 + 6] && R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[5][6][UP45P] = (!R[5*8 + 6] && !B[5*8 + 6]) && 

                 (
                 (R[5*8 + 5] && B[5*8 + 4]) ||
                 (R[5*8 + 5] && R[5*8 + 4] && B[5*8 + 3]) ||
                 (R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && B[5*8 + 2]) ||
                 (R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && B[5*8 + 1]) ||
                 (R[5*8 + 5] && R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && R[5*8 + 1] && B[5*8 + 0]) 
                 );
    M[6][5][ZEROP] = 1'b0;
    M[6][5][DOWN45P] = 1'b0;
    M[6][5][DOWN] = (!R[6*8 + 5] && !B[6*8 + 5]) && 

                 (
                 (R[5*8 + 4] && B[4*8 + 3]) ||
                 (R[5*8 + 4] && R[4*8 + 3] && B[3*8 + 2]) ||
                 (R[5*8 + 4] && R[4*8 + 3] && R[3*8 + 2] && B[2*8 + 1]) ||
                 (R[5*8 + 4] && R[4*8 + 3] && R[3*8 + 2] && R[2*8 + 1] && B[1*8 + 0]) 
                 );
    M[6][5][DOWN45M] = (!R[6*8 + 5] && !B[6*8 + 5]) && 

                 (
                 (R[5*8 + 6] && B[4*8 + 7]) 
                 );
    M[6][5][ZEROM] = (!R[6*8 + 5] && !B[6*8 + 5]) && 

                 (
                 (R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][5][UP45M] = 1'b0;
    M[6][5][UP] = (!R[6*8 + 5] && !B[6*8 + 5]) && 

                 (
                 (R[5*8 + 5] && B[4*8 + 5]) ||
                 (R[5*8 + 5] && R[4*8 + 5] && B[3*8 + 5]) ||
                 (R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && B[2*8 + 5]) ||
                 (R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && B[1*8 + 5]) ||
                 (R[5*8 + 5] && R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[6][5][UP45P] = (!R[6*8 + 5] && !B[6*8 + 5]) && 

                 (
                 (R[6*8 + 4] && B[6*8 + 3]) ||
                 (R[6*8 + 4] && R[6*8 + 3] && B[6*8 + 2]) ||
                 (R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && B[6*8 + 1]) ||
                 (R[6*8 + 4] && R[6*8 + 3] && R[6*8 + 2] && R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[6][2][ZEROP] = 1'b0;
    M[6][2][DOWN45P] = 1'b0;
    M[6][2][DOWN] = (!R[6*8 + 2] && !B[6*8 + 2]) && 

                 (
                 (R[5*8 + 1] && B[4*8 + 0]) 
                 );
    M[6][2][DOWN45M] = (!R[6*8 + 2] && !B[6*8 + 2]) && 

                 (
                 (R[5*8 + 3] && B[4*8 + 4]) ||
                 (R[5*8 + 3] && R[4*8 + 4] && B[3*8 + 5]) ||
                 (R[5*8 + 3] && R[4*8 + 4] && R[3*8 + 5] && B[2*8 + 6]) ||
                 (R[5*8 + 3] && R[4*8 + 4] && R[3*8 + 5] && R[2*8 + 6] && B[1*8 + 7]) 
                 );
    M[6][2][ZEROM] = (!R[6*8 + 2] && !B[6*8 + 2]) && 

                 (
                 (R[6*8 + 3] && B[6*8 + 4]) ||
                 (R[6*8 + 3] && R[6*8 + 4] && B[6*8 + 5]) ||
                 (R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && B[6*8 + 6]) ||
                 (R[6*8 + 3] && R[6*8 + 4] && R[6*8 + 5] && R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][2][UP45M] = 1'b0;
    M[6][2][UP] = (!R[6*8 + 2] && !B[6*8 + 2]) && 

                 (
                 (R[5*8 + 2] && B[4*8 + 2]) ||
                 (R[5*8 + 2] && R[4*8 + 2] && B[3*8 + 2]) ||
                 (R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && B[2*8 + 2]) ||
                 (R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && B[1*8 + 2]) ||
                 (R[5*8 + 2] && R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[6][2][UP45P] = (!R[6*8 + 2] && !B[6*8 + 2]) && 

                 (
                 (R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[5][1][ZEROP] = (!R[5*8 + 1] && !B[5*8 + 1]) && 

                 (
                 (R[6*8 + 2] && B[7*8 + 3]) 
                 );
    M[5][1][DOWN45P] = 1'b0;
    M[5][1][DOWN] = 1'b0;
    M[5][1][DOWN45M] = (!R[5*8 + 1] && !B[5*8 + 1]) && 

                 (
                 (R[4*8 + 2] && B[3*8 + 3]) ||
                 (R[4*8 + 2] && R[3*8 + 3] && B[2*8 + 4]) ||
                 (R[4*8 + 2] && R[3*8 + 3] && R[2*8 + 4] && B[1*8 + 5]) ||
                 (R[4*8 + 2] && R[3*8 + 3] && R[2*8 + 4] && R[1*8 + 5] && B[0*8 + 6]) 
                 );
    M[5][1][ZEROM] = (!R[5*8 + 1] && !B[5*8 + 1]) && 

                 (
                 (R[5*8 + 2] && B[5*8 + 3]) ||
                 (R[5*8 + 2] && R[5*8 + 3] && B[5*8 + 4]) ||
                 (R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && B[5*8 + 5]) ||
                 (R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && B[5*8 + 6]) ||
                 (R[5*8 + 2] && R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][1][UP45M] = (!R[5*8 + 1] && !B[5*8 + 1]) && 

                 (
                 (R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[5][1][UP] = (!R[5*8 + 1] && !B[5*8 + 1]) && 

                 (
                 (R[4*8 + 1] && B[3*8 + 1]) ||
                 (R[4*8 + 1] && R[3*8 + 1] && B[2*8 + 1]) ||
                 (R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && B[1*8 + 1]) ||
                 (R[4*8 + 1] && R[3*8 + 1] && R[2*8 + 1] && R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[5][1][UP45P] = 1'b0;
    M[2][1][ZEROP] = (!R[2*8 + 1] && !B[2*8 + 1]) && 

                 (
                 (R[3*8 + 2] && B[4*8 + 3]) ||
                 (R[3*8 + 2] && R[4*8 + 3] && B[5*8 + 4]) ||
                 (R[3*8 + 2] && R[4*8 + 3] && R[5*8 + 4] && B[6*8 + 5]) ||
                 (R[3*8 + 2] && R[4*8 + 3] && R[5*8 + 4] && R[6*8 + 5] && B[7*8 + 6]) 
                 );
    M[2][1][DOWN45P] = 1'b0;
    M[2][1][DOWN] = 1'b0;
    M[2][1][DOWN45M] = (!R[2*8 + 1] && !B[2*8 + 1]) && 

                 (
                 (R[1*8 + 2] && B[0*8 + 3]) 
                 );
    M[2][1][ZEROM] = (!R[2*8 + 1] && !B[2*8 + 1]) && 

                 (
                 (R[2*8 + 2] && B[2*8 + 3]) ||
                 (R[2*8 + 2] && R[2*8 + 3] && B[2*8 + 4]) ||
                 (R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && B[2*8 + 5]) ||
                 (R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && B[2*8 + 6]) ||
                 (R[2*8 + 2] && R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][1][UP45M] = (!R[2*8 + 1] && !B[2*8 + 1]) && 

                 (
                 (R[3*8 + 1] && B[4*8 + 1]) ||
                 (R[3*8 + 1] && R[4*8 + 1] && B[5*8 + 1]) ||
                 (R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && B[6*8 + 1]) ||
                 (R[3*8 + 1] && R[4*8 + 1] && R[5*8 + 1] && R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[2][1][UP] = (!R[2*8 + 1] && !B[2*8 + 1]) && 

                 (
                 (R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[2][1][UP45P] = 1'b0;


// Expresii generate pentru patrate G
    M[1][3][ZEROP] = (!R[1*8 + 3] && !B[1*8 + 3]) && 

                 (
                 (R[2*8 + 4] && B[3*8 + 5]) ||
                 (R[2*8 + 4] && R[3*8 + 5] && B[4*8 + 6]) ||
                 (R[2*8 + 4] && R[3*8 + 5] && R[4*8 + 6] && B[5*8 + 7]) 
                 );
    M[1][3][DOWN45P] = (!R[1*8 + 3] && !B[1*8 + 3]) && 

                 (
                 (R[2*8 + 2] && B[3*8 + 1]) ||
                 (R[2*8 + 2] && R[3*8 + 1] && B[4*8 + 0]) 
                 );
    M[1][3][DOWN] = 1'b0;
    M[1][3][DOWN45M] = 1'b0;
    M[1][3][ZEROM] = (!R[1*8 + 3] && !B[1*8 + 3]) && 

                 (
                 (R[1*8 + 4] && B[1*8 + 5]) ||
                 (R[1*8 + 4] && R[1*8 + 5] && B[1*8 + 6]) ||
                 (R[1*8 + 4] && R[1*8 + 5] && R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][3][UP45M] = (!R[1*8 + 3] && !B[1*8 + 3]) && 

                 (
                 (R[2*8 + 3] && B[3*8 + 3]) ||
                 (R[2*8 + 3] && R[3*8 + 3] && B[4*8 + 3]) ||
                 (R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && B[5*8 + 3]) ||
                 (R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && B[6*8 + 3]) ||
                 (R[2*8 + 3] && R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && R[6*8 + 3] && B[7*8 + 3]) 
                 );
    M[1][3][UP] = 1'b0;
    M[1][3][UP45P] = (!R[1*8 + 3] && !B[1*8 + 3]) && 

                 (
                 (R[1*8 + 2] && B[1*8 + 1]) ||
                 (R[1*8 + 2] && R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[1][4][ZEROP] = (!R[1*8 + 4] && !B[1*8 + 4]) && 

                 (
                 (R[2*8 + 5] && B[3*8 + 6]) ||
                 (R[2*8 + 5] && R[3*8 + 6] && B[4*8 + 7]) 
                 );
    M[1][4][DOWN45P] = (!R[1*8 + 4] && !B[1*8 + 4]) && 

                 (
                 (R[2*8 + 3] && B[3*8 + 2]) ||
                 (R[2*8 + 3] && R[3*8 + 2] && B[4*8 + 1]) ||
                 (R[2*8 + 3] && R[3*8 + 2] && R[4*8 + 1] && B[5*8 + 0]) 
                 );
    M[1][4][DOWN] = 1'b0;
    M[1][4][DOWN45M] = 1'b0;
    M[1][4][ZEROM] = (!R[1*8 + 4] && !B[1*8 + 4]) && 

                 (
                 (R[1*8 + 5] && B[1*8 + 6]) ||
                 (R[1*8 + 5] && R[1*8 + 6] && B[1*8 + 7]) 
                 );
    M[1][4][UP45M] = (!R[1*8 + 4] && !B[1*8 + 4]) && 

                 (
                 (R[2*8 + 4] && B[3*8 + 4]) ||
                 (R[2*8 + 4] && R[3*8 + 4] && B[4*8 + 4]) ||
                 (R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && B[5*8 + 4]) ||
                 (R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && B[6*8 + 4]) ||
                 (R[2*8 + 4] && R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && R[6*8 + 4] && B[7*8 + 4]) 
                 );
    M[1][4][UP] = 1'b0;
    M[1][4][UP45P] = (!R[1*8 + 4] && !B[1*8 + 4]) && 

                 (
                 (R[1*8 + 3] && B[1*8 + 2]) ||
                 (R[1*8 + 3] && R[1*8 + 2] && B[1*8 + 1]) ||
                 (R[1*8 + 3] && R[1*8 + 2] && R[1*8 + 1] && B[1*8 + 0]) 
                 );
    M[3][6][ZEROP] = 1'b0;
    M[3][6][DOWN45P] = (!R[3*8 + 6] && !B[3*8 + 6]) && 

                 (
                 (R[4*8 + 5] && B[5*8 + 4]) ||
                 (R[4*8 + 5] && R[5*8 + 4] && B[6*8 + 3]) ||
                 (R[4*8 + 5] && R[5*8 + 4] && R[6*8 + 3] && B[7*8 + 2]) 
                 );
    M[3][6][DOWN] = (!R[3*8 + 6] && !B[3*8 + 6]) && 

                 (
                 (R[2*8 + 5] && B[1*8 + 4]) ||
                 (R[2*8 + 5] && R[1*8 + 4] && B[0*8 + 3]) 
                 );
    M[3][6][DOWN45M] = 1'b0;
    M[3][6][ZEROM] = 1'b0;
    M[3][6][UP45M] = (!R[3*8 + 6] && !B[3*8 + 6]) && 

                 (
                 (R[4*8 + 6] && B[5*8 + 6]) ||
                 (R[4*8 + 6] && R[5*8 + 6] && B[6*8 + 6]) ||
                 (R[4*8 + 6] && R[5*8 + 6] && R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[3][6][UP] = (!R[3*8 + 6] && !B[3*8 + 6]) && 

                 (
                 (R[2*8 + 6] && B[1*8 + 6]) ||
                 (R[2*8 + 6] && R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[3][6][UP45P] = (!R[3*8 + 6] && !B[3*8 + 6]) && 

                 (
                 (R[3*8 + 5] && B[3*8 + 4]) ||
                 (R[3*8 + 5] && R[3*8 + 4] && B[3*8 + 3]) ||
                 (R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && B[3*8 + 2]) ||
                 (R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && B[3*8 + 1]) ||
                 (R[3*8 + 5] && R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && R[3*8 + 1] && B[3*8 + 0]) 
                 );
    M[4][6][ZEROP] = 1'b0;
    M[4][6][DOWN45P] = (!R[4*8 + 6] && !B[4*8 + 6]) && 

                 (
                 (R[5*8 + 5] && B[6*8 + 4]) ||
                 (R[5*8 + 5] && R[6*8 + 4] && B[7*8 + 3]) 
                 );
    M[4][6][DOWN] = (!R[4*8 + 6] && !B[4*8 + 6]) && 

                 (
                 (R[3*8 + 5] && B[2*8 + 4]) ||
                 (R[3*8 + 5] && R[2*8 + 4] && B[1*8 + 3]) ||
                 (R[3*8 + 5] && R[2*8 + 4] && R[1*8 + 3] && B[0*8 + 2]) 
                 );
    M[4][6][DOWN45M] = 1'b0;
    M[4][6][ZEROM] = 1'b0;
    M[4][6][UP45M] = (!R[4*8 + 6] && !B[4*8 + 6]) && 

                 (
                 (R[5*8 + 6] && B[6*8 + 6]) ||
                 (R[5*8 + 6] && R[6*8 + 6] && B[7*8 + 6]) 
                 );
    M[4][6][UP] = (!R[4*8 + 6] && !B[4*8 + 6]) && 

                 (
                 (R[3*8 + 6] && B[2*8 + 6]) ||
                 (R[3*8 + 6] && R[2*8 + 6] && B[1*8 + 6]) ||
                 (R[3*8 + 6] && R[2*8 + 6] && R[1*8 + 6] && B[0*8 + 6]) 
                 );
    M[4][6][UP45P] = (!R[4*8 + 6] && !B[4*8 + 6]) && 

                 (
                 (R[4*8 + 5] && B[4*8 + 4]) ||
                 (R[4*8 + 5] && R[4*8 + 4] && B[4*8 + 3]) ||
                 (R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && B[4*8 + 2]) ||
                 (R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && B[4*8 + 1]) ||
                 (R[4*8 + 5] && R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && R[4*8 + 1] && B[4*8 + 0]) 
                 );
    M[6][4][ZEROP] = 1'b0;
    M[6][4][DOWN45P] = 1'b0;
    M[6][4][DOWN] = (!R[6*8 + 4] && !B[6*8 + 4]) && 

                 (
                 (R[5*8 + 3] && B[4*8 + 2]) ||
                 (R[5*8 + 3] && R[4*8 + 2] && B[3*8 + 1]) ||
                 (R[5*8 + 3] && R[4*8 + 2] && R[3*8 + 1] && B[2*8 + 0]) 
                 );
    M[6][4][DOWN45M] = (!R[6*8 + 4] && !B[6*8 + 4]) && 

                 (
                 (R[5*8 + 5] && B[4*8 + 6]) ||
                 (R[5*8 + 5] && R[4*8 + 6] && B[3*8 + 7]) 
                 );
    M[6][4][ZEROM] = (!R[6*8 + 4] && !B[6*8 + 4]) && 

                 (
                 (R[6*8 + 5] && B[6*8 + 6]) ||
                 (R[6*8 + 5] && R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][4][UP45M] = 1'b0;
    M[6][4][UP] = (!R[6*8 + 4] && !B[6*8 + 4]) && 

                 (
                 (R[5*8 + 4] && B[4*8 + 4]) ||
                 (R[5*8 + 4] && R[4*8 + 4] && B[3*8 + 4]) ||
                 (R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && B[2*8 + 4]) ||
                 (R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && B[1*8 + 4]) ||
                 (R[5*8 + 4] && R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && R[1*8 + 4] && B[0*8 + 4]) 
                 );
    M[6][4][UP45P] = (!R[6*8 + 4] && !B[6*8 + 4]) && 

                 (
                 (R[6*8 + 3] && B[6*8 + 2]) ||
                 (R[6*8 + 3] && R[6*8 + 2] && B[6*8 + 1]) ||
                 (R[6*8 + 3] && R[6*8 + 2] && R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[6][3][ZEROP] = 1'b0;
    M[6][3][DOWN45P] = 1'b0;
    M[6][3][DOWN] = (!R[6*8 + 3] && !B[6*8 + 3]) && 

                 (
                 (R[5*8 + 2] && B[4*8 + 1]) ||
                 (R[5*8 + 2] && R[4*8 + 1] && B[3*8 + 0]) 
                 );
    M[6][3][DOWN45M] = (!R[6*8 + 3] && !B[6*8 + 3]) && 

                 (
                 (R[5*8 + 4] && B[4*8 + 5]) ||
                 (R[5*8 + 4] && R[4*8 + 5] && B[3*8 + 6]) ||
                 (R[5*8 + 4] && R[4*8 + 5] && R[3*8 + 6] && B[2*8 + 7]) 
                 );
    M[6][3][ZEROM] = (!R[6*8 + 3] && !B[6*8 + 3]) && 

                 (
                 (R[6*8 + 4] && B[6*8 + 5]) ||
                 (R[6*8 + 4] && R[6*8 + 5] && B[6*8 + 6]) ||
                 (R[6*8 + 4] && R[6*8 + 5] && R[6*8 + 6] && B[6*8 + 7]) 
                 );
    M[6][3][UP45M] = 1'b0;
    M[6][3][UP] = (!R[6*8 + 3] && !B[6*8 + 3]) && 

                 (
                 (R[5*8 + 3] && B[4*8 + 3]) ||
                 (R[5*8 + 3] && R[4*8 + 3] && B[3*8 + 3]) ||
                 (R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && B[2*8 + 3]) ||
                 (R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && B[1*8 + 3]) ||
                 (R[5*8 + 3] && R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && R[1*8 + 3] && B[0*8 + 3]) 
                 );
    M[6][3][UP45P] = (!R[6*8 + 3] && !B[6*8 + 3]) && 

                 (
                 (R[6*8 + 2] && B[6*8 + 1]) ||
                 (R[6*8 + 2] && R[6*8 + 1] && B[6*8 + 0]) 
                 );
    M[4][1][ZEROP] = (!R[4*8 + 1] && !B[4*8 + 1]) && 

                 (
                 (R[5*8 + 2] && B[6*8 + 3]) ||
                 (R[5*8 + 2] && R[6*8 + 3] && B[7*8 + 4]) 
                 );
    M[4][1][DOWN45P] = 1'b0;
    M[4][1][DOWN] = 1'b0;
    M[4][1][DOWN45M] = (!R[4*8 + 1] && !B[4*8 + 1]) && 

                 (
                 (R[3*8 + 2] && B[2*8 + 3]) ||
                 (R[3*8 + 2] && R[2*8 + 3] && B[1*8 + 4]) ||
                 (R[3*8 + 2] && R[2*8 + 3] && R[1*8 + 4] && B[0*8 + 5]) 
                 );
    M[4][1][ZEROM] = (!R[4*8 + 1] && !B[4*8 + 1]) && 

                 (
                 (R[4*8 + 2] && B[4*8 + 3]) ||
                 (R[4*8 + 2] && R[4*8 + 3] && B[4*8 + 4]) ||
                 (R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && B[4*8 + 5]) ||
                 (R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && B[4*8 + 6]) ||
                 (R[4*8 + 2] && R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && R[4*8 + 6] && B[4*8 + 7]) 
                 );
    M[4][1][UP45M] = (!R[4*8 + 1] && !B[4*8 + 1]) && 

                 (
                 (R[5*8 + 1] && B[6*8 + 1]) ||
                 (R[5*8 + 1] && R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[4][1][UP] = (!R[4*8 + 1] && !B[4*8 + 1]) && 

                 (
                 (R[3*8 + 1] && B[2*8 + 1]) ||
                 (R[3*8 + 1] && R[2*8 + 1] && B[1*8 + 1]) ||
                 (R[3*8 + 1] && R[2*8 + 1] && R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[4][1][UP45P] = 1'b0;
    M[3][1][ZEROP] = (!R[3*8 + 1] && !B[3*8 + 1]) && 

                 (
                 (R[4*8 + 2] && B[5*8 + 3]) ||
                 (R[4*8 + 2] && R[5*8 + 3] && B[6*8 + 4]) ||
                 (R[4*8 + 2] && R[5*8 + 3] && R[6*8 + 4] && B[7*8 + 5]) 
                 );
    M[3][1][DOWN45P] = 1'b0;
    M[3][1][DOWN] = 1'b0;
    M[3][1][DOWN45M] = (!R[3*8 + 1] && !B[3*8 + 1]) && 

                 (
                 (R[2*8 + 2] && B[1*8 + 3]) ||
                 (R[2*8 + 2] && R[1*8 + 3] && B[0*8 + 4]) 
                 );
    M[3][1][ZEROM] = (!R[3*8 + 1] && !B[3*8 + 1]) && 

                 (
                 (R[3*8 + 2] && B[3*8 + 3]) ||
                 (R[3*8 + 2] && R[3*8 + 3] && B[3*8 + 4]) ||
                 (R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && B[3*8 + 5]) ||
                 (R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && B[3*8 + 6]) ||
                 (R[3*8 + 2] && R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && R[3*8 + 6] && B[3*8 + 7]) 
                 );
    M[3][1][UP45M] = (!R[3*8 + 1] && !B[3*8 + 1]) && 

                 (
                 (R[4*8 + 1] && B[5*8 + 1]) ||
                 (R[4*8 + 1] && R[5*8 + 1] && B[6*8 + 1]) ||
                 (R[4*8 + 1] && R[5*8 + 1] && R[6*8 + 1] && B[7*8 + 1]) 
                 );
    M[3][1][UP] = (!R[3*8 + 1] && !B[3*8 + 1]) && 

                 (
                 (R[2*8 + 1] && B[1*8 + 1]) ||
                 (R[2*8 + 1] && R[1*8 + 1] && B[0*8 + 1]) 
                 );
    M[3][1][UP45P] = 1'b0;


// Expresii generate pentru patrate H
    M[2][2][ZEROP] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[3*8 + 3] && B[4*8 + 4]) ||
                 (R[3*8 + 3] && R[4*8 + 4] && B[5*8 + 5]) ||
                 (R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && B[6*8 + 6]) ||
                 (R[3*8 + 3] && R[4*8 + 4] && R[5*8 + 5] && R[6*8 + 6] && B[7*8 + 7]) 
                 );
    M[2][2][DOWN45P] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[3*8 + 1] && B[4*8 + 0]) 
                 );
    M[2][2][DOWN] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[1*8 + 1] && B[0*8 + 0]) 
                 );
    M[2][2][DOWN45M] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[1*8 + 3] && B[0*8 + 4]) 
                 );
    M[2][2][ZEROM] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[2*8 + 3] && B[2*8 + 4]) ||
                 (R[2*8 + 3] && R[2*8 + 4] && B[2*8 + 5]) ||
                 (R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && B[2*8 + 6]) ||
                 (R[2*8 + 3] && R[2*8 + 4] && R[2*8 + 5] && R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][2][UP45M] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[3*8 + 2] && B[4*8 + 2]) ||
                 (R[3*8 + 2] && R[4*8 + 2] && B[5*8 + 2]) ||
                 (R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && B[6*8 + 2]) ||
                 (R[3*8 + 2] && R[4*8 + 2] && R[5*8 + 2] && R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[2][2][UP] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[2][2][UP45P] = (!R[2*8 + 2] && !B[2*8 + 2]) && 

                 (
                 (R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[2][5][ZEROP] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[3*8 + 6] && B[4*8 + 7]) 
                 );
    M[2][5][DOWN45P] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[3*8 + 4] && B[4*8 + 3]) ||
                 (R[3*8 + 4] && R[4*8 + 3] && B[5*8 + 2]) ||
                 (R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && B[6*8 + 1]) ||
                 (R[3*8 + 4] && R[4*8 + 3] && R[5*8 + 2] && R[6*8 + 1] && B[7*8 + 0]) 
                 );
    M[2][5][DOWN] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[1*8 + 4] && B[0*8 + 3]) 
                 );
    M[2][5][DOWN45M] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[1*8 + 6] && B[0*8 + 7]) 
                 );
    M[2][5][ZEROM] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][5][UP45M] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[3*8 + 5] && B[4*8 + 5]) ||
                 (R[3*8 + 5] && R[4*8 + 5] && B[5*8 + 5]) ||
                 (R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && B[6*8 + 5]) ||
                 (R[3*8 + 5] && R[4*8 + 5] && R[5*8 + 5] && R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[2][5][UP] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[2][5][UP45P] = (!R[2*8 + 5] && !B[2*8 + 5]) && 

                 (
                 (R[2*8 + 4] && B[2*8 + 3]) ||
                 (R[2*8 + 4] && R[2*8 + 3] && B[2*8 + 2]) ||
                 (R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && B[2*8 + 1]) ||
                 (R[2*8 + 4] && R[2*8 + 3] && R[2*8 + 2] && R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[5][5][ZEROP] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[6*8 + 6] && B[7*8 + 7]) 
                 );
    M[5][5][DOWN45P] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[6*8 + 4] && B[7*8 + 3]) 
                 );
    M[5][5][DOWN] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[4*8 + 4] && B[3*8 + 3]) ||
                 (R[4*8 + 4] && R[3*8 + 3] && B[2*8 + 2]) ||
                 (R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && B[1*8 + 1]) ||
                 (R[4*8 + 4] && R[3*8 + 3] && R[2*8 + 2] && R[1*8 + 1] && B[0*8 + 0]) 
                 );
    M[5][5][DOWN45M] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[4*8 + 6] && B[3*8 + 7]) 
                 );
    M[5][5][ZEROM] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][5][UP45M] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[5][5][UP] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[4*8 + 5] && B[3*8 + 5]) ||
                 (R[4*8 + 5] && R[3*8 + 5] && B[2*8 + 5]) ||
                 (R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && B[1*8 + 5]) ||
                 (R[4*8 + 5] && R[3*8 + 5] && R[2*8 + 5] && R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[5][5][UP45P] = (!R[5*8 + 5] && !B[5*8 + 5]) && 

                 (
                 (R[5*8 + 4] && B[5*8 + 3]) ||
                 (R[5*8 + 4] && R[5*8 + 3] && B[5*8 + 2]) ||
                 (R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && B[5*8 + 1]) ||
                 (R[5*8 + 4] && R[5*8 + 3] && R[5*8 + 2] && R[5*8 + 1] && B[5*8 + 0]) 
                 );
    M[5][2][ZEROP] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[6*8 + 3] && B[7*8 + 4]) 
                 );
    M[5][2][DOWN45P] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[6*8 + 1] && B[7*8 + 0]) 
                 );
    M[5][2][DOWN] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[4*8 + 1] && B[3*8 + 0]) 
                 );
    M[5][2][DOWN45M] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[4*8 + 3] && B[3*8 + 4]) ||
                 (R[4*8 + 3] && R[3*8 + 4] && B[2*8 + 5]) ||
                 (R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && B[1*8 + 6]) ||
                 (R[4*8 + 3] && R[3*8 + 4] && R[2*8 + 5] && R[1*8 + 6] && B[0*8 + 7]) 
                 );
    M[5][2][ZEROM] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[5*8 + 3] && B[5*8 + 4]) ||
                 (R[5*8 + 3] && R[5*8 + 4] && B[5*8 + 5]) ||
                 (R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && B[5*8 + 6]) ||
                 (R[5*8 + 3] && R[5*8 + 4] && R[5*8 + 5] && R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][2][UP45M] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[5][2][UP] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[4*8 + 2] && B[3*8 + 2]) ||
                 (R[4*8 + 2] && R[3*8 + 2] && B[2*8 + 2]) ||
                 (R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && B[1*8 + 2]) ||
                 (R[4*8 + 2] && R[3*8 + 2] && R[2*8 + 2] && R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[5][2][UP45P] = (!R[5*8 + 2] && !B[5*8 + 2]) && 

                 (
                 (R[5*8 + 1] && B[5*8 + 0]) 
                 );


// Expresii generate pentru patrate I
    M[2][3][ZEROP] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[3*8 + 4] && B[4*8 + 5]) ||
                 (R[3*8 + 4] && R[4*8 + 5] && B[5*8 + 6]) ||
                 (R[3*8 + 4] && R[4*8 + 5] && R[5*8 + 6] && B[6*8 + 7]) 
                 );
    M[2][3][DOWN45P] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[3*8 + 2] && B[4*8 + 1]) ||
                 (R[3*8 + 2] && R[4*8 + 1] && B[5*8 + 0]) 
                 );
    M[2][3][DOWN] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[1*8 + 2] && B[0*8 + 1]) 
                 );
    M[2][3][DOWN45M] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[1*8 + 4] && B[0*8 + 5]) 
                 );
    M[2][3][ZEROM] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[2*8 + 4] && B[2*8 + 5]) ||
                 (R[2*8 + 4] && R[2*8 + 5] && B[2*8 + 6]) ||
                 (R[2*8 + 4] && R[2*8 + 5] && R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][3][UP45M] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[3*8 + 3] && B[4*8 + 3]) ||
                 (R[3*8 + 3] && R[4*8 + 3] && B[5*8 + 3]) ||
                 (R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && B[6*8 + 3]) ||
                 (R[3*8 + 3] && R[4*8 + 3] && R[5*8 + 3] && R[6*8 + 3] && B[7*8 + 3]) 
                 );
    M[2][3][UP] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[1*8 + 3] && B[0*8 + 3]) 
                 );
    M[2][3][UP45P] = (!R[2*8 + 3] && !B[2*8 + 3]) && 

                 (
                 (R[2*8 + 2] && B[2*8 + 1]) ||
                 (R[2*8 + 2] && R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[2][4][ZEROP] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[3*8 + 5] && B[4*8 + 6]) ||
                 (R[3*8 + 5] && R[4*8 + 6] && B[5*8 + 7]) 
                 );
    M[2][4][DOWN45P] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[3*8 + 3] && B[4*8 + 2]) ||
                 (R[3*8 + 3] && R[4*8 + 2] && B[5*8 + 1]) ||
                 (R[3*8 + 3] && R[4*8 + 2] && R[5*8 + 1] && B[6*8 + 0]) 
                 );
    M[2][4][DOWN] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[1*8 + 3] && B[0*8 + 2]) 
                 );
    M[2][4][DOWN45M] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[1*8 + 5] && B[0*8 + 6]) 
                 );
    M[2][4][ZEROM] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[2*8 + 5] && B[2*8 + 6]) ||
                 (R[2*8 + 5] && R[2*8 + 6] && B[2*8 + 7]) 
                 );
    M[2][4][UP45M] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[3*8 + 4] && B[4*8 + 4]) ||
                 (R[3*8 + 4] && R[4*8 + 4] && B[5*8 + 4]) ||
                 (R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && B[6*8 + 4]) ||
                 (R[3*8 + 4] && R[4*8 + 4] && R[5*8 + 4] && R[6*8 + 4] && B[7*8 + 4]) 
                 );
    M[2][4][UP] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[1*8 + 4] && B[0*8 + 4]) 
                 );
    M[2][4][UP45P] = (!R[2*8 + 4] && !B[2*8 + 4]) && 

                 (
                 (R[2*8 + 3] && B[2*8 + 2]) ||
                 (R[2*8 + 3] && R[2*8 + 2] && B[2*8 + 1]) ||
                 (R[2*8 + 3] && R[2*8 + 2] && R[2*8 + 1] && B[2*8 + 0]) 
                 );
    M[3][5][ZEROP] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[4*8 + 6] && B[5*8 + 7]) 
                 );
    M[3][5][DOWN45P] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[4*8 + 4] && B[5*8 + 3]) ||
                 (R[4*8 + 4] && R[5*8 + 3] && B[6*8 + 2]) ||
                 (R[4*8 + 4] && R[5*8 + 3] && R[6*8 + 2] && B[7*8 + 1]) 
                 );
    M[3][5][DOWN] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[2*8 + 4] && B[1*8 + 3]) ||
                 (R[2*8 + 4] && R[1*8 + 3] && B[0*8 + 2]) 
                 );
    M[3][5][DOWN45M] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[2*8 + 6] && B[1*8 + 7]) 
                 );
    M[3][5][ZEROM] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[3*8 + 6] && B[3*8 + 7]) 
                 );
    M[3][5][UP45M] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[4*8 + 5] && B[5*8 + 5]) ||
                 (R[4*8 + 5] && R[5*8 + 5] && B[6*8 + 5]) ||
                 (R[4*8 + 5] && R[5*8 + 5] && R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[3][5][UP] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[2*8 + 5] && B[1*8 + 5]) ||
                 (R[2*8 + 5] && R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[3][5][UP45P] = (!R[3*8 + 5] && !B[3*8 + 5]) && 

                 (
                 (R[3*8 + 4] && B[3*8 + 3]) ||
                 (R[3*8 + 4] && R[3*8 + 3] && B[3*8 + 2]) ||
                 (R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && B[3*8 + 1]) ||
                 (R[3*8 + 4] && R[3*8 + 3] && R[3*8 + 2] && R[3*8 + 1] && B[3*8 + 0]) 
                 );
    M[4][5][ZEROP] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[5*8 + 6] && B[6*8 + 7]) 
                 );
    M[4][5][DOWN45P] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[5*8 + 4] && B[6*8 + 3]) ||
                 (R[5*8 + 4] && R[6*8 + 3] && B[7*8 + 2]) 
                 );
    M[4][5][DOWN] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[3*8 + 4] && B[2*8 + 3]) ||
                 (R[3*8 + 4] && R[2*8 + 3] && B[1*8 + 2]) ||
                 (R[3*8 + 4] && R[2*8 + 3] && R[1*8 + 2] && B[0*8 + 1]) 
                 );
    M[4][5][DOWN45M] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[3*8 + 6] && B[2*8 + 7]) 
                 );
    M[4][5][ZEROM] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[4*8 + 6] && B[4*8 + 7]) 
                 );
    M[4][5][UP45M] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[5*8 + 5] && B[6*8 + 5]) ||
                 (R[5*8 + 5] && R[6*8 + 5] && B[7*8 + 5]) 
                 );
    M[4][5][UP] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[3*8 + 5] && B[2*8 + 5]) ||
                 (R[3*8 + 5] && R[2*8 + 5] && B[1*8 + 5]) ||
                 (R[3*8 + 5] && R[2*8 + 5] && R[1*8 + 5] && B[0*8 + 5]) 
                 );
    M[4][5][UP45P] = (!R[4*8 + 5] && !B[4*8 + 5]) && 

                 (
                 (R[4*8 + 4] && B[4*8 + 3]) ||
                 (R[4*8 + 4] && R[4*8 + 3] && B[4*8 + 2]) ||
                 (R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && B[4*8 + 1]) ||
                 (R[4*8 + 4] && R[4*8 + 3] && R[4*8 + 2] && R[4*8 + 1] && B[4*8 + 0]) 
                 );
    M[5][4][ZEROP] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[6*8 + 5] && B[7*8 + 6]) 
                 );
    M[5][4][DOWN45P] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[6*8 + 3] && B[7*8 + 2]) 
                 );
    M[5][4][DOWN] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[4*8 + 3] && B[3*8 + 2]) ||
                 (R[4*8 + 3] && R[3*8 + 2] && B[2*8 + 1]) ||
                 (R[4*8 + 3] && R[3*8 + 2] && R[2*8 + 1] && B[1*8 + 0]) 
                 );
    M[5][4][DOWN45M] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[4*8 + 5] && B[3*8 + 6]) ||
                 (R[4*8 + 5] && R[3*8 + 6] && B[2*8 + 7]) 
                 );
    M[5][4][ZEROM] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[5*8 + 5] && B[5*8 + 6]) ||
                 (R[5*8 + 5] && R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][4][UP45M] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[6*8 + 4] && B[7*8 + 4]) 
                 );
    M[5][4][UP] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[4*8 + 4] && B[3*8 + 4]) ||
                 (R[4*8 + 4] && R[3*8 + 4] && B[2*8 + 4]) ||
                 (R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && B[1*8 + 4]) ||
                 (R[4*8 + 4] && R[3*8 + 4] && R[2*8 + 4] && R[1*8 + 4] && B[0*8 + 4]) 
                 );
    M[5][4][UP45P] = (!R[5*8 + 4] && !B[5*8 + 4]) && 

                 (
                 (R[5*8 + 3] && B[5*8 + 2]) ||
                 (R[5*8 + 3] && R[5*8 + 2] && B[5*8 + 1]) ||
                 (R[5*8 + 3] && R[5*8 + 2] && R[5*8 + 1] && B[5*8 + 0]) 
                 );
    M[5][3][ZEROP] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[6*8 + 4] && B[7*8 + 5]) 
                 );
    M[5][3][DOWN45P] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[6*8 + 2] && B[7*8 + 1]) 
                 );
    M[5][3][DOWN] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[4*8 + 2] && B[3*8 + 1]) ||
                 (R[4*8 + 2] && R[3*8 + 1] && B[2*8 + 0]) 
                 );
    M[5][3][DOWN45M] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[4*8 + 4] && B[3*8 + 5]) ||
                 (R[4*8 + 4] && R[3*8 + 5] && B[2*8 + 6]) ||
                 (R[4*8 + 4] && R[3*8 + 5] && R[2*8 + 6] && B[1*8 + 7]) 
                 );
    M[5][3][ZEROM] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[5*8 + 4] && B[5*8 + 5]) ||
                 (R[5*8 + 4] && R[5*8 + 5] && B[5*8 + 6]) ||
                 (R[5*8 + 4] && R[5*8 + 5] && R[5*8 + 6] && B[5*8 + 7]) 
                 );
    M[5][3][UP45M] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[6*8 + 3] && B[7*8 + 3]) 
                 );
    M[5][3][UP] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[4*8 + 3] && B[3*8 + 3]) ||
                 (R[4*8 + 3] && R[3*8 + 3] && B[2*8 + 3]) ||
                 (R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && B[1*8 + 3]) ||
                 (R[4*8 + 3] && R[3*8 + 3] && R[2*8 + 3] && R[1*8 + 3] && B[0*8 + 3]) 
                 );
    M[5][3][UP45P] = (!R[5*8 + 3] && !B[5*8 + 3]) && 

                 (
                 (R[5*8 + 2] && B[5*8 + 1]) ||
                 (R[5*8 + 2] && R[5*8 + 1] && B[5*8 + 0]) 
                 );
    M[4][2][ZEROP] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[5*8 + 3] && B[6*8 + 4]) ||
                 (R[5*8 + 3] && R[6*8 + 4] && B[7*8 + 5]) 
                 );
    M[4][2][DOWN45P] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[5*8 + 1] && B[6*8 + 0]) 
                 );
    M[4][2][DOWN] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[3*8 + 1] && B[2*8 + 0]) 
                 );
    M[4][2][DOWN45M] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[3*8 + 3] && B[2*8 + 4]) ||
                 (R[3*8 + 3] && R[2*8 + 4] && B[1*8 + 5]) ||
                 (R[3*8 + 3] && R[2*8 + 4] && R[1*8 + 5] && B[0*8 + 6]) 
                 );
    M[4][2][ZEROM] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[4*8 + 3] && B[4*8 + 4]) ||
                 (R[4*8 + 3] && R[4*8 + 4] && B[4*8 + 5]) ||
                 (R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && B[4*8 + 6]) ||
                 (R[4*8 + 3] && R[4*8 + 4] && R[4*8 + 5] && R[4*8 + 6] && B[4*8 + 7]) 
                 );
    M[4][2][UP45M] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[5*8 + 2] && B[6*8 + 2]) ||
                 (R[5*8 + 2] && R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[4][2][UP] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[3*8 + 2] && B[2*8 + 2]) ||
                 (R[3*8 + 2] && R[2*8 + 2] && B[1*8 + 2]) ||
                 (R[3*8 + 2] && R[2*8 + 2] && R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[4][2][UP45P] = (!R[4*8 + 2] && !B[4*8 + 2]) && 

                 (
                 (R[4*8 + 1] && B[4*8 + 0]) 
                 );
    M[3][2][ZEROP] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[4*8 + 3] && B[5*8 + 4]) ||
                 (R[4*8 + 3] && R[5*8 + 4] && B[6*8 + 5]) ||
                 (R[4*8 + 3] && R[5*8 + 4] && R[6*8 + 5] && B[7*8 + 6]) 
                 );
    M[3][2][DOWN45P] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[4*8 + 1] && B[5*8 + 0]) 
                 );
    M[3][2][DOWN] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[2*8 + 1] && B[1*8 + 0]) 
                 );
    M[3][2][DOWN45M] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[2*8 + 3] && B[1*8 + 4]) ||
                 (R[2*8 + 3] && R[1*8 + 4] && B[0*8 + 5]) 
                 );
    M[3][2][ZEROM] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[3*8 + 3] && B[3*8 + 4]) ||
                 (R[3*8 + 3] && R[3*8 + 4] && B[3*8 + 5]) ||
                 (R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && B[3*8 + 6]) ||
                 (R[3*8 + 3] && R[3*8 + 4] && R[3*8 + 5] && R[3*8 + 6] && B[3*8 + 7]) 
                 );
    M[3][2][UP45M] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[4*8 + 2] && B[5*8 + 2]) ||
                 (R[4*8 + 2] && R[5*8 + 2] && B[6*8 + 2]) ||
                 (R[4*8 + 2] && R[5*8 + 2] && R[6*8 + 2] && B[7*8 + 2]) 
                 );
    M[3][2][UP] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[2*8 + 2] && B[1*8 + 2]) ||
                 (R[2*8 + 2] && R[1*8 + 2] && B[0*8 + 2]) 
                 );
    M[3][2][UP45P] = (!R[3*8 + 2] && !B[3*8 + 2]) && 

                 (
                 (R[3*8 + 1] && B[3*8 + 0]) 
                 );
    M[3][3][7:0] = 8'b00000000;
    M[3][4][7:0] = 8'b00000000;
    M[4][3][7:0] = 8'b00000000;
    M[4][4][7:0] = 8'b00000000;
	 
	RES_D[1*7 + 0 : 0*7 + 0] = {|M[0][7], |M[0][6], |M[0][5], |M[0][4], |M[0][3], |M[0][2], |M[0][1], |M[0][0]};
	RES_D[2*7 + 1 : 1*7 + 1] = {|M[1][7], |M[1][6], |M[1][5], |M[1][4], |M[1][3], |M[1][2], |M[1][1], |M[1][0]};
	RES_D[3*7 + 2 : 2*7 + 2] = {|M[2][7], |M[2][6], |M[2][5], |M[2][4], |M[2][3], |M[2][2], |M[2][1], |M[2][0]};
	RES_D[4*7 + 3 : 3*7 + 3] = {|M[3][7], |M[3][6], |M[3][5], |M[3][4], |M[3][3], |M[3][2], |M[3][1], |M[3][0]};
	RES_D[5*7 + 4 : 4*7 + 4] = {|M[4][7], |M[4][6], |M[4][5], |M[4][4], |M[4][3], |M[4][2], |M[4][1], |M[4][0]};
	RES_D[6*7 + 5 : 5*7 + 5] = {|M[5][7], |M[5][6], |M[5][5], |M[5][4], |M[5][3], |M[5][2], |M[5][1], |M[5][0]};
	RES_D[7*7 + 6 : 6*7 + 6] = {|M[6][7], |M[6][6], |M[6][5], |M[6][4], |M[6][3], |M[6][2], |M[6][1], |M[6][0]};
	RES_D[8*7 + 7 : 7*7 + 7] = {|M[7][7], |M[7][6], |M[7][5], |M[7][4], |M[7][3], |M[7][2], |M[7][1], |M[7][0]};	
  end
       
assign M_ = RES_Q;

endmodule
