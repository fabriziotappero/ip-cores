-- GRCAN 2.0 interface
  constant CFG_GRCAN      : integer := CONFIG_GRCAN_ENABLE;
  constant CFG_GRCAN_NUM  : integer := CONFIG_GRCAN_NUM;
  constant CFG_GRCANSEP   : integer := CONFIG_GRCANSEP;
  constant CFG_GRCANIRQ   : integer := CONFIG_GRCANIRQ;

