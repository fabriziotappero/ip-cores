-------------------------------------------------------------------------------------------------100
--| Modular Oscilloscope
--| UNSL - Argentine
--|
--| File: dual_port_memory_wb.vhd
--| Version: 0.1
--| Tested in: Actel A3PE1500
--|-------------------------------------------------------------------------------------------------
--| Description:
--|   MEMORY - Dual Port Memory Wishbone Interface
--|   An interface designed for a dual port memory generated by Actel SmartGen tool. It may not work 
--|   with other than ProASIC3 Family FPGA.
--|   
--|-------------------------------------------------------------------------------------------------
--| File history:
--|   0.1   | jun-2009 | First testing
--|   0.11  | aug-2009 | Corrected error in ACK_O from port B
----------------------------------------------------------------------------------------------------
--| Copyright � 2009, Facundo Aguilera.
--|
--| This VHDL design file is an open design; you can redistribute it and/or
--| modify it and/or implement it after contacting the author.

--| Wishbone Rev. B.3 compatible
----------------------------------------------------------------------------------------------------

-- La memoria solo puede accederse desde la direcci�n 0 hasta la 15360 (0011 11000 0000 0000). No 
-- est�n especificados los valores obtenidos fuera de ese rango. 


library ieee;
use ieee.std_logic_1164.all;

entity dual_port_memory_wb is
	port(
		-- Puerto A (Higer prioriry)
		RST_I_a: in std_logic;  
		CLK_I_a: in std_logic;  
		DAT_I_a: in std_logic_vector (15 downto 0);
		DAT_O_a: out std_logic_vector (15 downto 0);
		ADR_I_a: in std_logic_vector (13 downto 0);
		CYC_I_a: in std_logic;  
		STB_I_a: in std_logic;  
		ACK_O_a: out std_logic ;
		WE_I_a: in std_logic;
		
    
    -- Puerto B (Lower prioriry)
		RST_I_b: in std_logic;  
		CLK_I_b: in std_logic;  
		DAT_I_b: in std_logic_vector (15 downto 0);
		DAT_O_b: out std_logic_vector (15 downto 0);
		ADR_I_b: in std_logic_vector (13 downto 0);
		CYC_I_b: in std_logic;  
		STB_I_b: in std_logic;  
		ACK_O_b: out std_logic ;
		WE_I_b: in std_logic
	);
end entity dual_port_memory_wb;



architecture arch01  of dual_port_memory_wb is 
	---- Componentes ----
  component dual_port_memory is 
    port( 
      DINA:   in    std_logic_vector(15 downto 0); 
      DOUTA:  out   std_logic_vector(15 downto 0);  
      ADDRA:  in    std_logic_vector(13 downto 0);  -- Only available up to 15360 (11110000000000)
      RWA:    in    std_logic;                      -- '1' Read, '0' Write
      BLKA:   in    std_logic;                      -- '1' Block select
      CLKA:   in    std_logic;                      -- Rising edge

      DINB:   in    std_logic_vector(15 downto 0); 
      DOUTB:  out   std_logic_vector(15 downto 0); 
      ADDRB:  in    std_logic_vector(13 downto 0);
      RWB:    in    std_logic; 
      BLKB:   in    std_logic; 
      CLKB:   in    std_logic;

      RESET:  in    std_logic                       -- '1' Reset
    ) ;
        
	end component dual_port_memory;
	
  ---- Se�ales ----
	signal RST_I_common: std_logic;
  signal enable_BLK, to_BLKB, to_BLKA : std_logic;
  signal pre_ACK_O_a_read, pre_ACK_O_a_write: std_logic;
  signal pre_ACK_O_b_read, pre_ACK_O_b_write: std_logic;
  signal to_RWB, to_RWA: std_logic; -- para entradas negadas

	
begin	

  RST_I_common <= RST_I_b or RST_I_a;

  
  -- Correcci�n de escritura en la misma direcci�n
  to_BLKB <= CYC_I_b and STB_I_b and enable_BLK;
  to_BLKA <= CYC_I_a and STB_I_a;
   
  enable_BLK <= '1' when ADR_I_a /= ADR_I_b or to_BLKA = '0' else
                '0';
  
  
  -- Soluci�n de ACK en puerto A
  ACK_O_a <= pre_ACK_O_a_write or pre_ACK_O_a_read;
  pre_ACK_O_a_write <= STB_I_a and CYC_I_a and WE_I_a;
    -- la primera respuesta para el ciclo de lectura debe retrasarse un ciclo
  P_ACK_a_resolution: process (STB_I_a, CYC_I_a, RST_I_a, CLK_I_a, WE_I_a)
  begin
    if STB_I_a = '0' or CYC_I_a = '0' then
      pre_ACK_O_a_read <= '0';      
    elsif CLK_I_a'event and CLK_I_a = '1' then
      if RST_I_a = '1' then
        pre_ACK_O_a_read <= '0';
      elsif STB_I_a = '1' and CYC_I_a = '1' and WE_I_a = '0' then
        pre_ACK_O_a_read <= '1';
      end if;
    end if;
  end process;
  
   -- Soluci�n de ACK en puerto B
  ACK_O_b <= (pre_ACK_O_b_write or pre_ACK_O_b_read) and enable_BLK;
  pre_ACK_O_b_write <= STB_I_b and CYC_I_b and WE_I_b;
    -- la primera respuesta para el ciclo de lectura debe retrasarse un ciclo
  P_ACK_b_resolution: process (STB_I_b, CYC_I_b, RST_I_b, CLK_I_b)
  begin
    if STB_I_b = '0' or CYC_I_b = '0' then
      pre_ACK_O_b_read <= '0';      
    elsif CLK_I_b'event and CLK_I_b = '1' then
      if RST_I_b = '1' then
        pre_ACK_O_b_read <= '0';
      elsif STB_I_b = '1' and CYC_I_b = '1' and WE_I_b = '0'  then
        pre_ACK_O_b_read <= '1';
      end if;
    end if;
  end process;
  
  
  -- Instancia
  to_RWA <= not(WE_I_a);
  to_RWB <= not(WE_I_b);
	MEM: dual_port_memory port map (
			DINA => DAT_I_a,
			DOUTA => DAT_O_a,
			ADDRA => ADR_I_a,
			RWA => to_RWA,
			BLKA => to_BLKA,
			CLKA => CLK_I_a,

			DINB => DAT_I_b,
			DOUTB => DAT_O_b,
			ADDRB => ADR_I_b,
			RWB => to_RWB,
			BLKB => to_BLKB,
			CLKB => CLK_I_b,

			RESET => RST_I_common
	);
  

end architecture;
