-- ADCDAC enable 
  constant CFG_ADCDAC  : integer := CONFIG_ADCDAC_ENABLE;

