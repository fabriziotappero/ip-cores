/*
 Asynchronous SDM NoC
 (C)2011 Wei Song
 Advanced Processor Technologies Group
 Computer Science, the Univ. of Manchester, UK
 
 Authors: 
 Wei Song     wsong83@gmail.com
 
 License: LGPL 3.0 or later
 
 The SystemC to keep a module of the simulation analysis object. 
 
 History:
 27/02/2011  Initial version. <wsong83@gmail.com>
 30/05/2011  Clean up for opensource. <wsong83@gmail.com>
 
*/

module AnaProc ()
   //
   // The foreign attribute string value must be a SystemC value.
   //
   (* integer foreign = "SystemC";
    *);
   //
   // Verilog port names must match port names exactly as they appear in the
   // sc_module class in SystemC; they must also match in order, mode, and type.
   //
   
endmodule
   