-- GRLIB debugging
  constant CFG_DUART    : integer := CONFIG_DEBUG_UART;

