-------------------------------------------------------------------------------
--
-- A testbench model for the
-- GCpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: gcpad_mod-c.vhd 41 2009-04-01 19:58:04Z arniml $
--
-------------------------------------------------------------------------------

configuration gcpad_mod_behav_c0 of gcpad_mod is

  for behav
  end for;

end gcpad_mod_behav_c0;
