
--------------------------------------------------------------------------------
-- Designer:      Paolo Fulgoni <pfulgoni@opencores.org>
--
-- Create Date:   01/22/2008
-- Last Update:   01/22/2008
-- Project Name:  camellia-vhdl
-- Description:   Asynchronous SBOX1
--
-- Copyright (C) 2008  Paolo Fulgoni
-- This file is part of camellia-vhdl.
-- camellia-vhdl is free software; you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation; either version 3 of the License, or
-- (at your option) any later version.
-- camellia-vhdl is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
-- The Camellia cipher algorithm is 128 bit cipher developed by NTT and
-- Mitsubishi Electric researchers.
-- http://info.isl.ntt.co.jp/crypt/eng/camellia/
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;


entity SBOX1 is
    port  (
            data_in  : IN STD_LOGIC_VECTOR(0 to 7);
            data_out : OUT STD_LOGIC_VECTOR(0 to 7)
            );
end SBOX1;

architecture RTL of SBOX1 is
begin

    with data_in select
        data_out <= X"70" when X"00",
                    X"82" when X"01",
                    X"2C" when X"02",
                    X"EC" when X"03",
                    X"B3" when X"04",
                    X"27" when X"05",
                    X"C0" when X"06",
                    X"E5" when X"07",
                    X"E4" when X"08",
                    X"85" when X"09",
                    X"57" when X"0A",
                    X"35" when X"0B",
                    X"EA" when X"0C",
                    X"0C" when X"0D",
                    X"AE" when X"0E",
                    X"41" when X"0F",
                    X"23" when X"10",
                    X"EF" when X"11",
                    X"6B" when X"12",
                    X"93" when X"13",
                    X"45" when X"14",
                    X"19" when X"15",
                    X"A5" when X"16",
                    X"21" when X"17",
                    X"ED" when X"18",
                    X"0E" when X"19",
                    X"4F" when X"1A",
                    X"4E" when X"1B",
                    X"1D" when X"1C",
                    X"65" when X"1D",
                    X"92" when X"1E",
                    X"BD" when X"1F",
                    X"86" when X"20",
                    X"B8" when X"21",
                    X"AF" when X"22",
                    X"8F" when X"23",
                    X"7C" when X"24",
                    X"EB" when X"25",
                    X"1F" when X"26",
                    X"CE" when X"27",
                    X"3E" when X"28",
                    X"30" when X"29",
                    X"DC" when X"2A",
                    X"5F" when X"2B",
                    X"5E" when X"2C",
                    X"C5" when X"2D",
                    X"0B" when X"2E",
                    X"1A" when X"2F",
                    X"A6" when X"30",
                    X"E1" when X"31",
                    X"39" when X"32",
                    X"CA" when X"33",
                    X"D5" when X"34",
                    X"47" when X"35",
                    X"5D" when X"36",
                    X"3D" when X"37",
                    X"D9" when X"38",
                    X"01" when X"39",
                    X"5A" when X"3A",
                    X"D6" when X"3B",
                    X"51" when X"3C",
                    X"56" when X"3D",
                    X"6C" when X"3E",
                    X"4D" when X"3F",
                    X"8B" when X"40",
                    X"0D" when X"41",
                    X"9A" when X"42",
                    X"66" when X"43",
                    X"FB" when X"44",
                    X"CC" when X"45",
                    X"B0" when X"46",
                    X"2D" when X"47",
                    X"74" when X"48",
                    X"12" when X"49",
                    X"2B" when X"4A",
                    X"20" when X"4B",
                    X"F0" when X"4C",
                    X"B1" when X"4D",
                    X"84" when X"4E",
                    X"99" when X"4F",
                    X"DF" when X"50",
                    X"4C" when X"51",
                    X"CB" when X"52",
                    X"C2" when X"53",
                    X"34" when X"54",
                    X"7E" when X"55",
                    X"76" when X"56",
                    X"05" when X"57",
                    X"6D" when X"58",
                    X"B7" when X"59",
                    X"A9" when X"5A",
                    X"31" when X"5B",
                    X"D1" when X"5C",
                    X"17" when X"5D",
                    X"04" when X"5E",
                    X"D7" when X"5F",
                    X"14" when X"60",
                    X"58" when X"61",
                    X"3A" when X"62",
                    X"61" when X"63",
                    X"DE" when X"64",
                    X"1B" when X"65",
                    X"11" when X"66",
                    X"1C" when X"67",
                    X"32" when X"68",
                    X"0F" when X"69",
                    X"9C" when X"6A",
                    X"16" when X"6B",
                    X"53" when X"6C",
                    X"18" when X"6D",
                    X"F2" when X"6E",
                    X"22" when X"6F",
                    X"FE" when X"70",
                    X"44" when X"71",
                    X"CF" when X"72",
                    X"B2" when X"73",
                    X"C3" when X"74",
                    X"B5" when X"75",
                    X"7A" when X"76",
                    X"91" when X"77",
                    X"24" when X"78",
                    X"08" when X"79",
                    X"E8" when X"7A",
                    X"A8" when X"7B",
                    X"60" when X"7C",
                    X"FC" when X"7D",
                    X"69" when X"7E",
                    X"50" when X"7F",
                    X"AA" when X"80",
                    X"D0" when X"81",
                    X"A0" when X"82",
                    X"7D" when X"83",
                    X"A1" when X"84",
                    X"89" when X"85",
                    X"62" when X"86",
                    X"97" when X"87",
                    X"54" when X"88",
                    X"5B" when X"89",
                    X"1E" when X"8A",
                    X"95" when X"8B",
                    X"E0" when X"8C",
                    X"FF" when X"8D",
                    X"64" when X"8E",
                    X"D2" when X"8F",
                    X"10" when X"90",
                    X"C4" when X"91",
                    X"00" when X"92",
                    X"48" when X"93",
                    X"A3" when X"94",
                    X"F7" when X"95",
                    X"75" when X"96",
                    X"DB" when X"97",
                    X"8A" when X"98",
                    X"03" when X"99",
                    X"E6" when X"9A",
                    X"DA" when X"9B",
                    X"09" when X"9C",
                    X"3F" when X"9D",
                    X"DD" when X"9E",
                    X"94" when X"9F",
                    X"87" when X"A0",
                    X"5C" when X"A1",
                    X"83" when X"A2",
                    X"02" when X"A3",
                    X"CD" when X"A4",
                    X"4A" when X"A5",
                    X"90" when X"A6",
                    X"33" when X"A7",
                    X"73" when X"A8",
                    X"67" when X"A9",
                    X"F6" when X"AA",
                    X"F3" when X"AB",
                    X"9D" when X"AC",
                    X"7F" when X"AD",
                    X"BF" when X"AE",
                    X"E2" when X"AF",
                    X"52" when X"B0",
                    X"9B" when X"B1",
                    X"D8" when X"B2",
                    X"26" when X"B3",
                    X"C8" when X"B4",
                    X"37" when X"B5",
                    X"C6" when X"B6",
                    X"3B" when X"B7",
                    X"81" when X"B8",
                    X"96" when X"B9",
                    X"6F" when X"BA",
                    X"4B" when X"BB",
                    X"13" when X"BC",
                    X"BE" when X"BD",
                    X"63" when X"BE",
                    X"2E" when X"BF",
                    X"E9" when X"C0",
                    X"79" when X"C1",
                    X"A7" when X"C2",
                    X"8C" when X"C3",
                    X"9F" when X"C4",
                    X"6E" when X"C5",
                    X"BC" when X"C6",
                    X"8E" when X"C7",
                    X"29" when X"C8",
                    X"F5" when X"C9",
                    X"F9" when X"CA",
                    X"B6" when X"CB",
                    X"2F" when X"CC",
                    X"FD" when X"CD",
                    X"B4" when X"CE",
                    X"59" when X"CF",
                    X"78" when X"D0",
                    X"98" when X"D1",
                    X"06" when X"D2",
                    X"6A" when X"D3",
                    X"E7" when X"D4",
                    X"46" when X"D5",
                    X"71" when X"D6",
                    X"BA" when X"D7",
                    X"D4" when X"D8",
                    X"25" when X"D9",
                    X"AB" when X"DA",
                    X"42" when X"DB",
                    X"88" when X"DC",
                    X"A2" when X"DD",
                    X"8D" when X"DE",
                    X"FA" when X"DF",
                    X"72" when X"E0",
                    X"07" when X"E1",
                    X"B9" when X"E2",
                    X"55" when X"E3",
                    X"F8" when X"E4",
                    X"EE" when X"E5",
                    X"AC" when X"E6",
                    X"0A" when X"E7",
                    X"36" when X"E8",
                    X"49" when X"E9",
                    X"2A" when X"EA",
                    X"68" when X"EB",
                    X"3C" when X"EC",
                    X"38" when X"ED",
                    X"F1" when X"EE",
                    X"A4" when X"EF",
                    X"40" when X"F0",
                    X"28" when X"F1",
                    X"D3" when X"F2",
                    X"7B" when X"F3",
                    X"BB" when X"F4",
                    X"C9" when X"F5",
                    X"43" when X"F6",
                    X"C1" when X"F7",
                    X"15" when X"F8",
                    X"E3" when X"F9",
                    X"AD" when X"FA",
                    X"F4" when X"FB",
                    X"77" when X"FC",
                    X"C7" when X"FD",
                    X"80" when X"FE",
                    X"9E" when X"FF",
                    "--------" when others;

end RTL;
