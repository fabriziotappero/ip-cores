-- I2C master
  constant CFG_I2C_ENABLE : integer := CONFIG_I2C_ENABLE;

