-----------------------------------------------------------------
--                                                             --
-----------------------------------------------------------------
--                                                             --
-- Copyright (C) 2013 Stefano Tonello                          --
--                                                             --
-- This source file may be used and distributed without        --
-- restriction provided that this copyright statement is not   --
-- removed from the file and that any derivative work contains --
-- the original copyright notice and the associated disclaimer.--
--                                                             --
-- THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY         --
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   --
-- TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   --
-- FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      --
-- OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         --
-- INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    --
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   --
-- GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        --
-- BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  --
-- LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  --
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  --
-- OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         --
-- POSSIBILITY OF SUCH DAMAGE.                                 --
--                                                             --
-----------------------------------------------------------------

---------------------------------------------------------------
-- G.729a Codec Self-test ROMs package
---------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library WORK;
use work.G729A_ASIP_PKG.all;
use work.G729A_ASIP_CFG_PKG.all;

package G729A_CODEC_ST_ROM_PKG is

  subtype ROM_WORD_T is std_logic_vector(SDLEN-1 downto 0);

  type ROM_DATA_T is array (0 to 425-1) of ROM_WORD_T;

  constant STI_ROM_INIT_DATA : ROM_DATA_T := (
    to_std_logic_vector(to_signed(-5752,SDLEN)),
    to_std_logic_vector(to_signed(160,SDLEN)),
    to_std_logic_vector(to_signed(250,SDLEN)),
    to_std_logic_vector(to_signed(-15681,SDLEN)),
    to_std_logic_vector(to_signed(-18462,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(86,SDLEN)),
    to_std_logic_vector(to_signed(94,SDLEN)),
    to_std_logic_vector(to_signed(102,SDLEN)),
    to_std_logic_vector(to_signed(109,SDLEN)),
    to_std_logic_vector(to_signed(117,SDLEN)),
    to_std_logic_vector(to_signed(125,SDLEN)),
    to_std_logic_vector(to_signed(133,SDLEN)),
    to_std_logic_vector(to_signed(141,SDLEN)),
    to_std_logic_vector(to_signed(148,SDLEN)),
    to_std_logic_vector(to_signed(155,SDLEN)),
    to_std_logic_vector(to_signed(162,SDLEN)),
    to_std_logic_vector(to_signed(169,SDLEN)),
    to_std_logic_vector(to_signed(174,SDLEN)),
    to_std_logic_vector(to_signed(179,SDLEN)),
    to_std_logic_vector(to_signed(184,SDLEN)),
    to_std_logic_vector(to_signed(187,SDLEN)),
    to_std_logic_vector(to_signed(189,SDLEN)),
    to_std_logic_vector(to_signed(191,SDLEN)),
    to_std_logic_vector(to_signed(190,SDLEN)),
    to_std_logic_vector(to_signed(189,SDLEN)),
    to_std_logic_vector(to_signed(186,SDLEN)),
    to_std_logic_vector(to_signed(181,SDLEN)),
    to_std_logic_vector(to_signed(174,SDLEN)),
    to_std_logic_vector(to_signed(166,SDLEN)),
    to_std_logic_vector(to_signed(156,SDLEN)),
    to_std_logic_vector(to_signed(143,SDLEN)),
    to_std_logic_vector(to_signed(129,SDLEN)),
    to_std_logic_vector(to_signed(113,SDLEN)),
    to_std_logic_vector(to_signed(95,SDLEN)),
    to_std_logic_vector(to_signed(75,SDLEN)),
    to_std_logic_vector(to_signed(54,SDLEN)),
    to_std_logic_vector(to_signed(31,SDLEN)),
    to_std_logic_vector(to_signed(6,SDLEN)),
    to_std_logic_vector(to_signed(-19,SDLEN)),
    to_std_logic_vector(to_signed(-46,SDLEN)),
    to_std_logic_vector(to_signed(-74,SDLEN)),
    to_std_logic_vector(to_signed(-102,SDLEN)),
    to_std_logic_vector(to_signed(-131,SDLEN)),
    to_std_logic_vector(to_signed(-159,SDLEN)),
    to_std_logic_vector(to_signed(-186,SDLEN)),
    to_std_logic_vector(to_signed(-212,SDLEN)),
    to_std_logic_vector(to_signed(-236,SDLEN)),
    to_std_logic_vector(to_signed(-258,SDLEN)),
    to_std_logic_vector(to_signed(-277,SDLEN)),
    to_std_logic_vector(to_signed(-293,SDLEN)),
    to_std_logic_vector(to_signed(-306,SDLEN)),
    to_std_logic_vector(to_signed(-314,SDLEN)),
    to_std_logic_vector(to_signed(-318,SDLEN)),
    to_std_logic_vector(to_signed(-317,SDLEN)),
    to_std_logic_vector(to_signed(-311,SDLEN)),
    to_std_logic_vector(to_signed(-29314,SDLEN)),
    to_std_logic_vector(to_signed(6197,SDLEN)),
    to_std_logic_vector(to_signed(7439,SDLEN)),
    to_std_logic_vector(to_signed(-11681,SDLEN)),
    to_std_logic_vector(to_signed(22234,SDLEN)),
    to_std_logic_vector(to_signed(-300,SDLEN)),
    to_std_logic_vector(to_signed(-283,SDLEN)),
    to_std_logic_vector(to_signed(-260,SDLEN)),
    to_std_logic_vector(to_signed(-232,SDLEN)),
    to_std_logic_vector(to_signed(-199,SDLEN)),
    to_std_logic_vector(to_signed(-160,SDLEN)),
    to_std_logic_vector(to_signed(-118,SDLEN)),
    to_std_logic_vector(to_signed(-71,SDLEN)),
    to_std_logic_vector(to_signed(-22,SDLEN)),
    to_std_logic_vector(to_signed(28,SDLEN)),
    to_std_logic_vector(to_signed(81,SDLEN)),
    to_std_logic_vector(to_signed(134,SDLEN)),
    to_std_logic_vector(to_signed(185,SDLEN)),
    to_std_logic_vector(to_signed(235,SDLEN)),
    to_std_logic_vector(to_signed(280,SDLEN)),
    to_std_logic_vector(to_signed(320,SDLEN)),
    to_std_logic_vector(to_signed(355,SDLEN)),
    to_std_logic_vector(to_signed(382,SDLEN)),
    to_std_logic_vector(to_signed(400,SDLEN)),
    to_std_logic_vector(to_signed(409,SDLEN)),
    to_std_logic_vector(to_signed(408,SDLEN)),
    to_std_logic_vector(to_signed(396,SDLEN)),
    to_std_logic_vector(to_signed(374,SDLEN)),
    to_std_logic_vector(to_signed(341,SDLEN)),
    to_std_logic_vector(to_signed(298,SDLEN)),
    to_std_logic_vector(to_signed(245,SDLEN)),
    to_std_logic_vector(to_signed(183,SDLEN)),
    to_std_logic_vector(to_signed(115,SDLEN)),
    to_std_logic_vector(to_signed(41,SDLEN)),
    to_std_logic_vector(to_signed(-35,SDLEN)),
    to_std_logic_vector(to_signed(-113,SDLEN)),
    to_std_logic_vector(to_signed(-190,SDLEN)),
    to_std_logic_vector(to_signed(-262,SDLEN)),
    to_std_logic_vector(to_signed(-329,SDLEN)),
    to_std_logic_vector(to_signed(-386,SDLEN)),
    to_std_logic_vector(to_signed(-432,SDLEN)),
    to_std_logic_vector(to_signed(-465,SDLEN)),
    to_std_logic_vector(to_signed(-482,SDLEN)),
    to_std_logic_vector(to_signed(-483,SDLEN)),
    to_std_logic_vector(to_signed(-467,SDLEN)),
    to_std_logic_vector(to_signed(-434,SDLEN)),
    to_std_logic_vector(to_signed(-384,SDLEN)),
    to_std_logic_vector(to_signed(-318,SDLEN)),
    to_std_logic_vector(to_signed(-239,SDLEN)),
    to_std_logic_vector(to_signed(-148,SDLEN)),
    to_std_logic_vector(to_signed(-50,SDLEN)),
    to_std_logic_vector(to_signed(52,SDLEN)),
    to_std_logic_vector(to_signed(155,SDLEN)),
    to_std_logic_vector(to_signed(254,SDLEN)),
    to_std_logic_vector(to_signed(345,SDLEN)),
    to_std_logic_vector(to_signed(424,SDLEN)),
    to_std_logic_vector(to_signed(486,SDLEN)),
    to_std_logic_vector(to_signed(528,SDLEN)),
    to_std_logic_vector(to_signed(548,SDLEN)),
    to_std_logic_vector(to_signed(544,SDLEN)),
    to_std_logic_vector(to_signed(515,SDLEN)),
    to_std_logic_vector(to_signed(461,SDLEN)),
    to_std_logic_vector(to_signed(385,SDLEN)),
    to_std_logic_vector(to_signed(289,SDLEN)),
    to_std_logic_vector(to_signed(177,SDLEN)),
    to_std_logic_vector(to_signed(53,SDLEN)),
    to_std_logic_vector(to_signed(-74,SDLEN)),
    to_std_logic_vector(to_signed(-202,SDLEN)),
    to_std_logic_vector(to_signed(-322,SDLEN)),
    to_std_logic_vector(to_signed(-428,SDLEN)),
    to_std_logic_vector(to_signed(-513,SDLEN)),
    to_std_logic_vector(to_signed(-573,SDLEN)),
    to_std_logic_vector(to_signed(-604,SDLEN)),
    to_std_logic_vector(to_signed(-602,SDLEN)),
    to_std_logic_vector(to_signed(-567,SDLEN)),
    to_std_logic_vector(to_signed(-500,SDLEN)),
    to_std_logic_vector(to_signed(-402,SDLEN)),
    to_std_logic_vector(to_signed(-280,SDLEN)),
    to_std_logic_vector(to_signed(-139,SDLEN)),
    to_std_logic_vector(to_signed(12,SDLEN)),
    to_std_logic_vector(to_signed(166,SDLEN)),
    to_std_logic_vector(to_signed(313,SDLEN)),
    to_std_logic_vector(to_signed(444,SDLEN)),
    to_std_logic_vector(to_signed(550,SDLEN)),
    to_std_logic_vector(to_signed(623,SDLEN)),
    to_std_logic_vector(to_signed(-24229,SDLEN)),
    to_std_logic_vector(to_signed(18148,SDLEN)),
    to_std_logic_vector(to_signed(7402,SDLEN)),
    to_std_logic_vector(to_signed(25047,SDLEN)),
    to_std_logic_vector(to_signed(-10473,SDLEN)),
    to_std_logic_vector(to_signed(658,SDLEN)),
    to_std_logic_vector(to_signed(651,SDLEN)),
    to_std_logic_vector(to_signed(602,SDLEN)),
    to_std_logic_vector(to_signed(512,SDLEN)),
    to_std_logic_vector(to_signed(386,SDLEN)),
    to_std_logic_vector(to_signed(232,SDLEN)),
    to_std_logic_vector(to_signed(59,SDLEN)),
    to_std_logic_vector(to_signed(-120,SDLEN)),
    to_std_logic_vector(to_signed(-295,SDLEN)),
    to_std_logic_vector(to_signed(-452,SDLEN)),
    to_std_logic_vector(to_signed(-579,SDLEN)),
    to_std_logic_vector(to_signed(-667,SDLEN)),
    to_std_logic_vector(to_signed(-707,SDLEN)),
    to_std_logic_vector(to_signed(-696,SDLEN)),
    to_std_logic_vector(to_signed(-632,SDLEN)),
    to_std_logic_vector(to_signed(-519,SDLEN)),
    to_std_logic_vector(to_signed(-364,SDLEN)),
    to_std_logic_vector(to_signed(-179,SDLEN)),
    to_std_logic_vector(to_signed(23,SDLEN)),
    to_std_logic_vector(to_signed(227,SDLEN)),
    to_std_logic_vector(to_signed(417,SDLEN)),
    to_std_logic_vector(to_signed(575,SDLEN)),
    to_std_logic_vector(to_signed(690,SDLEN)),
    to_std_logic_vector(to_signed(748,SDLEN)),
    to_std_logic_vector(to_signed(745,SDLEN)),
    to_std_logic_vector(to_signed(679,SDLEN)),
    to_std_logic_vector(to_signed(554,SDLEN)),
    to_std_logic_vector(to_signed(379,SDLEN)),
    to_std_logic_vector(to_signed(168,SDLEN)),
    to_std_logic_vector(to_signed(-61,SDLEN)),
    to_std_logic_vector(to_signed(-288,SDLEN)),
    to_std_logic_vector(to_signed(-493,SDLEN)),
    to_std_logic_vector(to_signed(-656,SDLEN)),
    to_std_logic_vector(to_signed(-762,SDLEN)),
    to_std_logic_vector(to_signed(-798,SDLEN)),
    to_std_logic_vector(to_signed(-760,SDLEN)),
    to_std_logic_vector(to_signed(-649,SDLEN)),
    to_std_logic_vector(to_signed(-474,SDLEN)),
    to_std_logic_vector(to_signed(-251,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(255,SDLEN)),
    to_std_logic_vector(to_signed(488,SDLEN)),
    to_std_logic_vector(to_signed(676,SDLEN)),
    to_std_logic_vector(to_signed(797,SDLEN)),
    to_std_logic_vector(to_signed(839,SDLEN)),
    to_std_logic_vector(to_signed(794,SDLEN)),
    to_std_logic_vector(to_signed(666,SDLEN)),
    to_std_logic_vector(to_signed(465,SDLEN)),
    to_std_logic_vector(to_signed(212,SDLEN)),
    to_std_logic_vector(to_signed(-67,SDLEN)),
    to_std_logic_vector(to_signed(-343,SDLEN)),
    to_std_logic_vector(to_signed(-586,SDLEN)),
    to_std_logic_vector(to_signed(-767,SDLEN)),
    to_std_logic_vector(to_signed(-865,SDLEN)),
    to_std_logic_vector(to_signed(-866,SDLEN)),
    to_std_logic_vector(to_signed(-769,SDLEN)),
    to_std_logic_vector(to_signed(-583,SDLEN)),
    to_std_logic_vector(to_signed(-326,SDLEN)),
    to_std_logic_vector(to_signed(-27,SDLEN)),
    to_std_logic_vector(to_signed(278,SDLEN)),
    to_std_logic_vector(to_signed(555,SDLEN)),
    to_std_logic_vector(to_signed(769,SDLEN)),
    to_std_logic_vector(to_signed(892,SDLEN)),
    to_std_logic_vector(to_signed(908,SDLEN)),
    to_std_logic_vector(to_signed(812,SDLEN)),
    to_std_logic_vector(to_signed(614,SDLEN)),
    to_std_logic_vector(to_signed(336,SDLEN)),
    to_std_logic_vector(to_signed(11,SDLEN)),
    to_std_logic_vector(to_signed(-318,SDLEN)),
    to_std_logic_vector(to_signed(-611,SDLEN)),
    to_std_logic_vector(to_signed(-829,SDLEN)),
    to_std_logic_vector(to_signed(-941,SDLEN)),
    to_std_logic_vector(to_signed(-929,SDLEN)),
    to_std_logic_vector(to_signed(-794,SDLEN)),
    to_std_logic_vector(to_signed(-550,SDLEN)),
    to_std_logic_vector(to_signed(-228,SDLEN)),
    to_std_logic_vector(to_signed(128,SDLEN)),
    to_std_logic_vector(to_signed(472,SDLEN)),
    to_std_logic_vector(to_signed(754,SDLEN)),
    to_std_logic_vector(to_signed(934,SDLEN)),
    to_std_logic_vector(to_signed(-24141,SDLEN)),
    to_std_logic_vector(to_signed(16505,SDLEN)),
    to_std_logic_vector(to_signed(-28462,SDLEN)),
    to_std_logic_vector(to_signed(-16873,SDLEN)),
    to_std_logic_vector(to_signed(20964,SDLEN)),
    to_std_logic_vector(to_signed(985,SDLEN)),
    to_std_logic_vector(to_signed(895,SDLEN)),
    to_std_logic_vector(to_signed(676,SDLEN)),
    to_std_logic_vector(to_signed(356,SDLEN)),
    to_std_logic_vector(to_signed(-19,SDLEN)),
    to_std_logic_vector(to_signed(-397,SDLEN)),
    to_std_logic_vector(to_signed(-720,SDLEN)),
    to_std_logic_vector(to_signed(-939,SDLEN)),
    to_std_logic_vector(to_signed(-1019,SDLEN)),
    to_std_logic_vector(to_signed(-946,SDLEN)),
    to_std_logic_vector(to_signed(-726,SDLEN)),
    to_std_logic_vector(to_signed(-392,SDLEN)),
    to_std_logic_vector(to_signed(7,SDLEN)),
    to_std_logic_vector(to_signed(410,SDLEN)),
    to_std_logic_vector(to_signed(752,SDLEN)),
    to_std_logic_vector(to_signed(979,SDLEN)),
    to_std_logic_vector(to_signed(1051,SDLEN)),
    to_std_logic_vector(to_signed(954,SDLEN)),
    to_std_logic_vector(to_signed(700,SDLEN)),
    to_std_logic_vector(to_signed(329,SDLEN)),
    to_std_logic_vector(to_signed(-101,SDLEN)),
    to_std_logic_vector(to_signed(-519,SDLEN)),
    to_std_logic_vector(to_signed(-855,SDLEN)),
    to_std_logic_vector(to_signed(-1050,SDLEN)),
    to_std_logic_vector(to_signed(-1068,SDLEN)),
    to_std_logic_vector(to_signed(-903,SDLEN)),
    to_std_logic_vector(to_signed(-579,SDLEN)),
    to_std_logic_vector(to_signed(-151,SDLEN)),
    to_std_logic_vector(to_signed(308,SDLEN)),
    to_std_logic_vector(to_signed(718,SDLEN)),
    to_std_logic_vector(to_signed(1004,SDLEN)),
    to_std_logic_vector(to_signed(1114,SDLEN)),
    to_std_logic_vector(to_signed(1023,SDLEN)),
    to_std_logic_vector(to_signed(744,SDLEN)),
    to_std_logic_vector(to_signed(326,SDLEN)),
    to_std_logic_vector(to_signed(-155,SDLEN)),
    to_std_logic_vector(to_signed(-614,SDLEN)),
    to_std_logic_vector(to_signed(-963,SDLEN)),
    to_std_logic_vector(to_signed(-1133,SDLEN)),
    to_std_logic_vector(to_signed(-1090,SDLEN)),
    to_std_logic_vector(to_signed(-838,SDLEN)),
    to_std_logic_vector(to_signed(-421,SDLEN)),
    to_std_logic_vector(to_signed(80,SDLEN)),
    to_std_logic_vector(to_signed(573,SDLEN)),
    to_std_logic_vector(to_signed(957,SDLEN)),
    to_std_logic_vector(to_signed(1156,SDLEN)),
    to_std_logic_vector(to_signed(1126,SDLEN)),
    to_std_logic_vector(to_signed(870,SDLEN)),
    to_std_logic_vector(to_signed(434,SDLEN)),
    to_std_logic_vector(to_signed(-93,SDLEN)),
    to_std_logic_vector(to_signed(-607,SDLEN)),
    to_std_logic_vector(to_signed(-1001,SDLEN)),
    to_std_logic_vector(to_signed(-1191,SDLEN)),
    to_std_logic_vector(to_signed(-1134,SDLEN)),
    to_std_logic_vector(to_signed(-837,SDLEN)),
    to_std_logic_vector(to_signed(-360,SDLEN)),
    to_std_logic_vector(to_signed(198,SDLEN)),
    to_std_logic_vector(to_signed(720,SDLEN)),
    to_std_logic_vector(to_signed(1091,SDLEN)),
    to_std_logic_vector(to_signed(1228,SDLEN)),
    to_std_logic_vector(to_signed(1098,SDLEN)),
    to_std_logic_vector(to_signed(723,SDLEN)),
    to_std_logic_vector(to_signed(185,SDLEN)),
    to_std_logic_vector(to_signed(-399,SDLEN)),
    to_std_logic_vector(to_signed(-900,SDLEN)),
    to_std_logic_vector(to_signed(-1202,SDLEN)),
    to_std_logic_vector(to_signed(-1233,SDLEN)),
    to_std_logic_vector(to_signed(-982,SDLEN)),
    to_std_logic_vector(to_signed(-501,SDLEN)),
    to_std_logic_vector(to_signed(99,SDLEN)),
    to_std_logic_vector(to_signed(683,SDLEN)),
    to_std_logic_vector(to_signed(1112,SDLEN)),
    to_std_logic_vector(to_signed(1281,SDLEN)),
    to_std_logic_vector(to_signed(1147,SDLEN)),
    to_std_logic_vector(to_signed(737,SDLEN)),
    to_std_logic_vector(to_signed(146,SDLEN)),
    to_std_logic_vector(to_signed(-486,SDLEN)),
    to_std_logic_vector(to_signed(-1006,SDLEN)),
    to_std_logic_vector(to_signed(-1283,SDLEN)),
    to_std_logic_vector(to_signed(-1246,SDLEN)),
    to_std_logic_vector(to_signed(-32313,SDLEN)),
    to_std_logic_vector(to_signed(-14461,SDLEN)),
    to_std_logic_vector(to_signed(-23925,SDLEN)),
    to_std_logic_vector(to_signed(-15334,SDLEN)),
    to_std_logic_vector(to_signed(15774,SDLEN)),
    to_std_logic_vector(to_signed(-899,SDLEN)),
    to_std_logic_vector(to_signed(-323,SDLEN)),
    to_std_logic_vector(to_signed(338,SDLEN)),
    to_std_logic_vector(to_signed(920,SDLEN)),
    to_std_logic_vector(to_signed(1273,SDLEN)),
    to_std_logic_vector(to_signed(1304,SDLEN)),
    to_std_logic_vector(to_signed(998,SDLEN)),
    to_std_logic_vector(to_signed(431,SDLEN)),
    to_std_logic_vector(to_signed(-253,SDLEN)),
    to_std_logic_vector(to_signed(-877,SDLEN)),
    to_std_logic_vector(to_signed(-1275,SDLEN)),
    to_std_logic_vector(to_signed(-1338,SDLEN)),
    to_std_logic_vector(to_signed(-1044,SDLEN)),
    to_std_logic_vector(to_signed(-467,SDLEN)),
    to_std_logic_vector(to_signed(241,SDLEN)),
    to_std_logic_vector(to_signed(890,SDLEN)),
    to_std_logic_vector(to_signed(1302,SDLEN)),
    to_std_logic_vector(to_signed(1359,SDLEN)),
    to_std_logic_vector(to_signed(1040,SDLEN)),
    to_std_logic_vector(to_signed(430,SDLEN)),
    to_std_logic_vector(to_signed(-305,SDLEN)),
    to_std_logic_vector(to_signed(-962,SDLEN)),
    to_std_logic_vector(to_signed(-1351,SDLEN)),
    to_std_logic_vector(to_signed(-1360,SDLEN)),
    to_std_logic_vector(to_signed(-979,SDLEN)),
    to_std_logic_vector(to_signed(-313,SDLEN)),
    to_std_logic_vector(to_signed(448,SDLEN)),
    to_std_logic_vector(to_signed(1086,SDLEN)),
    to_std_logic_vector(to_signed(1412,SDLEN)),
    to_std_logic_vector(to_signed(1324,SDLEN)),
    to_std_logic_vector(to_signed(844,SDLEN)),
    to_std_logic_vector(to_signed(108,SDLEN)),
    to_std_logic_vector(to_signed(-665,SDLEN)),
    to_std_logic_vector(to_signed(-1245,SDLEN)),
    to_std_logic_vector(to_signed(-1453,SDLEN)),
    to_std_logic_vector(to_signed(-1221,SDLEN)),
    to_std_logic_vector(to_signed(-613,SDLEN)),
    to_std_logic_vector(to_signed(188,SDLEN)),
    to_std_logic_vector(to_signed(938,SDLEN)),
    to_std_logic_vector(to_signed(1402,SDLEN)),
    to_std_logic_vector(to_signed(1431,SDLEN)),
    to_std_logic_vector(to_signed(1011,SDLEN)),
    to_std_logic_vector(to_signed(268,SDLEN)),
    to_std_logic_vector(to_signed(-566,SDLEN)),
    to_std_logic_vector(to_signed(-1226,SDLEN)),
    to_std_logic_vector(to_signed(-1498,SDLEN)),
    to_std_logic_vector(to_signed(-1288,SDLEN)),
    to_std_logic_vector(to_signed(-658,SDLEN)),
    to_std_logic_vector(to_signed(190,SDLEN)),
    to_std_logic_vector(to_signed(984,SDLEN)),
    to_std_logic_vector(to_signed(1459,SDLEN)),
    to_std_logic_vector(to_signed(1454,SDLEN)),
    to_std_logic_vector(to_signed(965,SDLEN)),
    to_std_logic_vector(to_signed(148,SDLEN)),
    to_std_logic_vector(to_signed(-724,SDLEN)),
    to_std_logic_vector(to_signed(-1358,SDLEN)),
    to_std_logic_vector(to_signed(-1536,SDLEN)),
    to_std_logic_vector(to_signed(-1189,SDLEN)),
    to_std_logic_vector(to_signed(-431,SDLEN)),
    to_std_logic_vector(to_signed(480,SDLEN)),
    to_std_logic_vector(to_signed(1233,SDLEN)),
    to_std_logic_vector(to_signed(1561,SDLEN)),
    to_std_logic_vector(to_signed(1344,SDLEN)),
    to_std_logic_vector(to_signed(651,SDLEN)),
    to_std_logic_vector(to_signed(-277,SDLEN)),
    to_std_logic_vector(to_signed(-1114,SDLEN)),
    to_std_logic_vector(to_signed(-1559,SDLEN)),
    to_std_logic_vector(to_signed(-1446,SDLEN)),
    to_std_logic_vector(to_signed(-810,SDLEN)),
    to_std_logic_vector(to_signed(125,SDLEN)),
    to_std_logic_vector(to_signed(1021,SDLEN)),
    to_std_logic_vector(to_signed(1550,SDLEN)),
    to_std_logic_vector(to_signed(1510,SDLEN)),
    to_std_logic_vector(to_signed(911,SDLEN)),
    to_std_logic_vector(to_signed(-31,SDLEN)),
    to_std_logic_vector(to_signed(-969,SDLEN)),
    to_std_logic_vector(to_signed(-1550,SDLEN)),
    to_std_logic_vector(to_signed(-1548,SDLEN)),
    to_std_logic_vector(to_signed(-959,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN))
  );

  constant STO_ROM_INIT_DATA : ROM_DATA_T := (
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(4,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(3,SDLEN)),
    to_std_logic_vector(to_signed(1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(0,SDLEN)),
    to_std_logic_vector(to_signed(15,SDLEN)),
    to_std_logic_vector(to_signed(33,SDLEN)),
    to_std_logic_vector(to_signed(51,SDLEN)),
    to_std_logic_vector(to_signed(51,SDLEN)),
    to_std_logic_vector(to_signed(52,SDLEN)),
    to_std_logic_vector(to_signed(51,SDLEN)),
    to_std_logic_vector(to_signed(51,SDLEN)),
    to_std_logic_vector(to_signed(47,SDLEN)),
    to_std_logic_vector(to_signed(56,SDLEN)),
    to_std_logic_vector(to_signed(50,SDLEN)),
    to_std_logic_vector(to_signed(43,SDLEN)),
    to_std_logic_vector(to_signed(-5752,SDLEN)),
    to_std_logic_vector(to_signed(160,SDLEN)),
    to_std_logic_vector(to_signed(250,SDLEN)),
    to_std_logic_vector(to_signed(-15681,SDLEN)),
    to_std_logic_vector(to_signed(-18462,SDLEN)),
    to_std_logic_vector(to_signed(37,SDLEN)),
    to_std_logic_vector(to_signed(26,SDLEN)),
    to_std_logic_vector(to_signed(19,SDLEN)),
    to_std_logic_vector(to_signed(5,SDLEN)),
    to_std_logic_vector(to_signed(-5,SDLEN)),
    to_std_logic_vector(to_signed(-16,SDLEN)),
    to_std_logic_vector(to_signed(-27,SDLEN)),
    to_std_logic_vector(to_signed(-38,SDLEN)),
    to_std_logic_vector(to_signed(-45,SDLEN)),
    to_std_logic_vector(to_signed(-51,SDLEN)),
    to_std_logic_vector(to_signed(-54,SDLEN)),
    to_std_logic_vector(to_signed(-56,SDLEN)),
    to_std_logic_vector(to_signed(-57,SDLEN)),
    to_std_logic_vector(to_signed(-56,SDLEN)),
    to_std_logic_vector(to_signed(-53,SDLEN)),
    to_std_logic_vector(to_signed(-50,SDLEN)),
    to_std_logic_vector(to_signed(-75,SDLEN)),
    to_std_logic_vector(to_signed(-78,SDLEN)),
    to_std_logic_vector(to_signed(-86,SDLEN)),
    to_std_logic_vector(to_signed(-85,SDLEN)),
    to_std_logic_vector(to_signed(-85,SDLEN)),
    to_std_logic_vector(to_signed(-82,SDLEN)),
    to_std_logic_vector(to_signed(-100,SDLEN)),
    to_std_logic_vector(to_signed(-96,SDLEN)),
    to_std_logic_vector(to_signed(-94,SDLEN)),
    to_std_logic_vector(to_signed(-116,SDLEN)),
    to_std_logic_vector(to_signed(-114,SDLEN)),
    to_std_logic_vector(to_signed(-113,SDLEN)),
    to_std_logic_vector(to_signed(-131,SDLEN)),
    to_std_logic_vector(to_signed(-123,SDLEN)),
    to_std_logic_vector(to_signed(-117,SDLEN)),
    to_std_logic_vector(to_signed(-102,SDLEN)),
    to_std_logic_vector(to_signed(-82,SDLEN)),
    to_std_logic_vector(to_signed(-57,SDLEN)),
    to_std_logic_vector(to_signed(-30,SDLEN)),
    to_std_logic_vector(to_signed(-1,SDLEN)),
    to_std_logic_vector(to_signed(25,SDLEN)),
    to_std_logic_vector(to_signed(52,SDLEN)),
    to_std_logic_vector(to_signed(74,SDLEN)),
    to_std_logic_vector(to_signed(94,SDLEN)),
    to_std_logic_vector(to_signed(118,SDLEN)),
    to_std_logic_vector(to_signed(145,SDLEN)),
    to_std_logic_vector(to_signed(171,SDLEN)),
    to_std_logic_vector(to_signed(196,SDLEN)),
    to_std_logic_vector(to_signed(218,SDLEN)),
    to_std_logic_vector(to_signed(240,SDLEN)),
    to_std_logic_vector(to_signed(255,SDLEN)),
    to_std_logic_vector(to_signed(264,SDLEN)),
    to_std_logic_vector(to_signed(267,SDLEN)),
    to_std_logic_vector(to_signed(260,SDLEN)),
    to_std_logic_vector(to_signed(264,SDLEN)),
    to_std_logic_vector(to_signed(254,SDLEN)),
    to_std_logic_vector(to_signed(240,SDLEN)),
    to_std_logic_vector(to_signed(220,SDLEN)),
    to_std_logic_vector(to_signed(214,SDLEN)),
    to_std_logic_vector(to_signed(194,SDLEN)),
    to_std_logic_vector(to_signed(172,SDLEN)),
    to_std_logic_vector(to_signed(145,SDLEN)),
    to_std_logic_vector(to_signed(112,SDLEN)),
    to_std_logic_vector(to_signed(79,SDLEN)),
    to_std_logic_vector(to_signed(38,SDLEN)),
    to_std_logic_vector(to_signed(-5,SDLEN)),
    to_std_logic_vector(to_signed(-48,SDLEN)),
    to_std_logic_vector(to_signed(-90,SDLEN)),
    to_std_logic_vector(to_signed(-144,SDLEN)),
    to_std_logic_vector(to_signed(-188,SDLEN)),
    to_std_logic_vector(to_signed(-244,SDLEN)),
    to_std_logic_vector(to_signed(-296,SDLEN)),
    to_std_logic_vector(to_signed(-343,SDLEN)),
    to_std_logic_vector(to_signed(-381,SDLEN)),
    to_std_logic_vector(to_signed(-421,SDLEN)),
    to_std_logic_vector(to_signed(-443,SDLEN)),
    to_std_logic_vector(to_signed(-450,SDLEN)),
    to_std_logic_vector(to_signed(-463,SDLEN)),
    to_std_logic_vector(to_signed(-454,SDLEN)),
    to_std_logic_vector(to_signed(-428,SDLEN)),
    to_std_logic_vector(to_signed(-415,SDLEN)),
    to_std_logic_vector(to_signed(-359,SDLEN)),
    to_std_logic_vector(to_signed(-303,SDLEN)),
    to_std_logic_vector(to_signed(-249,SDLEN)),
    to_std_logic_vector(to_signed(-29314,SDLEN)),
    to_std_logic_vector(to_signed(6197,SDLEN)),
    to_std_logic_vector(to_signed(7439,SDLEN)),
    to_std_logic_vector(to_signed(-11681,SDLEN)),
    to_std_logic_vector(to_signed(22234,SDLEN)),
    to_std_logic_vector(to_signed(-138,SDLEN)),
    to_std_logic_vector(to_signed(-34,SDLEN)),
    to_std_logic_vector(to_signed(96,SDLEN)),
    to_std_logic_vector(to_signed(210,SDLEN)),
    to_std_logic_vector(to_signed(310,SDLEN)),
    to_std_logic_vector(to_signed(405,SDLEN)),
    to_std_logic_vector(to_signed(475,SDLEN)),
    to_std_logic_vector(to_signed(521,SDLEN)),
    to_std_logic_vector(to_signed(561,SDLEN)),
    to_std_logic_vector(to_signed(570,SDLEN)),
    to_std_logic_vector(to_signed(558,SDLEN)),
    to_std_logic_vector(to_signed(529,SDLEN)),
    to_std_logic_vector(to_signed(473,SDLEN)),
    to_std_logic_vector(to_signed(405,SDLEN)),
    to_std_logic_vector(to_signed(310,SDLEN)),
    to_std_logic_vector(to_signed(196,SDLEN)),
    to_std_logic_vector(to_signed(92,SDLEN)),
    to_std_logic_vector(to_signed(-28,SDLEN)),
    to_std_logic_vector(to_signed(-142,SDLEN)),
    to_std_logic_vector(to_signed(-246,SDLEN)),
    to_std_logic_vector(to_signed(-347,SDLEN)),
    to_std_logic_vector(to_signed(-431,SDLEN)),
    to_std_logic_vector(to_signed(-505,SDLEN)),
    to_std_logic_vector(to_signed(-548,SDLEN)),
    to_std_logic_vector(to_signed(-583,SDLEN)),
    to_std_logic_vector(to_signed(-586,SDLEN)),
    to_std_logic_vector(to_signed(-549,SDLEN)),
    to_std_logic_vector(to_signed(-512,SDLEN)),
    to_std_logic_vector(to_signed(-437,SDLEN)),
    to_std_logic_vector(to_signed(-355,SDLEN)),
    to_std_logic_vector(to_signed(-244,SDLEN)),
    to_std_logic_vector(to_signed(-120,SDLEN)),
    to_std_logic_vector(to_signed(2,SDLEN)),
    to_std_logic_vector(to_signed(140,SDLEN)),
    to_std_logic_vector(to_signed(264,SDLEN)),
    to_std_logic_vector(to_signed(375,SDLEN)),
    to_std_logic_vector(to_signed(480,SDLEN)),
    to_std_logic_vector(to_signed(551,SDLEN)),
    to_std_logic_vector(to_signed(600,SDLEN)),
    to_std_logic_vector(to_signed(629,SDLEN)),
    to_std_logic_vector(to_signed(573,SDLEN)),
    to_std_logic_vector(to_signed(491,SDLEN)),
    to_std_logic_vector(to_signed(373,SDLEN)),
    to_std_logic_vector(to_signed(225,SDLEN)),
    to_std_logic_vector(to_signed(63,SDLEN)),
    to_std_logic_vector(to_signed(-103,SDLEN)),
    to_std_logic_vector(to_signed(-247,SDLEN)),
    to_std_logic_vector(to_signed(-383,SDLEN)),
    to_std_logic_vector(to_signed(-468,SDLEN)),
    to_std_logic_vector(to_signed(-509,SDLEN)),
    to_std_logic_vector(to_signed(-530,SDLEN)),
    to_std_logic_vector(to_signed(-510,SDLEN)),
    to_std_logic_vector(to_signed(-460,SDLEN)),
    to_std_logic_vector(to_signed(-355,SDLEN)),
    to_std_logic_vector(to_signed(-229,SDLEN)),
    to_std_logic_vector(to_signed(-82,SDLEN)),
    to_std_logic_vector(to_signed(74,SDLEN)),
    to_std_logic_vector(to_signed(232,SDLEN)),
    to_std_logic_vector(to_signed(373,SDLEN)),
    to_std_logic_vector(to_signed(502,SDLEN)),
    to_std_logic_vector(to_signed(593,SDLEN)),
    to_std_logic_vector(to_signed(655,SDLEN)),
    to_std_logic_vector(to_signed(670,SDLEN)),
    to_std_logic_vector(to_signed(638,SDLEN)),
    to_std_logic_vector(to_signed(571,SDLEN)),
    to_std_logic_vector(to_signed(455,SDLEN)),
    to_std_logic_vector(to_signed(310,SDLEN)),
    to_std_logic_vector(to_signed(138,SDLEN)),
    to_std_logic_vector(to_signed(-43,SDLEN)),
    to_std_logic_vector(to_signed(-221,SDLEN)),
    to_std_logic_vector(to_signed(-380,SDLEN)),
    to_std_logic_vector(to_signed(-488,SDLEN)),
    to_std_logic_vector(to_signed(-555,SDLEN)),
    to_std_logic_vector(to_signed(-595,SDLEN)),
    to_std_logic_vector(to_signed(-581,SDLEN)),
    to_std_logic_vector(to_signed(-521,SDLEN)),
    to_std_logic_vector(to_signed(-396,SDLEN)),
    to_std_logic_vector(to_signed(-246,SDLEN)),
    to_std_logic_vector(to_signed(-72,SDLEN)),
    to_std_logic_vector(to_signed(111,SDLEN)),
    to_std_logic_vector(to_signed(-24229,SDLEN)),
    to_std_logic_vector(to_signed(18148,SDLEN)),
    to_std_logic_vector(to_signed(7402,SDLEN)),
    to_std_logic_vector(to_signed(25047,SDLEN)),
    to_std_logic_vector(to_signed(-10473,SDLEN)),
    to_std_logic_vector(to_signed(303,SDLEN)),
    to_std_logic_vector(to_signed(451,SDLEN)),
    to_std_logic_vector(to_signed(545,SDLEN)),
    to_std_logic_vector(to_signed(579,SDLEN)),
    to_std_logic_vector(to_signed(534,SDLEN)),
    to_std_logic_vector(to_signed(409,SDLEN)),
    to_std_logic_vector(to_signed(228,SDLEN)),
    to_std_logic_vector(to_signed(10,SDLEN)),
    to_std_logic_vector(to_signed(-214,SDLEN)),
    to_std_logic_vector(to_signed(-421,SDLEN)),
    to_std_logic_vector(to_signed(-569,SDLEN)),
    to_std_logic_vector(to_signed(-659,SDLEN)),
    to_std_logic_vector(to_signed(-698,SDLEN)),
    to_std_logic_vector(to_signed(-674,SDLEN)),
    to_std_logic_vector(to_signed(-584,SDLEN)),
    to_std_logic_vector(to_signed(-414,SDLEN)),
    to_std_logic_vector(to_signed(-184,SDLEN)),
    to_std_logic_vector(to_signed(68,SDLEN)),
    to_std_logic_vector(to_signed(333,SDLEN)),
    to_std_logic_vector(to_signed(566,SDLEN)),
    to_std_logic_vector(to_signed(752,SDLEN)),
    to_std_logic_vector(to_signed(854,SDLEN)),
    to_std_logic_vector(to_signed(868,SDLEN)),
    to_std_logic_vector(to_signed(800,SDLEN)),
    to_std_logic_vector(to_signed(635,SDLEN)),
    to_std_logic_vector(to_signed(398,SDLEN)),
    to_std_logic_vector(to_signed(112,SDLEN)),
    to_std_logic_vector(to_signed(-183,SDLEN)),
    to_std_logic_vector(to_signed(-456,SDLEN)),
    to_std_logic_vector(to_signed(-674,SDLEN)),
    to_std_logic_vector(to_signed(-800,SDLEN)),
    to_std_logic_vector(to_signed(-851,SDLEN)),
    to_std_logic_vector(to_signed(-815,SDLEN)),
    to_std_logic_vector(to_signed(-686,SDLEN)),
    to_std_logic_vector(to_signed(-476,SDLEN)),
    to_std_logic_vector(to_signed(-184,SDLEN)),
    to_std_logic_vector(to_signed(134,SDLEN)),
    to_std_logic_vector(to_signed(445,SDLEN)),
    to_std_logic_vector(to_signed(715,SDLEN)),
    to_std_logic_vector(to_signed(897,SDLEN)),
    to_std_logic_vector(to_signed(944,SDLEN)),
    to_std_logic_vector(to_signed(851,SDLEN)),
    to_std_logic_vector(to_signed(641,SDLEN)),
    to_std_logic_vector(to_signed(351,SDLEN)),
    to_std_logic_vector(to_signed(-65,SDLEN)),
    to_std_logic_vector(to_signed(-454,SDLEN)),
    to_std_logic_vector(to_signed(-807,SDLEN)),
    to_std_logic_vector(to_signed(-1051,SDLEN)),
    to_std_logic_vector(to_signed(-1156,SDLEN)),
    to_std_logic_vector(to_signed(-1087,SDLEN)),
    to_std_logic_vector(to_signed(-774,SDLEN)),
    to_std_logic_vector(to_signed(-354,SDLEN)),
    to_std_logic_vector(to_signed(152,SDLEN)),
    to_std_logic_vector(to_signed(637,SDLEN)),
    to_std_logic_vector(to_signed(1012,SDLEN)),
    to_std_logic_vector(to_signed(1191,SDLEN)),
    to_std_logic_vector(to_signed(1161,SDLEN)),
    to_std_logic_vector(to_signed(847,SDLEN)),
    to_std_logic_vector(to_signed(392,SDLEN)),
    to_std_logic_vector(to_signed(-150,SDLEN)),
    to_std_logic_vector(to_signed(-646,SDLEN)),
    to_std_logic_vector(to_signed(-1006,SDLEN)),
    to_std_logic_vector(to_signed(-1141,SDLEN)),
    to_std_logic_vector(to_signed(-1046,SDLEN)),
    to_std_logic_vector(to_signed(-755,SDLEN)),
    to_std_logic_vector(to_signed(-346,SDLEN)),
    to_std_logic_vector(to_signed(177,SDLEN)),
    to_std_logic_vector(to_signed(626,SDLEN)),
    to_std_logic_vector(to_signed(967,SDLEN)),
    to_std_logic_vector(to_signed(1133,SDLEN)),
    to_std_logic_vector(to_signed(1112,SDLEN)),
    to_std_logic_vector(to_signed(909,SDLEN)),
    to_std_logic_vector(to_signed(591,SDLEN)),
    to_std_logic_vector(to_signed(156,SDLEN)),
    to_std_logic_vector(to_signed(-256,SDLEN)),
    to_std_logic_vector(to_signed(-612,SDLEN)),
    to_std_logic_vector(to_signed(-844,SDLEN)),
    to_std_logic_vector(to_signed(-934,SDLEN)),
    to_std_logic_vector(to_signed(-870,SDLEN)),
    to_std_logic_vector(to_signed(-616,SDLEN)),
    to_std_logic_vector(to_signed(-24141,SDLEN)),
    to_std_logic_vector(to_signed(16505,SDLEN)),
    to_std_logic_vector(to_signed(-28462,SDLEN)),
    to_std_logic_vector(to_signed(-16873,SDLEN)),
    to_std_logic_vector(to_signed(20964,SDLEN)),
    to_std_logic_vector(to_signed(-220,SDLEN)),
    to_std_logic_vector(to_signed(225,SDLEN)),
    to_std_logic_vector(to_signed(618,SDLEN)),
    to_std_logic_vector(to_signed(854,SDLEN)),
    to_std_logic_vector(to_signed(909,SDLEN)),
    to_std_logic_vector(to_signed(738,SDLEN)),
    to_std_logic_vector(to_signed(394,SDLEN)),
    to_std_logic_vector(to_signed(-60,SDLEN)),
    to_std_logic_vector(to_signed(-498,SDLEN)),
    to_std_logic_vector(to_signed(-846,SDLEN)),
    to_std_logic_vector(to_signed(-1033,SDLEN)),
    to_std_logic_vector(to_signed(-1018,SDLEN)),
    to_std_logic_vector(to_signed(-818,SDLEN)),
    to_std_logic_vector(to_signed(-484,SDLEN)),
    to_std_logic_vector(to_signed(-59,SDLEN)),
    to_std_logic_vector(to_signed(367,SDLEN)),
    to_std_logic_vector(to_signed(721,SDLEN)),
    to_std_logic_vector(to_signed(932,SDLEN)),
    to_std_logic_vector(to_signed(977,SDLEN)),
    to_std_logic_vector(to_signed(837,SDLEN)),
    to_std_logic_vector(to_signed(554,SDLEN)),
    to_std_logic_vector(to_signed(146,SDLEN)),
    to_std_logic_vector(to_signed(-288,SDLEN)),
    to_std_logic_vector(to_signed(-685,SDLEN)),
    to_std_logic_vector(to_signed(-947,SDLEN)),
    to_std_logic_vector(to_signed(-1035,SDLEN)),
    to_std_logic_vector(to_signed(-918,SDLEN)),
    to_std_logic_vector(to_signed(-615,SDLEN)),
    to_std_logic_vector(to_signed(-182,SDLEN)),
    to_std_logic_vector(to_signed(305,SDLEN)),
    to_std_logic_vector(to_signed(729,SDLEN)),
    to_std_logic_vector(to_signed(1004,SDLEN)),
    to_std_logic_vector(to_signed(1050,SDLEN)),
    to_std_logic_vector(to_signed(874,SDLEN)),
    to_std_logic_vector(to_signed(502,SDLEN)),
    to_std_logic_vector(to_signed(13,SDLEN)),
    to_std_logic_vector(to_signed(-483,SDLEN)),
    to_std_logic_vector(to_signed(-863,SDLEN)),
    to_std_logic_vector(to_signed(-1063,SDLEN)),
    to_std_logic_vector(to_signed(-1037,SDLEN)),
    to_std_logic_vector(to_signed(-665,SDLEN)),
    to_std_logic_vector(to_signed(-124,SDLEN)),
    to_std_logic_vector(to_signed(447,SDLEN)),
    to_std_logic_vector(to_signed(880,SDLEN)),
    to_std_logic_vector(to_signed(1065,SDLEN)),
    to_std_logic_vector(to_signed(932,SDLEN)),
    to_std_logic_vector(to_signed(529,SDLEN)),
    to_std_logic_vector(to_signed(-39,SDLEN)),
    to_std_logic_vector(to_signed(-614,SDLEN)),
    to_std_logic_vector(to_signed(-1032,SDLEN)),
    to_std_logic_vector(to_signed(-1167,SDLEN)),
    to_std_logic_vector(to_signed(-985,SDLEN)),
    to_std_logic_vector(to_signed(-527,SDLEN)),
    to_std_logic_vector(to_signed(105,SDLEN)),
    to_std_logic_vector(to_signed(728,SDLEN)),
    to_std_logic_vector(to_signed(1176,SDLEN)),
    to_std_logic_vector(to_signed(1306,SDLEN)),
    to_std_logic_vector(to_signed(1079,SDLEN)),
    to_std_logic_vector(to_signed(572,SDLEN)),
    to_std_logic_vector(to_signed(-88,SDLEN)),
    to_std_logic_vector(to_signed(-723,SDLEN)),
    to_std_logic_vector(to_signed(-1162,SDLEN)),
    to_std_logic_vector(to_signed(-1280,SDLEN)),
    to_std_logic_vector(to_signed(-1073,SDLEN)),
    to_std_logic_vector(to_signed(-575,SDLEN)),
    to_std_logic_vector(to_signed(86,SDLEN)),
    to_std_logic_vector(to_signed(727,SDLEN)),
    to_std_logic_vector(to_signed(1173,SDLEN)),
    to_std_logic_vector(to_signed(1319,SDLEN)),
    to_std_logic_vector(to_signed(1113,SDLEN)),
    to_std_logic_vector(to_signed(610,SDLEN)),
    to_std_logic_vector(to_signed(-56,SDLEN)),
    to_std_logic_vector(to_signed(-705,SDLEN)),
    to_std_logic_vector(to_signed(-1155,SDLEN)),
    to_std_logic_vector(to_signed(-1279,SDLEN)),
    to_std_logic_vector(to_signed(-1024,SDLEN)),
    to_std_logic_vector(to_signed(-485,SDLEN)),
    to_std_logic_vector(to_signed(209,SDLEN)),
    to_std_logic_vector(to_signed(862,SDLEN)),
    to_std_logic_vector(to_signed(1280,SDLEN)),
    to_std_logic_vector(to_signed(-32313,SDLEN)),
    to_std_logic_vector(to_signed(-14461,SDLEN)),
    to_std_logic_vector(to_signed(-23925,SDLEN)),
    to_std_logic_vector(to_signed(-15334,SDLEN)),
    to_std_logic_vector(to_signed(15774,SDLEN))
  );

end G729A_CODEC_ST_ROM_PKG;

package body G729A_CODEC_ST_ROM_PKG is

  -- empty package body

end G729A_CODEC_ST_ROM_PKG;
