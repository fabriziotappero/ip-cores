

`define VENDOR_FPGA



