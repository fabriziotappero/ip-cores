--  Copyright (C) 2004-2005 Digish Pandya <digish.pandya@gmail.com>

--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.

-- VHDL Test Bench Created from source file tf_lms.vhd -- 14:23:32 02/24/2005
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends 
-- that these types always be used for the top-level I/O of a design in order 
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

LIBRARY ieee;
USE IEEE.STD_LOGIC_TEXTIO.ALL;
USE STD.TEXTIO.ALL;

ENTITY testbench IS
END testbench;

ARCHITECTURE behavior OF testbench IS 
    FILE RESULTS: TEXT IS OUT "yout.txt";
    FILE ERRF: TEXT IS OUT "error.txt";

    FUNCTION to_hex( x : IN std_logic_vector) RETURN string IS
    VARIABLE result  : STRING(1 TO 8); -- 1024 bits max
    VARIABLE i       : INTEGER;
    VARIABLE imod    : INTEGER;
    VARIABLE j       : INTEGER;
    VARIABLE newx    : std_logic_vector(1023 DOWNTO 0);
    BEGIN
      newx := (OTHERS => '0');
      newx(x'RANGE) := x;
      i := 7;
      j := 1;

      WHILE i >= 0 LOOP
        IF    newx(i) = '0' THEN result(j) := '0';
	   elsif newx(i) = '1' THEN result(j) := '1';
        ELSE result(j) := 'X';
        END IF;

        i := i-1;
	   j := j+1;
      END LOOP;
      RETURN result(1 TO j-1);
    END;

	COMPONENT tf_lms
	PORT(
		xin : IN std_logic_vector(7 downto 0);
		dxin : IN std_logic_vector(7 downto 0);
		clock : IN std_logic;
		err: out std_logic_vector(7 downto 0);
      	adapt_en: in std_logic;		 
		yout : OUT std_logic_vector(7 downto 0)
		);
	END COMPONENT;

	SIGNAL xin :  std_logic_vector(7 downto 0);
	SIGNAL dxin :  std_logic_vector(7 downto 0);
	SIGNAL clock :  std_logic;
	SIGNAL yout :  std_logic_vector(7 downto 0);
	signal err: std_logic_vector(7 downto 0);
	signal adapt_en : std_logic;
	CONSTANT clk_high   : time := 10 ns;
	CONSTANT clk_low    : time := 10 ns;
	CONSTANT clk_period : time := 20 ns;
	CONSTANT clk_hold   : time := 4 ns;



	  TYPE filter_data IS ARRAY (0 TO 999) OF std_logic_vector(7 downto 0);
	  TYPE filter_out_table IS ARRAY (0 TO 999)OF std_logic_vector(7 downto 0);

	  -- Constants
	  CONSTANT filter_dx_in : filter_data :=
	    (    	

"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000",
"01000000",
"11000000"
		
);
	  CONSTANT filter_x_in : filter_data :=
	    (

"11110011",
"00100110",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010",
"10100110",
"01011010"

);



BEGIN

	uut: tf_lms PORT MAP(
		xin => xin,
		dxin => dxin,
		clock => clock,
		err => err,
     	adapt_en => adapt_en,		 
		yout => yout
	);


-- *** Test Bench - User Defined Section ***
   clk_gen: PROCESS
   BEGIN
	    clock <= '1';
	    WAIT FOR clk_high;
	    clock <= '0';
	    WAIT FOR clk_low;

   END PROCESS clk_gen;

   tb:
   PROCESS
    		variable IN_x,IN_dx:std_logic_vector(7 downto 0); 
		VARIABLE TX_STR : String(1 to 512);
		VARIABLE TX_LOC : LINE;
		VARIABLE RX_LOC : LINE;

  
   BEGIN					    
				   
		adapt_en <= '1';

		FOR n IN 0 TO 500 LOOP
--			readline(F_XIN,xin);
			--xin <= IN_X;
			--Deallocate(RX_LOC);
			xin  <= filter_x_in(n);
	   		dxin <= filter_dx_in(n);
			wait for clk_period;
			write(TX_LOC,string'("'"));
			write(TX_LOC, yout);	
			write(TX_LOC,string'("'"));
			writeline(results, TX_LOC);
			Deallocate(TX_LOC);
			write(TX_LOC,string'("'"));
			write(TX_LOC, err);	
			write(TX_LOC,string'("'"));
			writeline(ERRF, TX_LOC);
			Deallocate(TX_LOC);
		end loop;

	--	adapt_en <= '0';

		FOR n IN 501 TO 999 LOOP
--			readline(F_XIN,xin);
			--xin <= IN_X;
			--Deallocate(RX_LOC);
			xin  <= filter_x_in(n);
	   		dxin <= filter_dx_in(n);
			wait for clk_period;
			write(TX_LOC,string'("'"));
			write(TX_LOC, yout);	
			write(TX_LOC,string'("'"));
			writeline(results, TX_LOC);
			Deallocate(TX_LOC);
			write(TX_LOC,string'("'"));
			write(TX_LOC, err);	
			write(TX_LOC,string'("'"));
			writeline(ERRF, TX_LOC);
			Deallocate(TX_LOC);
		end loop;

		
   wait; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
