// alu controller defines
// `define  addAB     00
// `define  subAB     01
// `define  incA      02
// `define  incB      03
// `define  decA      04
// `define  decB      05
// `define  cmpAB     06
// `define  andAB     07
// `define  orAB      08
// `define  xorAB     09
// `define  cplB      10
// `define  cplA      11
// `define  slAB      12
// `define  srAB      13
// `define  clrALL    14


`define  clrZ       0

`define  clrV       1
`define  clrC       2
       
`define  cADD_AB    0
`define  cINC_A     1
`define  cINC_B     9
`define  cSUB_AB    2
`define  cCMP_AB    3
`define  cASL_AbyB  4
`define  cASR_AbyB  5
`define  cCLR       6
`define  cDEC_A     7
`define  cDEC_B     8
`define  cMUL_AB   10
`define  cCPL_A    11
`define  cAND_AB   12
`define  cOR_AB    13
`define  cXOR_AB   14
`define  cCPL_B    15
