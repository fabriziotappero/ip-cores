---------------------------------------------------------------------
----                                                             ----
----  DCT IP core                                                ----
----                                                             ----
----  Authors: Anatoliy Sergienko, Volodya Lepeha                ----
----  Company: Unicore Systems http://unicore.co.ua              ----
----                                                             ----
----  Downloaded from: http://www.opencores.org                  ----
----                                                             ----
---------------------------------------------------------------------
----                                                             ----
---- Copyright (C) 2006-2010 Unicore Systems LTD                 ----
---- www.unicore.co.ua                                           ----
---- o.uzenkov@unicore.co.ua                                     ----
----                                                             ----
---- This source file may be used and distributed without        ----
---- restriction provided that this copyright statement is not   ----
---- removed from the file and that any derivative work contains ----
---- the original copyright notice and the associated disclaimer.----
----                                                             ----
---- THIS SOFTWARE IS PROVIDED "AS IS"                           ----
---- AND ANY EXPRESSED OR IMPLIED WARRANTIES,                    ----
---- INCLUDING, BUT NOT LIMITED TO, THE IMPLIED                  ----
---- WARRANTIES OF MERCHANTABILITY, NONINFRINGEMENT              ----
---- AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.        ----
---- IN NO EVENT SHALL THE UNICORE SYSTEMS OR ITS                ----
---- CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,            ----
---- INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL            ----
---- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT         ----
---- OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,               ----
---- DATA, OR PROFITS; OR BUSINESS INTERRUPTION)                 ----
---- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,              ----
---- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT              ----
---- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING                 ----
---- IN ANY WAY OUT OF THE USE OF THIS SOFTWARE,                 ----
---- EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.          ----
----                                                             ----
---------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.math_real.all;

entity BMP_GENERATOR is	 
	generic(  SIGNED_DATA : integer:= 0;   --  input data - 0 - unsigned, 1 - signed
		RANDOM:integer:=1 );
	port (
		CLK: in STD_LOGIC;
		RST: in STD_LOGIC;
		START: out STD_LOGIC;
		DATA: out STD_LOGIC_VECTOR (7 downto 0):=x"01"
		);
end BMP_GENERATOR;


architecture BMP_GENERATOR of BMP_GENERATOR is	   
	type TLUT is array(0 to 2047 ) of integer;	
	Constant ROMBMP:Tlut:=( ( 

	
	-- data patterns		
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	108,-25,-127,-72,72,127, 25,-109,
	
	127,127,127,127, 127,127,127,127,
	52,52,52,52,52,52,52,52,
	-52,-52,-52,-52,-52,-52,-52,-52,
	-127,-127,-127,-127,-127,-127,-127,-127,
	-127,-127,-127,-127,-127,-127,-127,-127,
	-52,-52,-52,-52,-52,-52,-52,-52,
	52,52,52,52,52,52,52,52,
	127,127,127,127, 127,127,127,127,
	
	
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,
	127,52,-52,-127,-127,-52,52, 127,  	
	
	
	
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52,   
	52,-127,127,-52,-52,127,-127,52, 
	
	
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	
	
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	127,-127,127,-127,127,-127,127,-127,
	
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	127,-117,90,-49,0,-49,90,117,
	
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	0,117,90,-49,-127,-49,90,117,
	
	
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90,
	127,-90, 0,90,-127,90,0,-90, 
	
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,
	127,-90,-90,127,-90,-90,127,-90,  
	
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	127,90,0,-90,-127,-90,0,90,
	
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,
	128,128,128,128, 128,128,128,128,	
	
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,
	127,127,127,127, 127,127,127,127,	   
	
	127,127,127,127,127,127,127,127,
	117,117,117,117,117,117,117,117,
	90,90,90,90, 90,90,90,90, 
	49,49,49,49,49,49,49,49,
	0,0,0,0,0,0,0,0,	
	49,49,49,49,49,49,49,49,
	90,90,90,90, 90,90,90,90, 
	117,117,117,117,117,117,117,117,
	
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,
	127, 117,	90, 49,00,49,90,117,   
	
	127,127,127,127,127,127,127,127,
	90,90,90,90, 90,90,90,90, 
	0,0,0,0,0,0,0,0,	   
	-90,-90,-90,-90, -90,-90,-90,-90,
	-127,-127,-127,-127,-127,-127,-127,-127,
	-90,-90,-90,-90, -90,-90,-90,-90,
	0,0,0,0,0,0,0,0,	   
	90,90,90,90, 90,90,90,90, 
	
	
	
	255, 255, 255, 255, 255, 255, 255, 255,  			
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255,   
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255,	  	
	--
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,
	0,255,0,255,0,255,0,255,			 
	
	
	
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127, 0,127,0,127,
	0,127,0,127,0,127,0,127,	 
	
	
	
	
	
	
	
	0,0,0,0,0,0,0,0,		 									  --3
	255,255,255,255,255,255,255,255,   		
	0,0,0,0,0,0,0,0,		 
	255,255,255,255,255,255,255,255,   		
	0,0,0,0,0,0,0,0,		 
	255,255,255,255,255,255,255,255,   		
	0,0,0,0,0,0,0,0,		 
	255,255,255,255,255,255,255,255,  
	
	
	255, 255, 255, 255, 255, 255, 255, 255,  			
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255, 
	255, 255, 255, 255, 255, 255, 255, 255,   	 
	0,0,0,0,0,0,0,0,		 								
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	
	
	183, 160, 94, 153, 194, 163, 132, 165, 	
	183, 153, 116, 176, 187, 166, 130, 169, 
	179, 168, 171, 182, 179, 165, 131, 167, 
	177, 177, 179, 177, 179, 165, 131, 167, 
	178, 178, 179, 176, 182, 164, 130, 171, 
	179, 180, 180, 179, 183, 169, 132, 169, 
	179, 179, 180, 182, 183, 170, 129, 172, 
	180, 179, 181, 179, 181, 170, 130, 169,    
	
	0,32,64,96,128, 160,192,224,	 	
	224,192,160,128,96, 64,32, 0,	
	0,32,64,96,128, 160,192,224,	 	
	224,192,160,128,96, 64,32, 0,
	0,32,64,96,128, 160,192,224,	 	
	224,192,160,128,96, 64,32, 0,
	0,32,64,96,128, 160,192,224,	 	
	224,192,160,128,96, 64,32, 0,
	
	128, 128, 128, 128, 128, 128, 128, 128, 
	128, 128, 128, 128, 128, 128, 128, 128,  
	128, 128, 192, 192, 192, 192, 128, 128, 
	128, 128, 192, 192, 192, 192, 128, 128,   
	128, 128, 192, 192, 192, 192, 128, 128, 
	128, 128, 192, 192, 192, 192, 128, 128, 
	128, 128, 128, 128, 128, 128, 128, 128, 
	128, 128, 128, 128, 128, 128, 128, 128, 
	
	90,100,110,120,130,140,150,160,	  
	91,101,111,121,131,141,151,161,			
	92,102,112,122,132,142,152,162,	  
	93,103,113,123,133,143,153,163,		
	90,100,110,120,130,140,150,160,	  
	91,101,111,121,131,141,151,161,			
	92,102,112,122,132,142,152,162,	  
	93,103,113,123,133,143,153,163,
	
	0,32,64,96,128, 160,192,224,	  
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	0,32,64,96,128, 160,192,224,
	
	183, 160, 94, 153, 194, 163, 132, 165, 	
	183, 153, 116, 176, 187, 166, 130, 169, 
	179, 168, 171, 182, 179, 165, 131, 167, 
	177, 177, 179, 177, 179, 165, 131, 167, 
	178, 178, 179, 176, 182, 164, 130, 171, 
	179, 180, 180, 179, 183, 169, 132, 169, 
	179, 179, 180, 182, 183, 170, 129, 173, 
	180, 179, 181, 179, 181, 170, 130, 169, 
	
	
	159, 128, 198, 128, 128, 128, 140, 128, 
	128, 128, 128, 128, 128, 128, 128, 128, 
	198, 128, 155, 128, 128, 128, 166, 128, 
	128, 128, 128, 128, 128, 128, 128, 128,   
	128, 128, 128, 128, 128, 128, 128, 128, 
	128, 128, 128, 128, 128, 128, 128, 128, 
	140, 128, 156, 128, 128, 128, 132, 128, 
	128, 128, 128, 128, 128, 128, 128, 128, 
	
	others=>127
	
	));	 			 
	
	signal dr,DATAi: STD_LOGIC_VECTOR (7 downto 0);
	signal 	index: integer range 0 to 2048; 					  
	
begin			
	
	process(clk)  --Generator of random images
		variable a,b:integer:=333;
		variable s:real;		 
		variable d,d1,d2,d3,d4,do:integer:=0;
	begin					
		if clk='1' then 
			UNIFORM(	a,b,s);	
			d4:=d3;
			d3:=d2;
			d2:=d1;				
			d1:=d;	  
			d:=integer(s*2.0**8);   
			--some LP filtering
			do :=(d +4*d1+ 6*d2+4*d3+d4)/16;
			dr<=conv_std_logic_vector(do,8)	;	 
		end if;  
		
	end process;
	
	
	DATA_OUTPUT:process(CLK,RST)
		
		variable delay: integer; 
		variable STARTi: STD_LOGIC;
		variable startdel:boolean;
	begin				
		if	 RST='1'  then
			startdel:=false;	
			STARTi:='0';
			delay:=0;
		elsif  CLK='1' and CLK'event and delay<10000 then 		 
			delay:=delay+1;
			if delay=10 or delay=11 then--or delay=500 or delay= 501  or delay=800 or delay= 801 then
				STARTi:='1' ;
			elsif delay=12  then --or delay= 502 or delay= 802 then		 
				STARTi:='0';
				startdel:=true;	  
			end if;
		end if;
		
		if RST='1'  then
			index<=0;
		elsif CLK='1' and CLK'event and startdel  then 
			if RANDOM=0 then   
				
				DATAi<=CONV_STD_LOGIC_VECTOR(INTEGER(ROMBMP(index)),8) after 7 ns;
				index<=(index+1) mod 2048;		 
			else
				DATAi<=dr;	
			end if;
		end if;			
		START<=STARTi after 5 ns;
		
	end process;
	
	DATA<= unsigned(DATAi)-UNSIGNED(X"80") when SIGNED_DATA=0 else DATAi; 
	
end BMP_GENERATOR;
