-- SDHC-SC-Core
-- Secure Digital High Capacity Self Configuring Core
-- 
-- (C) Copyright 2010, Rainer Kastl
-- All rights reserved.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the <organization> nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS  "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL <COPYRIGHT HOLDER> BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- File        : Counter-Rtl-a.vhdl
-- Owner       : Rainer Kastl
-- Description : Generic counter
-- Links       : 
-- 

architecture Rtl of Counter is

type aReg is record
	Counter : unsigned(gBitWidth - 1 downto 0);
	Enabled : std_ulogic;
end record aReg;

constant cDefaultReg : aReg := (
Counter => (others => '1'),
Enabled => cInactivated);

signal R : aReg := cDefaultReg;

begin

	Regs : process (iClk)
	begin
		if (iClk'event and iClk = cActivated) then
			if (iRstSync = cActivated) then
				R <= cDefaultReg;
			else
				oStrobe <= cInactivated;

				if (iDisable = cActivated) then
					R.Enabled <= cInactivated;
					R.Counter <= to_unsigned(0, R.Counter'length);

				elsif (iEnable = cActivated or R.Enabled = cActivated) then
					R.Enabled <= cActivated;

					if (R.Counter = iMax) then
						R.Counter <= to_unsigned(0, R.Counter'length);
						oStrobe   <= cActivated;
						R.Enabled <= cInactivated;

					else 
						R.Counter <= R.Counter + 1;
					end if;

				end if;
			end if;
		end if;
	end process Regs;

end architecture Rtl;
