@0
01
20
03
40
05
60
07
80
01
02
00
07
80
50
51
00
ff
ff
ff
ff
