--------------------------------------------------------------------------
-- Package of Direct Digital Synthesizer (DDS) sinewave generator components
--
-- NOTE: These components are for producing digital samples of sinewaves
--       by using sinewave lookup tables.  For modules which produce
--       single bit pulses of known frequency and/or duty cycle, please
--       refer to "dds_pack.vhd"
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package dds_sine_pack is

  component quadrature_oscillator
    generic(
      AMPL_BITS         : natural;
      AMPL_VALUE        : natural; -- Set to some value below full scale.  There is no saturation!
      SAMPLES_PER_CYCLE : natural
    );
    port(
      clk_i     : in  std_logic; -- System clock
      rst_n_i   : in  std_logic; -- Low asserted reset
      clk_en_i  : in  std_logic; -- clock enable, determines sample rate

      -- Sine and Cosine outputs
      sin_o     : out signed(AMPL_BITS-1 downto 0);
      cos_o     : out signed(AMPL_BITS-1 downto 0)
    );
  end component;

  component sine_generator_dds
    generic(
      PHI_BITS     : natural; -- Bits in phase accumulator, must be >= PHASE_BITS
      AMPL_BITS    : natural;
      PHASE_BITS   : natural
    );
    port(
      clk_i     : in  std_logic;
      rst_n_i   : in  std_logic;
      clk_en_i  : in  std_logic;

      -- Frequency Tuning Word input
      ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

      -- Outputs
      accum_o   : out unsigned(PHI_BITS-1 downto 0);
      sine_o    : out signed(AMPL_BITS-1 downto 0)
    );
  end component;

  component dds_sine
    generic(
      PHI_BITS     : natural; -- Bits in phase accumulator, must be >= PHASE_BITS
      AMPL_BITS    : natural;
      PHASE_BITS   : natural
    );
    port(
      clk_i     : in  std_logic;
      rst_n_i   : in  std_logic;
      clk_en_i  : in  std_logic;

      -- Look Up Table interface
      lut_adr_o : out unsigned(PHASE_BITS-3 downto 0); -- Quarter wave LUT
      lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

      -- Frequency Tuning Word input
      ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

      -- Outputs
      accum_o   : out unsigned(PHI_BITS-1 downto 0);
      sine_o    : out signed(AMPL_BITS-1 downto 0)
    );
  end component;

  component dds_sine_non_power_of_two
    generic(
      PHI_BITS     : natural; -- Bits in phase accumulator, must be >= PHASE_BITS
      AMPL_BITS    : natural;
      PHASE_LENGTH : natural;
      PHASE_BITS   : natural
    );
    port(
      clk_i     : in  std_logic;
      rst_n_i   : in  std_logic;
      clk_en_i  : in  std_logic;

      -- Look Up Table interface
      lut_adr_o : out unsigned(PHASE_BITS-3 downto 0); -- Quarter wave LUT
      lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

      -- Frequency Tuning Word input
      ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

      -- Outputs
      accum_o   : out unsigned(PHI_BITS-1 downto 0);
      sine_o    : out signed(AMPL_BITS-1 downto 0)
      );
  end component;

  component dds_arb
    generic(
      PHI_BITS     : natural; -- Bits in phase accumulator, must be >= PHASE_BITS
      AMPL_BITS    : natural;
      PHASE_BITS   : natural
    );
    port(
      clk_i     : in  std_logic;
      rst_n_i   : in  std_logic;
      clk_en_i  : in  std_logic;

      -- Look Up Table interface
      lut_adr_o : out unsigned(PHASE_BITS-1 downto 0); -- Full Wave LUT
      lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

      -- Frequency Tuning Word input
      ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

      -- Outputs
      accum_o   : out unsigned(PHI_BITS-1 downto 0);
      arb_o     : out signed(AMPL_BITS-1 downto 0)
    );
  end component;

-- Quarter sine lookup table
type lut_5000_x_16_type is array(0 to 1249) of unsigned(15 downto 0);
constant sine_lut_5000_x_16 : lut_5000_x_16_type := (
    to_unsigned(0,16),
    to_unsigned(41,16),
    to_unsigned(82,16),
    to_unsigned(124,16),
    to_unsigned(165,16),
    to_unsigned(206,16),
    to_unsigned(247,16),
    to_unsigned(288,16),
    to_unsigned(329,16),
    to_unsigned(371,16),
    to_unsigned(412,16),
    to_unsigned(453,16),
    to_unsigned(494,16),
    to_unsigned(535,16),
    to_unsigned(576,16),
    to_unsigned(618,16),
    to_unsigned(659,16),
    to_unsigned(700,16),
    to_unsigned(741,16),
    to_unsigned(782,16),
    to_unsigned(823,16),
    to_unsigned(865,16),
    to_unsigned(906,16),
    to_unsigned(947,16),
    to_unsigned(988,16),
    to_unsigned(1029,16),
    to_unsigned(1070,16),
    to_unsigned(1112,16),
    to_unsigned(1153,16),
    to_unsigned(1194,16),
    to_unsigned(1235,16),
    to_unsigned(1276,16),
    to_unsigned(1317,16),
    to_unsigned(1358,16),
    to_unsigned(1400,16),
    to_unsigned(1441,16),
    to_unsigned(1482,16),
    to_unsigned(1523,16),
    to_unsigned(1564,16),
    to_unsigned(1605,16),
    to_unsigned(1646,16),
    to_unsigned(1687,16),
    to_unsigned(1729,16),
    to_unsigned(1770,16),
    to_unsigned(1811,16),
    to_unsigned(1852,16),
    to_unsigned(1893,16),
    to_unsigned(1934,16),
    to_unsigned(1975,16),
    to_unsigned(2016,16),
    to_unsigned(2057,16),
    to_unsigned(2099,16),
    to_unsigned(2140,16),
    to_unsigned(2181,16),
    to_unsigned(2222,16),
    to_unsigned(2263,16),
    to_unsigned(2304,16),
    to_unsigned(2345,16),
    to_unsigned(2386,16),
    to_unsigned(2427,16),
    to_unsigned(2468,16),
    to_unsigned(2509,16),
    to_unsigned(2550,16),
    to_unsigned(2591,16),
    to_unsigned(2632,16),
    to_unsigned(2673,16),
    to_unsigned(2715,16),
    to_unsigned(2756,16),
    to_unsigned(2797,16),
    to_unsigned(2838,16),
    to_unsigned(2879,16),
    to_unsigned(2920,16),
    to_unsigned(2961,16),
    to_unsigned(3002,16),
    to_unsigned(3043,16),
    to_unsigned(3084,16),
    to_unsigned(3125,16),
    to_unsigned(3166,16),
    to_unsigned(3207,16),
    to_unsigned(3248,16),
    to_unsigned(3289,16),
    to_unsigned(3330,16),
    to_unsigned(3370,16),
    to_unsigned(3411,16),
    to_unsigned(3452,16),
    to_unsigned(3493,16),
    to_unsigned(3534,16),
    to_unsigned(3575,16),
    to_unsigned(3616,16),
    to_unsigned(3657,16),
    to_unsigned(3698,16),
    to_unsigned(3739,16),
    to_unsigned(3780,16),
    to_unsigned(3821,16),
    to_unsigned(3862,16),
    to_unsigned(3902,16),
    to_unsigned(3943,16),
    to_unsigned(3984,16),
    to_unsigned(4025,16),
    to_unsigned(4066,16),
    to_unsigned(4107,16),
    to_unsigned(4148,16),
    to_unsigned(4188,16),
    to_unsigned(4229,16),
    to_unsigned(4270,16),
    to_unsigned(4311,16),
    to_unsigned(4352,16),
    to_unsigned(4393,16),
    to_unsigned(4433,16),
    to_unsigned(4474,16),
    to_unsigned(4515,16),
    to_unsigned(4556,16),
    to_unsigned(4597,16),
    to_unsigned(4637,16),
    to_unsigned(4678,16),
    to_unsigned(4719,16),
    to_unsigned(4760,16),
    to_unsigned(4800,16),
    to_unsigned(4841,16),
    to_unsigned(4882,16),
    to_unsigned(4922,16),
    to_unsigned(4963,16),
    to_unsigned(5004,16),
    to_unsigned(5045,16),
    to_unsigned(5085,16),
    to_unsigned(5126,16),
    to_unsigned(5167,16),
    to_unsigned(5207,16),
    to_unsigned(5248,16),
    to_unsigned(5288,16),
    to_unsigned(5329,16),
    to_unsigned(5370,16),
    to_unsigned(5410,16),
    to_unsigned(5451,16),
    to_unsigned(5492,16),
    to_unsigned(5532,16),
    to_unsigned(5573,16),
    to_unsigned(5613,16),
    to_unsigned(5654,16),
    to_unsigned(5694,16),
    to_unsigned(5735,16),
    to_unsigned(5776,16),
    to_unsigned(5816,16),
    to_unsigned(5857,16),
    to_unsigned(5897,16),
    to_unsigned(5938,16),
    to_unsigned(5978,16),
    to_unsigned(6019,16),
    to_unsigned(6059,16),
    to_unsigned(6099,16),
    to_unsigned(6140,16),
    to_unsigned(6180,16),
    to_unsigned(6221,16),
    to_unsigned(6261,16),
    to_unsigned(6302,16),
    to_unsigned(6342,16),
    to_unsigned(6382,16),
    to_unsigned(6423,16),
    to_unsigned(6463,16),
    to_unsigned(6504,16),
    to_unsigned(6544,16),
    to_unsigned(6584,16),
    to_unsigned(6625,16),
    to_unsigned(6665,16),
    to_unsigned(6705,16),
    to_unsigned(6746,16),
    to_unsigned(6786,16),
    to_unsigned(6826,16),
    to_unsigned(6866,16),
    to_unsigned(6907,16),
    to_unsigned(6947,16),
    to_unsigned(6987,16),
    to_unsigned(7027,16),
    to_unsigned(7068,16),
    to_unsigned(7108,16),
    to_unsigned(7148,16),
    to_unsigned(7188,16),
    to_unsigned(7228,16),
    to_unsigned(7268,16),
    to_unsigned(7309,16),
    to_unsigned(7349,16),
    to_unsigned(7389,16),
    to_unsigned(7429,16),
    to_unsigned(7469,16),
    to_unsigned(7509,16),
    to_unsigned(7549,16),
    to_unsigned(7589,16),
    to_unsigned(7629,16),
    to_unsigned(7669,16),
    to_unsigned(7709,16),
    to_unsigned(7749,16),
    to_unsigned(7789,16),
    to_unsigned(7829,16),
    to_unsigned(7869,16),
    to_unsigned(7909,16),
    to_unsigned(7949,16),
    to_unsigned(7989,16),
    to_unsigned(8029,16),
    to_unsigned(8069,16),
    to_unsigned(8109,16),
    to_unsigned(8149,16),
    to_unsigned(8189,16),
    to_unsigned(8229,16),
    to_unsigned(8268,16),
    to_unsigned(8308,16),
    to_unsigned(8348,16),
    to_unsigned(8388,16),
    to_unsigned(8428,16),
    to_unsigned(8467,16),
    to_unsigned(8507,16),
    to_unsigned(8547,16),
    to_unsigned(8587,16),
    to_unsigned(8626,16),
    to_unsigned(8666,16),
    to_unsigned(8706,16),
    to_unsigned(8746,16),
    to_unsigned(8785,16),
    to_unsigned(8825,16),
    to_unsigned(8865,16),
    to_unsigned(8904,16),
    to_unsigned(8944,16),
    to_unsigned(8983,16),
    to_unsigned(9023,16),
    to_unsigned(9063,16),
    to_unsigned(9102,16),
    to_unsigned(9142,16),
    to_unsigned(9181,16),
    to_unsigned(9221,16),
    to_unsigned(9260,16),
    to_unsigned(9300,16),
    to_unsigned(9339,16),
    to_unsigned(9379,16),
    to_unsigned(9418,16),
    to_unsigned(9458,16),
    to_unsigned(9497,16),
    to_unsigned(9536,16),
    to_unsigned(9576,16),
    to_unsigned(9615,16),
    to_unsigned(9654,16),
    to_unsigned(9694,16),
    to_unsigned(9733,16),
    to_unsigned(9772,16),
    to_unsigned(9812,16),
    to_unsigned(9851,16),
    to_unsigned(9890,16),
    to_unsigned(9930,16),
    to_unsigned(9969,16),
    to_unsigned(10008,16),
    to_unsigned(10047,16),
    to_unsigned(10086,16),
    to_unsigned(10126,16),
    to_unsigned(10165,16),
    to_unsigned(10204,16),
    to_unsigned(10243,16),
    to_unsigned(10282,16),
    to_unsigned(10321,16),
    to_unsigned(10360,16),
    to_unsigned(10399,16),
    to_unsigned(10438,16),
    to_unsigned(10477,16),
    to_unsigned(10516,16),
    to_unsigned(10555,16),
    to_unsigned(10594,16),
    to_unsigned(10633,16),
    to_unsigned(10672,16),
    to_unsigned(10711,16),
    to_unsigned(10750,16),
    to_unsigned(10789,16),
    to_unsigned(10828,16),
    to_unsigned(10867,16),
    to_unsigned(10905,16),
    to_unsigned(10944,16),
    to_unsigned(10983,16),
    to_unsigned(11022,16),
    to_unsigned(11061,16),
    to_unsigned(11099,16),
    to_unsigned(11138,16),
    to_unsigned(11177,16),
    to_unsigned(11216,16),
    to_unsigned(11254,16),
    to_unsigned(11293,16),
    to_unsigned(11332,16),
    to_unsigned(11370,16),
    to_unsigned(11409,16),
    to_unsigned(11447,16),
    to_unsigned(11486,16),
    to_unsigned(11525,16),
    to_unsigned(11563,16),
    to_unsigned(11602,16),
    to_unsigned(11640,16),
    to_unsigned(11679,16),
    to_unsigned(11717,16),
    to_unsigned(11755,16),
    to_unsigned(11794,16),
    to_unsigned(11832,16),
    to_unsigned(11871,16),
    to_unsigned(11909,16),
    to_unsigned(11947,16),
    to_unsigned(11986,16),
    to_unsigned(12024,16),
    to_unsigned(12062,16),
    to_unsigned(12101,16),
    to_unsigned(12139,16),
    to_unsigned(12177,16),
    to_unsigned(12215,16),
    to_unsigned(12254,16),
    to_unsigned(12292,16),
    to_unsigned(12330,16),
    to_unsigned(12368,16),
    to_unsigned(12406,16),
    to_unsigned(12444,16),
    to_unsigned(12482,16),
    to_unsigned(12520,16),
    to_unsigned(12558,16),
    to_unsigned(12596,16),
    to_unsigned(12634,16),
    to_unsigned(12672,16),
    to_unsigned(12710,16),
    to_unsigned(12748,16),
    to_unsigned(12786,16),
    to_unsigned(12824,16),
    to_unsigned(12862,16),
    to_unsigned(12900,16),
    to_unsigned(12938,16),
    to_unsigned(12976,16),
    to_unsigned(13013,16),
    to_unsigned(13051,16),
    to_unsigned(13089,16),
    to_unsigned(13127,16),
    to_unsigned(13164,16),
    to_unsigned(13202,16),
    to_unsigned(13240,16),
    to_unsigned(13277,16),
    to_unsigned(13315,16),
    to_unsigned(13353,16),
    to_unsigned(13390,16),
    to_unsigned(13428,16),
    to_unsigned(13465,16),
    to_unsigned(13503,16),
    to_unsigned(13540,16),
    to_unsigned(13578,16),
    to_unsigned(13615,16),
    to_unsigned(13653,16),
    to_unsigned(13690,16),
    to_unsigned(13728,16),
    to_unsigned(13765,16),
    to_unsigned(13802,16),
    to_unsigned(13840,16),
    to_unsigned(13877,16),
    to_unsigned(13914,16),
    to_unsigned(13952,16),
    to_unsigned(13989,16),
    to_unsigned(14026,16),
    to_unsigned(14063,16),
    to_unsigned(14100,16),
    to_unsigned(14138,16),
    to_unsigned(14175,16),
    to_unsigned(14212,16),
    to_unsigned(14249,16),
    to_unsigned(14286,16),
    to_unsigned(14323,16),
    to_unsigned(14360,16),
    to_unsigned(14397,16),
    to_unsigned(14434,16),
    to_unsigned(14471,16),
    to_unsigned(14508,16),
    to_unsigned(14545,16),
    to_unsigned(14582,16),
    to_unsigned(14619,16),
    to_unsigned(14655,16),
    to_unsigned(14692,16),
    to_unsigned(14729,16),
    to_unsigned(14766,16),
    to_unsigned(14802,16),
    to_unsigned(14839,16),
    to_unsigned(14876,16),
    to_unsigned(14913,16),
    to_unsigned(14949,16),
    to_unsigned(14986,16),
    to_unsigned(15022,16),
    to_unsigned(15059,16),
    to_unsigned(15096,16),
    to_unsigned(15132,16),
    to_unsigned(15169,16),
    to_unsigned(15205,16),
    to_unsigned(15242,16),
    to_unsigned(15278,16),
    to_unsigned(15314,16),
    to_unsigned(15351,16),
    to_unsigned(15387,16),
    to_unsigned(15424,16),
    to_unsigned(15460,16),
    to_unsigned(15496,16),
    to_unsigned(15532,16),
    to_unsigned(15569,16),
    to_unsigned(15605,16),
    to_unsigned(15641,16),
    to_unsigned(15677,16),
    to_unsigned(15713,16),
    to_unsigned(15750,16),
    to_unsigned(15786,16),
    to_unsigned(15822,16),
    to_unsigned(15858,16),
    to_unsigned(15894,16),
    to_unsigned(15930,16),
    to_unsigned(15966,16),
    to_unsigned(16002,16),
    to_unsigned(16038,16),
    to_unsigned(16073,16),
    to_unsigned(16109,16),
    to_unsigned(16145,16),
    to_unsigned(16181,16),
    to_unsigned(16217,16),
    to_unsigned(16253,16),
    to_unsigned(16288,16),
    to_unsigned(16324,16),
    to_unsigned(16360,16),
    to_unsigned(16395,16),
    to_unsigned(16431,16),
    to_unsigned(16467,16),
    to_unsigned(16502,16),
    to_unsigned(16538,16),
    to_unsigned(16573,16),
    to_unsigned(16609,16),
    to_unsigned(16644,16),
    to_unsigned(16680,16),
    to_unsigned(16715,16),
    to_unsigned(16751,16),
    to_unsigned(16786,16),
    to_unsigned(16821,16),
    to_unsigned(16857,16),
    to_unsigned(16892,16),
    to_unsigned(16927,16),
    to_unsigned(16962,16),
    to_unsigned(16998,16),
    to_unsigned(17033,16),
    to_unsigned(17068,16),
    to_unsigned(17103,16),
    to_unsigned(17138,16),
    to_unsigned(17173,16),
    to_unsigned(17208,16),
    to_unsigned(17243,16),
    to_unsigned(17278,16),
    to_unsigned(17313,16),
    to_unsigned(17348,16),
    to_unsigned(17383,16),
    to_unsigned(17418,16),
    to_unsigned(17453,16),
    to_unsigned(17488,16),
    to_unsigned(17523,16),
    to_unsigned(17557,16),
    to_unsigned(17592,16),
    to_unsigned(17627,16),
    to_unsigned(17662,16),
    to_unsigned(17696,16),
    to_unsigned(17731,16),
    to_unsigned(17766,16),
    to_unsigned(17800,16),
    to_unsigned(17835,16),
    to_unsigned(17869,16),
    to_unsigned(17904,16),
    to_unsigned(17938,16),
    to_unsigned(17973,16),
    to_unsigned(18007,16),
    to_unsigned(18041,16),
    to_unsigned(18076,16),
    to_unsigned(18110,16),
    to_unsigned(18144,16),
    to_unsigned(18179,16),
    to_unsigned(18213,16),
    to_unsigned(18247,16),
    to_unsigned(18281,16),
    to_unsigned(18315,16),
    to_unsigned(18350,16),
    to_unsigned(18384,16),
    to_unsigned(18418,16),
    to_unsigned(18452,16),
    to_unsigned(18486,16),
    to_unsigned(18520,16),
    to_unsigned(18554,16),
    to_unsigned(18588,16),
    to_unsigned(18622,16),
    to_unsigned(18655,16),
    to_unsigned(18689,16),
    to_unsigned(18723,16),
    to_unsigned(18757,16),
    to_unsigned(18791,16),
    to_unsigned(18824,16),
    to_unsigned(18858,16),
    to_unsigned(18892,16),
    to_unsigned(18925,16),
    to_unsigned(18959,16),
    to_unsigned(18992,16),
    to_unsigned(19026,16),
    to_unsigned(19060,16),
    to_unsigned(19093,16),
    to_unsigned(19126,16),
    to_unsigned(19160,16),
    to_unsigned(19193,16),
    to_unsigned(19227,16),
    to_unsigned(19260,16),
    to_unsigned(19293,16),
    to_unsigned(19327,16),
    to_unsigned(19360,16),
    to_unsigned(19393,16),
    to_unsigned(19426,16),
    to_unsigned(19459,16),
    to_unsigned(19492,16),
    to_unsigned(19525,16),
    to_unsigned(19559,16),
    to_unsigned(19592,16),
    to_unsigned(19625,16),
    to_unsigned(19658,16),
    to_unsigned(19690,16),
    to_unsigned(19723,16),
    to_unsigned(19756,16),
    to_unsigned(19789,16),
    to_unsigned(19822,16),
    to_unsigned(19855,16),
    to_unsigned(19887,16),
    to_unsigned(19920,16),
    to_unsigned(19953,16),
    to_unsigned(19985,16),
    to_unsigned(20018,16),
    to_unsigned(20051,16),
    to_unsigned(20083,16),
    to_unsigned(20116,16),
    to_unsigned(20148,16),
    to_unsigned(20181,16),
    to_unsigned(20213,16),
    to_unsigned(20245,16),
    to_unsigned(20278,16),
    to_unsigned(20310,16),
    to_unsigned(20342,16),
    to_unsigned(20375,16),
    to_unsigned(20407,16),
    to_unsigned(20439,16),
    to_unsigned(20471,16),
    to_unsigned(20503,16),
    to_unsigned(20535,16),
    to_unsigned(20568,16),
    to_unsigned(20600,16),
    to_unsigned(20632,16),
    to_unsigned(20664,16),
    to_unsigned(20696,16),
    to_unsigned(20727,16),
    to_unsigned(20759,16),
    to_unsigned(20791,16),
    to_unsigned(20823,16),
    to_unsigned(20855,16),
    to_unsigned(20886,16),
    to_unsigned(20918,16),
    to_unsigned(20950,16),
    to_unsigned(20982,16),
    to_unsigned(21013,16),
    to_unsigned(21045,16),
    to_unsigned(21076,16),
    to_unsigned(21108,16),
    to_unsigned(21139,16),
    to_unsigned(21171,16),
    to_unsigned(21202,16),
    to_unsigned(21233,16),
    to_unsigned(21265,16),
    to_unsigned(21296,16),
    to_unsigned(21327,16),
    to_unsigned(21359,16),
    to_unsigned(21390,16),
    to_unsigned(21421,16),
    to_unsigned(21452,16),
    to_unsigned(21483,16),
    to_unsigned(21514,16),
    to_unsigned(21545,16),
    to_unsigned(21576,16),
    to_unsigned(21607,16),
    to_unsigned(21638,16),
    to_unsigned(21669,16),
    to_unsigned(21700,16),
    to_unsigned(21731,16),
    to_unsigned(21762,16),
    to_unsigned(21792,16),
    to_unsigned(21823,16),
    to_unsigned(21854,16),
    to_unsigned(21885,16),
    to_unsigned(21915,16),
    to_unsigned(21946,16),
    to_unsigned(21976,16),
    to_unsigned(22007,16),
    to_unsigned(22037,16),
    to_unsigned(22068,16),
    to_unsigned(22098,16),
    to_unsigned(22129,16),
    to_unsigned(22159,16),
    to_unsigned(22189,16),
    to_unsigned(22220,16),
    to_unsigned(22250,16),
    to_unsigned(22280,16),
    to_unsigned(22310,16),
    to_unsigned(22340,16),
    to_unsigned(22370,16),
    to_unsigned(22401,16),
    to_unsigned(22431,16),
    to_unsigned(22461,16),
    to_unsigned(22491,16),
    to_unsigned(22520,16),
    to_unsigned(22550,16),
    to_unsigned(22580,16),
    to_unsigned(22610,16),
    to_unsigned(22640,16),
    to_unsigned(22670,16),
    to_unsigned(22699,16),
    to_unsigned(22729,16),
    to_unsigned(22759,16),
    to_unsigned(22788,16),
    to_unsigned(22818,16),
    to_unsigned(22847,16),
    to_unsigned(22877,16),
    to_unsigned(22906,16),
    to_unsigned(22936,16),
    to_unsigned(22965,16),
    to_unsigned(22994,16),
    to_unsigned(23024,16),
    to_unsigned(23053,16),
    to_unsigned(23082,16),
    to_unsigned(23111,16),
    to_unsigned(23141,16),
    to_unsigned(23170,16),
    to_unsigned(23199,16),
    to_unsigned(23228,16),
    to_unsigned(23257,16),
    to_unsigned(23286,16),
    to_unsigned(23315,16),
    to_unsigned(23344,16),
    to_unsigned(23373,16),
    to_unsigned(23402,16),
    to_unsigned(23430,16),
    to_unsigned(23459,16),
    to_unsigned(23488,16),
    to_unsigned(23517,16),
    to_unsigned(23545,16),
    to_unsigned(23574,16),
    to_unsigned(23602,16),
    to_unsigned(23631,16),
    to_unsigned(23659,16),
    to_unsigned(23688,16),
    to_unsigned(23716,16),
    to_unsigned(23745,16),
    to_unsigned(23773,16),
    to_unsigned(23801,16),
    to_unsigned(23830,16),
    to_unsigned(23858,16),
    to_unsigned(23886,16),
    to_unsigned(23914,16),
    to_unsigned(23942,16),
    to_unsigned(23971,16),
    to_unsigned(23999,16),
    to_unsigned(24027,16),
    to_unsigned(24055,16),
    to_unsigned(24082,16),
    to_unsigned(24110,16),
    to_unsigned(24138,16),
    to_unsigned(24166,16),
    to_unsigned(24194,16),
    to_unsigned(24222,16),
    to_unsigned(24249,16),
    to_unsigned(24277,16),
    to_unsigned(24305,16),
    to_unsigned(24332,16),
    to_unsigned(24360,16),
    to_unsigned(24387,16),
    to_unsigned(24415,16),
    to_unsigned(24442,16),
    to_unsigned(24470,16),
    to_unsigned(24497,16),
    to_unsigned(24524,16),
    to_unsigned(24552,16),
    to_unsigned(24579,16),
    to_unsigned(24606,16),
    to_unsigned(24633,16),
    to_unsigned(24660,16),
    to_unsigned(24687,16),
    to_unsigned(24715,16),
    to_unsigned(24742,16),
    to_unsigned(24769,16),
    to_unsigned(24795,16),
    to_unsigned(24822,16),
    to_unsigned(24849,16),
    to_unsigned(24876,16),
    to_unsigned(24903,16),
    to_unsigned(24930,16),
    to_unsigned(24956,16),
    to_unsigned(24983,16),
    to_unsigned(25010,16),
    to_unsigned(25036,16),
    to_unsigned(25063,16),
    to_unsigned(25089,16),
    to_unsigned(25116,16),
    to_unsigned(25142,16),
    to_unsigned(25168,16),
    to_unsigned(25195,16),
    to_unsigned(25221,16),
    to_unsigned(25247,16),
    to_unsigned(25274,16),
    to_unsigned(25300,16),
    to_unsigned(25326,16),
    to_unsigned(25352,16),
    to_unsigned(25378,16),
    to_unsigned(25404,16),
    to_unsigned(25430,16),
    to_unsigned(25456,16),
    to_unsigned(25482,16),
    to_unsigned(25508,16),
    to_unsigned(25534,16),
    to_unsigned(25559,16),
    to_unsigned(25585,16),
    to_unsigned(25611,16),
    to_unsigned(25637,16),
    to_unsigned(25662,16),
    to_unsigned(25688,16),
    to_unsigned(25713,16),
    to_unsigned(25739,16),
    to_unsigned(25764,16),
    to_unsigned(25790,16),
    to_unsigned(25815,16),
    to_unsigned(25840,16),
    to_unsigned(25866,16),
    to_unsigned(25891,16),
    to_unsigned(25916,16),
    to_unsigned(25941,16),
    to_unsigned(25967,16),
    to_unsigned(25992,16),
    to_unsigned(26017,16),
    to_unsigned(26042,16),
    to_unsigned(26067,16),
    to_unsigned(26092,16),
    to_unsigned(26116,16),
    to_unsigned(26141,16),
    to_unsigned(26166,16),
    to_unsigned(26191,16),
    to_unsigned(26216,16),
    to_unsigned(26240,16),
    to_unsigned(26265,16),
    to_unsigned(26290,16),
    to_unsigned(26314,16),
    to_unsigned(26339,16),
    to_unsigned(26363,16),
    to_unsigned(26388,16),
    to_unsigned(26412,16),
    to_unsigned(26436,16),
    to_unsigned(26461,16),
    to_unsigned(26485,16),
    to_unsigned(26509,16),
    to_unsigned(26533,16),
    to_unsigned(26557,16),
    to_unsigned(26581,16),
    to_unsigned(26606,16),
    to_unsigned(26630,16),
    to_unsigned(26654,16),
    to_unsigned(26677,16),
    to_unsigned(26701,16),
    to_unsigned(26725,16),
    to_unsigned(26749,16),
    to_unsigned(26773,16),
    to_unsigned(26796,16),
    to_unsigned(26820,16),
    to_unsigned(26844,16),
    to_unsigned(26867,16),
    to_unsigned(26891,16),
    to_unsigned(26914,16),
    to_unsigned(26938,16),
    to_unsigned(26961,16),
    to_unsigned(26985,16),
    to_unsigned(27008,16),
    to_unsigned(27031,16),
    to_unsigned(27055,16),
    to_unsigned(27078,16),
    to_unsigned(27101,16),
    to_unsigned(27124,16),
    to_unsigned(27147,16),
    to_unsigned(27170,16),
    to_unsigned(27193,16),
    to_unsigned(27216,16),
    to_unsigned(27239,16),
    to_unsigned(27262,16),
    to_unsigned(27285,16),
    to_unsigned(27308,16),
    to_unsigned(27330,16),
    to_unsigned(27353,16),
    to_unsigned(27376,16),
    to_unsigned(27398,16),
    to_unsigned(27421,16),
    to_unsigned(27443,16),
    to_unsigned(27466,16),
    to_unsigned(27488,16),
    to_unsigned(27511,16),
    to_unsigned(27533,16),
    to_unsigned(27555,16),
    to_unsigned(27577,16),
    to_unsigned(27600,16),
    to_unsigned(27622,16),
    to_unsigned(27644,16),
    to_unsigned(27666,16),
    to_unsigned(27688,16),
    to_unsigned(27710,16),
    to_unsigned(27732,16),
    to_unsigned(27754,16),
    to_unsigned(27776,16),
    to_unsigned(27798,16),
    to_unsigned(27819,16),
    to_unsigned(27841,16),
    to_unsigned(27863,16),
    to_unsigned(27885,16),
    to_unsigned(27906,16),
    to_unsigned(27928,16),
    to_unsigned(27949,16),
    to_unsigned(27971,16),
    to_unsigned(27992,16),
    to_unsigned(28013,16),
    to_unsigned(28035,16),
    to_unsigned(28056,16),
    to_unsigned(28077,16),
    to_unsigned(28099,16),
    to_unsigned(28120,16),
    to_unsigned(28141,16),
    to_unsigned(28162,16),
    to_unsigned(28183,16),
    to_unsigned(28204,16),
    to_unsigned(28225,16),
    to_unsigned(28246,16),
    to_unsigned(28267,16),
    to_unsigned(28287,16),
    to_unsigned(28308,16),
    to_unsigned(28329,16),
    to_unsigned(28350,16),
    to_unsigned(28370,16),
    to_unsigned(28391,16),
    to_unsigned(28411,16),
    to_unsigned(28432,16),
    to_unsigned(28452,16),
    to_unsigned(28473,16),
    to_unsigned(28493,16),
    to_unsigned(28513,16),
    to_unsigned(28534,16),
    to_unsigned(28554,16),
    to_unsigned(28574,16),
    to_unsigned(28594,16),
    to_unsigned(28614,16),
    to_unsigned(28634,16),
    to_unsigned(28654,16),
    to_unsigned(28674,16),
    to_unsigned(28694,16),
    to_unsigned(28714,16),
    to_unsigned(28734,16),
    to_unsigned(28754,16),
    to_unsigned(28773,16),
    to_unsigned(28793,16),
    to_unsigned(28813,16),
    to_unsigned(28832,16),
    to_unsigned(28852,16),
    to_unsigned(28871,16),
    to_unsigned(28891,16),
    to_unsigned(28910,16),
    to_unsigned(28929,16),
    to_unsigned(28949,16),
    to_unsigned(28968,16),
    to_unsigned(28987,16),
    to_unsigned(29006,16),
    to_unsigned(29026,16),
    to_unsigned(29045,16),
    to_unsigned(29064,16),
    to_unsigned(29083,16),
    to_unsigned(29102,16),
    to_unsigned(29120,16),
    to_unsigned(29139,16),
    to_unsigned(29158,16),
    to_unsigned(29177,16),
    to_unsigned(29196,16),
    to_unsigned(29214,16),
    to_unsigned(29233,16),
    to_unsigned(29251,16),
    to_unsigned(29270,16),
    to_unsigned(29289,16),
    to_unsigned(29307,16),
    to_unsigned(29325,16),
    to_unsigned(29344,16),
    to_unsigned(29362,16),
    to_unsigned(29380,16),
    to_unsigned(29398,16),
    to_unsigned(29417,16),
    to_unsigned(29435,16),
    to_unsigned(29453,16),
    to_unsigned(29471,16),
    to_unsigned(29489,16),
    to_unsigned(29507,16),
    to_unsigned(29525,16),
    to_unsigned(29542,16),
    to_unsigned(29560,16),
    to_unsigned(29578,16),
    to_unsigned(29596,16),
    to_unsigned(29613,16),
    to_unsigned(29631,16),
    to_unsigned(29648,16),
    to_unsigned(29666,16),
    to_unsigned(29683,16),
    to_unsigned(29701,16),
    to_unsigned(29718,16),
    to_unsigned(29736,16),
    to_unsigned(29753,16),
    to_unsigned(29770,16),
    to_unsigned(29787,16),
    to_unsigned(29804,16),
    to_unsigned(29821,16),
    to_unsigned(29838,16),
    to_unsigned(29855,16),
    to_unsigned(29872,16),
    to_unsigned(29889,16),
    to_unsigned(29906,16),
    to_unsigned(29923,16),
    to_unsigned(29940,16),
    to_unsigned(29956,16),
    to_unsigned(29973,16),
    to_unsigned(29990,16),
    to_unsigned(30006,16),
    to_unsigned(30023,16),
    to_unsigned(30039,16),
    to_unsigned(30056,16),
    to_unsigned(30072,16),
    to_unsigned(30088,16),
    to_unsigned(30105,16),
    to_unsigned(30121,16),
    to_unsigned(30137,16),
    to_unsigned(30153,16),
    to_unsigned(30169,16),
    to_unsigned(30185,16),
    to_unsigned(30201,16),
    to_unsigned(30217,16),
    to_unsigned(30233,16),
    to_unsigned(30249,16),
    to_unsigned(30265,16),
    to_unsigned(30281,16),
    to_unsigned(30296,16),
    to_unsigned(30312,16),
    to_unsigned(30328,16),
    to_unsigned(30343,16),
    to_unsigned(30359,16),
    to_unsigned(30374,16),
    to_unsigned(30390,16),
    to_unsigned(30405,16),
    to_unsigned(30420,16),
    to_unsigned(30436,16),
    to_unsigned(30451,16),
    to_unsigned(30466,16),
    to_unsigned(30481,16),
    to_unsigned(30496,16),
    to_unsigned(30511,16),
    to_unsigned(30526,16),
    to_unsigned(30541,16),
    to_unsigned(30556,16),
    to_unsigned(30571,16),
    to_unsigned(30586,16),
    to_unsigned(30600,16),
    to_unsigned(30615,16),
    to_unsigned(30630,16),
    to_unsigned(30644,16),
    to_unsigned(30659,16),
    to_unsigned(30673,16),
    to_unsigned(30688,16),
    to_unsigned(30702,16),
    to_unsigned(30717,16),
    to_unsigned(30731,16),
    to_unsigned(30745,16),
    to_unsigned(30759,16),
    to_unsigned(30774,16),
    to_unsigned(30788,16),
    to_unsigned(30802,16),
    to_unsigned(30816,16),
    to_unsigned(30830,16),
    to_unsigned(30844,16),
    to_unsigned(30858,16),
    to_unsigned(30871,16),
    to_unsigned(30885,16),
    to_unsigned(30899,16),
    to_unsigned(30913,16),
    to_unsigned(30926,16),
    to_unsigned(30940,16),
    to_unsigned(30953,16),
    to_unsigned(30967,16),
    to_unsigned(30980,16),
    to_unsigned(30994,16),
    to_unsigned(31007,16),
    to_unsigned(31020,16),
    to_unsigned(31034,16),
    to_unsigned(31047,16),
    to_unsigned(31060,16),
    to_unsigned(31073,16),
    to_unsigned(31086,16),
    to_unsigned(31099,16),
    to_unsigned(31112,16),
    to_unsigned(31125,16),
    to_unsigned(31138,16),
    to_unsigned(31151,16),
    to_unsigned(31163,16),
    to_unsigned(31176,16),
    to_unsigned(31189,16),
    to_unsigned(31201,16),
    to_unsigned(31214,16),
    to_unsigned(31226,16),
    to_unsigned(31239,16),
    to_unsigned(31251,16),
    to_unsigned(31263,16),
    to_unsigned(31276,16),
    to_unsigned(31288,16),
    to_unsigned(31300,16),
    to_unsigned(31312,16),
    to_unsigned(31325,16),
    to_unsigned(31337,16),
    to_unsigned(31349,16),
    to_unsigned(31361,16),
    to_unsigned(31372,16),
    to_unsigned(31384,16),
    to_unsigned(31396,16),
    to_unsigned(31408,16),
    to_unsigned(31420,16),
    to_unsigned(31431,16),
    to_unsigned(31443,16),
    to_unsigned(31454,16),
    to_unsigned(31466,16),
    to_unsigned(31477,16),
    to_unsigned(31489,16),
    to_unsigned(31500,16),
    to_unsigned(31511,16),
    to_unsigned(31523,16),
    to_unsigned(31534,16),
    to_unsigned(31545,16),
    to_unsigned(31556,16),
    to_unsigned(31567,16),
    to_unsigned(31578,16),
    to_unsigned(31589,16),
    to_unsigned(31600,16),
    to_unsigned(31611,16),
    to_unsigned(31622,16),
    to_unsigned(31633,16),
    to_unsigned(31643,16),
    to_unsigned(31654,16),
    to_unsigned(31665,16),
    to_unsigned(31675,16),
    to_unsigned(31686,16),
    to_unsigned(31696,16),
    to_unsigned(31707,16),
    to_unsigned(31717,16),
    to_unsigned(31727,16),
    to_unsigned(31738,16),
    to_unsigned(31748,16),
    to_unsigned(31758,16),
    to_unsigned(31768,16),
    to_unsigned(31778,16),
    to_unsigned(31788,16),
    to_unsigned(31798,16),
    to_unsigned(31808,16),
    to_unsigned(31818,16),
    to_unsigned(31828,16),
    to_unsigned(31837,16),
    to_unsigned(31847,16),
    to_unsigned(31857,16),
    to_unsigned(31866,16),
    to_unsigned(31876,16),
    to_unsigned(31886,16),
    to_unsigned(31895,16),
    to_unsigned(31904,16),
    to_unsigned(31914,16),
    to_unsigned(31923,16),
    to_unsigned(31932,16),
    to_unsigned(31942,16),
    to_unsigned(31951,16),
    to_unsigned(31960,16),
    to_unsigned(31969,16),
    to_unsigned(31978,16),
    to_unsigned(31987,16),
    to_unsigned(31996,16),
    to_unsigned(32005,16),
    to_unsigned(32013,16),
    to_unsigned(32022,16),
    to_unsigned(32031,16),
    to_unsigned(32040,16),
    to_unsigned(32048,16),
    to_unsigned(32057,16),
    to_unsigned(32065,16),
    to_unsigned(32074,16),
    to_unsigned(32082,16),
    to_unsigned(32090,16),
    to_unsigned(32099,16),
    to_unsigned(32107,16),
    to_unsigned(32115,16),
    to_unsigned(32123,16),
    to_unsigned(32131,16),
    to_unsigned(32139,16),
    to_unsigned(32147,16),
    to_unsigned(32155,16),
    to_unsigned(32163,16),
    to_unsigned(32171,16),
    to_unsigned(32179,16),
    to_unsigned(32187,16),
    to_unsigned(32194,16),
    to_unsigned(32202,16),
    to_unsigned(32210,16),
    to_unsigned(32217,16),
    to_unsigned(32225,16),
    to_unsigned(32232,16),
    to_unsigned(32239,16),
    to_unsigned(32247,16),
    to_unsigned(32254,16),
    to_unsigned(32261,16),
    to_unsigned(32268,16),
    to_unsigned(32276,16),
    to_unsigned(32283,16),
    to_unsigned(32290,16),
    to_unsigned(32297,16),
    to_unsigned(32304,16),
    to_unsigned(32310,16),
    to_unsigned(32317,16),
    to_unsigned(32324,16),
    to_unsigned(32331,16),
    to_unsigned(32337,16),
    to_unsigned(32344,16),
    to_unsigned(32351,16),
    to_unsigned(32357,16),
    to_unsigned(32364,16),
    to_unsigned(32370,16),
    to_unsigned(32376,16),
    to_unsigned(32383,16),
    to_unsigned(32389,16),
    to_unsigned(32395,16),
    to_unsigned(32401,16),
    to_unsigned(32407,16),
    to_unsigned(32413,16),
    to_unsigned(32419,16),
    to_unsigned(32425,16),
    to_unsigned(32431,16),
    to_unsigned(32437,16),
    to_unsigned(32443,16),
    to_unsigned(32449,16),
    to_unsigned(32454,16),
    to_unsigned(32460,16),
    to_unsigned(32466,16),
    to_unsigned(32471,16),
    to_unsigned(32477,16),
    to_unsigned(32482,16),
    to_unsigned(32488,16),
    to_unsigned(32493,16),
    to_unsigned(32498,16),
    to_unsigned(32503,16),
    to_unsigned(32509,16),
    to_unsigned(32514,16),
    to_unsigned(32519,16),
    to_unsigned(32524,16),
    to_unsigned(32529,16),
    to_unsigned(32534,16),
    to_unsigned(32539,16),
    to_unsigned(32543,16),
    to_unsigned(32548,16),
    to_unsigned(32553,16),
    to_unsigned(32558,16),
    to_unsigned(32562,16),
    to_unsigned(32567,16),
    to_unsigned(32571,16),
    to_unsigned(32576,16),
    to_unsigned(32580,16),
    to_unsigned(32585,16),
    to_unsigned(32589,16),
    to_unsigned(32593,16),
    to_unsigned(32597,16),
    to_unsigned(32602,16),
    to_unsigned(32606,16),
    to_unsigned(32610,16),
    to_unsigned(32614,16),
    to_unsigned(32618,16),
    to_unsigned(32622,16),
    to_unsigned(32625,16),
    to_unsigned(32629,16),
    to_unsigned(32633,16),
    to_unsigned(32637,16),
    to_unsigned(32640,16),
    to_unsigned(32644,16),
    to_unsigned(32647,16),
    to_unsigned(32651,16),
    to_unsigned(32654,16),
    to_unsigned(32658,16),
    to_unsigned(32661,16),
    to_unsigned(32664,16),
    to_unsigned(32668,16),
    to_unsigned(32671,16),
    to_unsigned(32674,16),
    to_unsigned(32677,16),
    to_unsigned(32680,16),
    to_unsigned(32683,16),
    to_unsigned(32686,16),
    to_unsigned(32689,16),
    to_unsigned(32692,16),
    to_unsigned(32694,16),
    to_unsigned(32697,16),
    to_unsigned(32700,16),
    to_unsigned(32702,16),
    to_unsigned(32705,16),
    to_unsigned(32707,16),
    to_unsigned(32710,16),
    to_unsigned(32712,16),
    to_unsigned(32715,16),
    to_unsigned(32717,16),
    to_unsigned(32719,16),
    to_unsigned(32721,16),
    to_unsigned(32724,16),
    to_unsigned(32726,16),
    to_unsigned(32728,16),
    to_unsigned(32730,16),
    to_unsigned(32732,16),
    to_unsigned(32733,16),
    to_unsigned(32735,16),
    to_unsigned(32737,16),
    to_unsigned(32739,16),
    to_unsigned(32741,16),
    to_unsigned(32742,16),
    to_unsigned(32744,16),
    to_unsigned(32745,16),
    to_unsigned(32747,16),
    to_unsigned(32748,16),
    to_unsigned(32750,16),
    to_unsigned(32751,16),
    to_unsigned(32752,16),
    to_unsigned(32753,16),
    to_unsigned(32754,16),
    to_unsigned(32756,16),
    to_unsigned(32757,16),
    to_unsigned(32758,16),
    to_unsigned(32759,16),
    to_unsigned(32760,16),
    to_unsigned(32760,16),
    to_unsigned(32761,16),
    to_unsigned(32762,16),
    to_unsigned(32763,16),
    to_unsigned(32763,16),
    to_unsigned(32764,16),
    to_unsigned(32764,16),
    to_unsigned(32765,16),
    to_unsigned(32765,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16)
	);

-- Quarter sine lookup table
type lut_10000_type is array(0 to 2499) of unsigned(15 downto 0);
constant sine_lut_10000_x_16 : lut_10000_type := (
    to_unsigned(0,16),
    to_unsigned(21,16),
    to_unsigned(41,16),
    to_unsigned(62,16),
    to_unsigned(82,16),
    to_unsigned(103,16),
    to_unsigned(124,16),
    to_unsigned(144,16),
    to_unsigned(165,16),
    to_unsigned(185,16),
    to_unsigned(206,16),
    to_unsigned(226,16),
    to_unsigned(247,16),
    to_unsigned(268,16),
    to_unsigned(288,16),
    to_unsigned(309,16),
    to_unsigned(329,16),
    to_unsigned(350,16),
    to_unsigned(371,16),
    to_unsigned(391,16),
    to_unsigned(412,16),
    to_unsigned(432,16),
    to_unsigned(453,16),
    to_unsigned(474,16),
    to_unsigned(494,16),
    to_unsigned(515,16),
    to_unsigned(535,16),
    to_unsigned(556,16),
    to_unsigned(576,16),
    to_unsigned(597,16),
    to_unsigned(618,16),
    to_unsigned(638,16),
    to_unsigned(659,16),
    to_unsigned(679,16),
    to_unsigned(700,16),
    to_unsigned(721,16),
    to_unsigned(741,16),
    to_unsigned(762,16),
    to_unsigned(782,16),
    to_unsigned(803,16),
    to_unsigned(823,16),
    to_unsigned(844,16),
    to_unsigned(865,16),
    to_unsigned(885,16),
    to_unsigned(906,16),
    to_unsigned(926,16),
    to_unsigned(947,16),
    to_unsigned(968,16),
    to_unsigned(988,16),
    to_unsigned(1009,16),
    to_unsigned(1029,16),
    to_unsigned(1050,16),
    to_unsigned(1070,16),
    to_unsigned(1091,16),
    to_unsigned(1112,16),
    to_unsigned(1132,16),
    to_unsigned(1153,16),
    to_unsigned(1173,16),
    to_unsigned(1194,16),
    to_unsigned(1214,16),
    to_unsigned(1235,16),
    to_unsigned(1256,16),
    to_unsigned(1276,16),
    to_unsigned(1297,16),
    to_unsigned(1317,16),
    to_unsigned(1338,16),
    to_unsigned(1358,16),
    to_unsigned(1379,16),
    to_unsigned(1400,16),
    to_unsigned(1420,16),
    to_unsigned(1441,16),
    to_unsigned(1461,16),
    to_unsigned(1482,16),
    to_unsigned(1502,16),
    to_unsigned(1523,16),
    to_unsigned(1544,16),
    to_unsigned(1564,16),
    to_unsigned(1585,16),
    to_unsigned(1605,16),
    to_unsigned(1626,16),
    to_unsigned(1646,16),
    to_unsigned(1667,16),
    to_unsigned(1687,16),
    to_unsigned(1708,16),
    to_unsigned(1729,16),
    to_unsigned(1749,16),
    to_unsigned(1770,16),
    to_unsigned(1790,16),
    to_unsigned(1811,16),
    to_unsigned(1831,16),
    to_unsigned(1852,16),
    to_unsigned(1872,16),
    to_unsigned(1893,16),
    to_unsigned(1914,16),
    to_unsigned(1934,16),
    to_unsigned(1955,16),
    to_unsigned(1975,16),
    to_unsigned(1996,16),
    to_unsigned(2016,16),
    to_unsigned(2037,16),
    to_unsigned(2057,16),
    to_unsigned(2078,16),
    to_unsigned(2099,16),
    to_unsigned(2119,16),
    to_unsigned(2140,16),
    to_unsigned(2160,16),
    to_unsigned(2181,16),
    to_unsigned(2201,16),
    to_unsigned(2222,16),
    to_unsigned(2242,16),
    to_unsigned(2263,16),
    to_unsigned(2283,16),
    to_unsigned(2304,16),
    to_unsigned(2325,16),
    to_unsigned(2345,16),
    to_unsigned(2366,16),
    to_unsigned(2386,16),
    to_unsigned(2407,16),
    to_unsigned(2427,16),
    to_unsigned(2448,16),
    to_unsigned(2468,16),
    to_unsigned(2489,16),
    to_unsigned(2509,16),
    to_unsigned(2530,16),
    to_unsigned(2550,16),
    to_unsigned(2571,16),
    to_unsigned(2591,16),
    to_unsigned(2612,16),
    to_unsigned(2632,16),
    to_unsigned(2653,16),
    to_unsigned(2673,16),
    to_unsigned(2694,16),
    to_unsigned(2715,16),
    to_unsigned(2735,16),
    to_unsigned(2756,16),
    to_unsigned(2776,16),
    to_unsigned(2797,16),
    to_unsigned(2817,16),
    to_unsigned(2838,16),
    to_unsigned(2858,16),
    to_unsigned(2879,16),
    to_unsigned(2899,16),
    to_unsigned(2920,16),
    to_unsigned(2940,16),
    to_unsigned(2961,16),
    to_unsigned(2981,16),
    to_unsigned(3002,16),
    to_unsigned(3022,16),
    to_unsigned(3043,16),
    to_unsigned(3063,16),
    to_unsigned(3084,16),
    to_unsigned(3104,16),
    to_unsigned(3125,16),
    to_unsigned(3145,16),
    to_unsigned(3166,16),
    to_unsigned(3186,16),
    to_unsigned(3207,16),
    to_unsigned(3227,16),
    to_unsigned(3248,16),
    to_unsigned(3268,16),
    to_unsigned(3289,16),
    to_unsigned(3309,16),
    to_unsigned(3330,16),
    to_unsigned(3350,16),
    to_unsigned(3370,16),
    to_unsigned(3391,16),
    to_unsigned(3411,16),
    to_unsigned(3432,16),
    to_unsigned(3452,16),
    to_unsigned(3473,16),
    to_unsigned(3493,16),
    to_unsigned(3514,16),
    to_unsigned(3534,16),
    to_unsigned(3555,16),
    to_unsigned(3575,16),
    to_unsigned(3596,16),
    to_unsigned(3616,16),
    to_unsigned(3637,16),
    to_unsigned(3657,16),
    to_unsigned(3678,16),
    to_unsigned(3698,16),
    to_unsigned(3718,16),
    to_unsigned(3739,16),
    to_unsigned(3759,16),
    to_unsigned(3780,16),
    to_unsigned(3800,16),
    to_unsigned(3821,16),
    to_unsigned(3841,16),
    to_unsigned(3862,16),
    to_unsigned(3882,16),
    to_unsigned(3902,16),
    to_unsigned(3923,16),
    to_unsigned(3943,16),
    to_unsigned(3964,16),
    to_unsigned(3984,16),
    to_unsigned(4005,16),
    to_unsigned(4025,16),
    to_unsigned(4046,16),
    to_unsigned(4066,16),
    to_unsigned(4086,16),
    to_unsigned(4107,16),
    to_unsigned(4127,16),
    to_unsigned(4148,16),
    to_unsigned(4168,16),
    to_unsigned(4188,16),
    to_unsigned(4209,16),
    to_unsigned(4229,16),
    to_unsigned(4250,16),
    to_unsigned(4270,16),
    to_unsigned(4291,16),
    to_unsigned(4311,16),
    to_unsigned(4331,16),
    to_unsigned(4352,16),
    to_unsigned(4372,16),
    to_unsigned(4393,16),
    to_unsigned(4413,16),
    to_unsigned(4433,16),
    to_unsigned(4454,16),
    to_unsigned(4474,16),
    to_unsigned(4495,16),
    to_unsigned(4515,16),
    to_unsigned(4535,16),
    to_unsigned(4556,16),
    to_unsigned(4576,16),
    to_unsigned(4597,16),
    to_unsigned(4617,16),
    to_unsigned(4637,16),
    to_unsigned(4658,16),
    to_unsigned(4678,16),
    to_unsigned(4698,16),
    to_unsigned(4719,16),
    to_unsigned(4739,16),
    to_unsigned(4760,16),
    to_unsigned(4780,16),
    to_unsigned(4800,16),
    to_unsigned(4821,16),
    to_unsigned(4841,16),
    to_unsigned(4861,16),
    to_unsigned(4882,16),
    to_unsigned(4902,16),
    to_unsigned(4922,16),
    to_unsigned(4943,16),
    to_unsigned(4963,16),
    to_unsigned(4983,16),
    to_unsigned(5004,16),
    to_unsigned(5024,16),
    to_unsigned(5045,16),
    to_unsigned(5065,16),
    to_unsigned(5085,16),
    to_unsigned(5106,16),
    to_unsigned(5126,16),
    to_unsigned(5146,16),
    to_unsigned(5167,16),
    to_unsigned(5187,16),
    to_unsigned(5207,16),
    to_unsigned(5228,16),
    to_unsigned(5248,16),
    to_unsigned(5268,16),
    to_unsigned(5288,16),
    to_unsigned(5309,16),
    to_unsigned(5329,16),
    to_unsigned(5349,16),
    to_unsigned(5370,16),
    to_unsigned(5390,16),
    to_unsigned(5410,16),
    to_unsigned(5431,16),
    to_unsigned(5451,16),
    to_unsigned(5471,16),
    to_unsigned(5492,16),
    to_unsigned(5512,16),
    to_unsigned(5532,16),
    to_unsigned(5552,16),
    to_unsigned(5573,16),
    to_unsigned(5593,16),
    to_unsigned(5613,16),
    to_unsigned(5634,16),
    to_unsigned(5654,16),
    to_unsigned(5674,16),
    to_unsigned(5694,16),
    to_unsigned(5715,16),
    to_unsigned(5735,16),
    to_unsigned(5755,16),
    to_unsigned(5776,16),
    to_unsigned(5796,16),
    to_unsigned(5816,16),
    to_unsigned(5836,16),
    to_unsigned(5857,16),
    to_unsigned(5877,16),
    to_unsigned(5897,16),
    to_unsigned(5917,16),
    to_unsigned(5938,16),
    to_unsigned(5958,16),
    to_unsigned(5978,16),
    to_unsigned(5998,16),
    to_unsigned(6019,16),
    to_unsigned(6039,16),
    to_unsigned(6059,16),
    to_unsigned(6079,16),
    to_unsigned(6099,16),
    to_unsigned(6120,16),
    to_unsigned(6140,16),
    to_unsigned(6160,16),
    to_unsigned(6180,16),
    to_unsigned(6201,16),
    to_unsigned(6221,16),
    to_unsigned(6241,16),
    to_unsigned(6261,16),
    to_unsigned(6281,16),
    to_unsigned(6302,16),
    to_unsigned(6322,16),
    to_unsigned(6342,16),
    to_unsigned(6362,16),
    to_unsigned(6382,16),
    to_unsigned(6403,16),
    to_unsigned(6423,16),
    to_unsigned(6443,16),
    to_unsigned(6463,16),
    to_unsigned(6483,16),
    to_unsigned(6504,16),
    to_unsigned(6524,16),
    to_unsigned(6544,16),
    to_unsigned(6564,16),
    to_unsigned(6584,16),
    to_unsigned(6604,16),
    to_unsigned(6625,16),
    to_unsigned(6645,16),
    to_unsigned(6665,16),
    to_unsigned(6685,16),
    to_unsigned(6705,16),
    to_unsigned(6725,16),
    to_unsigned(6746,16),
    to_unsigned(6766,16),
    to_unsigned(6786,16),
    to_unsigned(6806,16),
    to_unsigned(6826,16),
    to_unsigned(6846,16),
    to_unsigned(6866,16),
    to_unsigned(6886,16),
    to_unsigned(6907,16),
    to_unsigned(6927,16),
    to_unsigned(6947,16),
    to_unsigned(6967,16),
    to_unsigned(6987,16),
    to_unsigned(7007,16),
    to_unsigned(7027,16),
    to_unsigned(7047,16),
    to_unsigned(7068,16),
    to_unsigned(7088,16),
    to_unsigned(7108,16),
    to_unsigned(7128,16),
    to_unsigned(7148,16),
    to_unsigned(7168,16),
    to_unsigned(7188,16),
    to_unsigned(7208,16),
    to_unsigned(7228,16),
    to_unsigned(7248,16),
    to_unsigned(7268,16),
    to_unsigned(7288,16),
    to_unsigned(7309,16),
    to_unsigned(7329,16),
    to_unsigned(7349,16),
    to_unsigned(7369,16),
    to_unsigned(7389,16),
    to_unsigned(7409,16),
    to_unsigned(7429,16),
    to_unsigned(7449,16),
    to_unsigned(7469,16),
    to_unsigned(7489,16),
    to_unsigned(7509,16),
    to_unsigned(7529,16),
    to_unsigned(7549,16),
    to_unsigned(7569,16),
    to_unsigned(7589,16),
    to_unsigned(7609,16),
    to_unsigned(7629,16),
    to_unsigned(7649,16),
    to_unsigned(7669,16),
    to_unsigned(7689,16),
    to_unsigned(7709,16),
    to_unsigned(7729,16),
    to_unsigned(7749,16),
    to_unsigned(7769,16),
    to_unsigned(7789,16),
    to_unsigned(7809,16),
    to_unsigned(7829,16),
    to_unsigned(7849,16),
    to_unsigned(7869,16),
    to_unsigned(7889,16),
    to_unsigned(7909,16),
    to_unsigned(7929,16),
    to_unsigned(7949,16),
    to_unsigned(7969,16),
    to_unsigned(7989,16),
    to_unsigned(8009,16),
    to_unsigned(8029,16),
    to_unsigned(8049,16),
    to_unsigned(8069,16),
    to_unsigned(8089,16),
    to_unsigned(8109,16),
    to_unsigned(8129,16),
    to_unsigned(8149,16),
    to_unsigned(8169,16),
    to_unsigned(8189,16),
    to_unsigned(8209,16),
    to_unsigned(8229,16),
    to_unsigned(8248,16),
    to_unsigned(8268,16),
    to_unsigned(8288,16),
    to_unsigned(8308,16),
    to_unsigned(8328,16),
    to_unsigned(8348,16),
    to_unsigned(8368,16),
    to_unsigned(8388,16),
    to_unsigned(8408,16),
    to_unsigned(8428,16),
    to_unsigned(8448,16),
    to_unsigned(8467,16),
    to_unsigned(8487,16),
    to_unsigned(8507,16),
    to_unsigned(8527,16),
    to_unsigned(8547,16),
    to_unsigned(8567,16),
    to_unsigned(8587,16),
    to_unsigned(8607,16),
    to_unsigned(8626,16),
    to_unsigned(8646,16),
    to_unsigned(8666,16),
    to_unsigned(8686,16),
    to_unsigned(8706,16),
    to_unsigned(8726,16),
    to_unsigned(8746,16),
    to_unsigned(8765,16),
    to_unsigned(8785,16),
    to_unsigned(8805,16),
    to_unsigned(8825,16),
    to_unsigned(8845,16),
    to_unsigned(8865,16),
    to_unsigned(8884,16),
    to_unsigned(8904,16),
    to_unsigned(8924,16),
    to_unsigned(8944,16),
    to_unsigned(8964,16),
    to_unsigned(8983,16),
    to_unsigned(9003,16),
    to_unsigned(9023,16),
    to_unsigned(9043,16),
    to_unsigned(9063,16),
    to_unsigned(9082,16),
    to_unsigned(9102,16),
    to_unsigned(9122,16),
    to_unsigned(9142,16),
    to_unsigned(9161,16),
    to_unsigned(9181,16),
    to_unsigned(9201,16),
    to_unsigned(9221,16),
    to_unsigned(9241,16),
    to_unsigned(9260,16),
    to_unsigned(9280,16),
    to_unsigned(9300,16),
    to_unsigned(9319,16),
    to_unsigned(9339,16),
    to_unsigned(9359,16),
    to_unsigned(9379,16),
    to_unsigned(9398,16),
    to_unsigned(9418,16),
    to_unsigned(9438,16),
    to_unsigned(9458,16),
    to_unsigned(9477,16),
    to_unsigned(9497,16),
    to_unsigned(9517,16),
    to_unsigned(9536,16),
    to_unsigned(9556,16),
    to_unsigned(9576,16),
    to_unsigned(9595,16),
    to_unsigned(9615,16),
    to_unsigned(9635,16),
    to_unsigned(9654,16),
    to_unsigned(9674,16),
    to_unsigned(9694,16),
    to_unsigned(9714,16),
    to_unsigned(9733,16),
    to_unsigned(9753,16),
    to_unsigned(9772,16),
    to_unsigned(9792,16),
    to_unsigned(9812,16),
    to_unsigned(9831,16),
    to_unsigned(9851,16),
    to_unsigned(9871,16),
    to_unsigned(9890,16),
    to_unsigned(9910,16),
    to_unsigned(9930,16),
    to_unsigned(9949,16),
    to_unsigned(9969,16),
    to_unsigned(9988,16),
    to_unsigned(10008,16),
    to_unsigned(10028,16),
    to_unsigned(10047,16),
    to_unsigned(10067,16),
    to_unsigned(10086,16),
    to_unsigned(10106,16),
    to_unsigned(10126,16),
    to_unsigned(10145,16),
    to_unsigned(10165,16),
    to_unsigned(10184,16),
    to_unsigned(10204,16),
    to_unsigned(10223,16),
    to_unsigned(10243,16),
    to_unsigned(10263,16),
    to_unsigned(10282,16),
    to_unsigned(10302,16),
    to_unsigned(10321,16),
    to_unsigned(10341,16),
    to_unsigned(10360,16),
    to_unsigned(10380,16),
    to_unsigned(10399,16),
    to_unsigned(10419,16),
    to_unsigned(10438,16),
    to_unsigned(10458,16),
    to_unsigned(10477,16),
    to_unsigned(10497,16),
    to_unsigned(10516,16),
    to_unsigned(10536,16),
    to_unsigned(10555,16),
    to_unsigned(10575,16),
    to_unsigned(10594,16),
    to_unsigned(10614,16),
    to_unsigned(10633,16),
    to_unsigned(10653,16),
    to_unsigned(10672,16),
    to_unsigned(10692,16),
    to_unsigned(10711,16),
    to_unsigned(10731,16),
    to_unsigned(10750,16),
    to_unsigned(10769,16),
    to_unsigned(10789,16),
    to_unsigned(10808,16),
    to_unsigned(10828,16),
    to_unsigned(10847,16),
    to_unsigned(10867,16),
    to_unsigned(10886,16),
    to_unsigned(10905,16),
    to_unsigned(10925,16),
    to_unsigned(10944,16),
    to_unsigned(10964,16),
    to_unsigned(10983,16),
    to_unsigned(11003,16),
    to_unsigned(11022,16),
    to_unsigned(11041,16),
    to_unsigned(11061,16),
    to_unsigned(11080,16),
    to_unsigned(11099,16),
    to_unsigned(11119,16),
    to_unsigned(11138,16),
    to_unsigned(11158,16),
    to_unsigned(11177,16),
    to_unsigned(11196,16),
    to_unsigned(11216,16),
    to_unsigned(11235,16),
    to_unsigned(11254,16),
    to_unsigned(11274,16),
    to_unsigned(11293,16),
    to_unsigned(11312,16),
    to_unsigned(11332,16),
    to_unsigned(11351,16),
    to_unsigned(11370,16),
    to_unsigned(11389,16),
    to_unsigned(11409,16),
    to_unsigned(11428,16),
    to_unsigned(11447,16),
    to_unsigned(11467,16),
    to_unsigned(11486,16),
    to_unsigned(11505,16),
    to_unsigned(11525,16),
    to_unsigned(11544,16),
    to_unsigned(11563,16),
    to_unsigned(11582,16),
    to_unsigned(11602,16),
    to_unsigned(11621,16),
    to_unsigned(11640,16),
    to_unsigned(11659,16),
    to_unsigned(11679,16),
    to_unsigned(11698,16),
    to_unsigned(11717,16),
    to_unsigned(11736,16),
    to_unsigned(11755,16),
    to_unsigned(11775,16),
    to_unsigned(11794,16),
    to_unsigned(11813,16),
    to_unsigned(11832,16),
    to_unsigned(11851,16),
    to_unsigned(11871,16),
    to_unsigned(11890,16),
    to_unsigned(11909,16),
    to_unsigned(11928,16),
    to_unsigned(11947,16),
    to_unsigned(11967,16),
    to_unsigned(11986,16),
    to_unsigned(12005,16),
    to_unsigned(12024,16),
    to_unsigned(12043,16),
    to_unsigned(12062,16),
    to_unsigned(12081,16),
    to_unsigned(12101,16),
    to_unsigned(12120,16),
    to_unsigned(12139,16),
    to_unsigned(12158,16),
    to_unsigned(12177,16),
    to_unsigned(12196,16),
    to_unsigned(12215,16),
    to_unsigned(12234,16),
    to_unsigned(12254,16),
    to_unsigned(12273,16),
    to_unsigned(12292,16),
    to_unsigned(12311,16),
    to_unsigned(12330,16),
    to_unsigned(12349,16),
    to_unsigned(12368,16),
    to_unsigned(12387,16),
    to_unsigned(12406,16),
    to_unsigned(12425,16),
    to_unsigned(12444,16),
    to_unsigned(12463,16),
    to_unsigned(12482,16),
    to_unsigned(12501,16),
    to_unsigned(12520,16),
    to_unsigned(12539,16),
    to_unsigned(12558,16),
    to_unsigned(12577,16),
    to_unsigned(12596,16),
    to_unsigned(12615,16),
    to_unsigned(12634,16),
    to_unsigned(12653,16),
    to_unsigned(12672,16),
    to_unsigned(12691,16),
    to_unsigned(12710,16),
    to_unsigned(12729,16),
    to_unsigned(12748,16),
    to_unsigned(12767,16),
    to_unsigned(12786,16),
    to_unsigned(12805,16),
    to_unsigned(12824,16),
    to_unsigned(12843,16),
    to_unsigned(12862,16),
    to_unsigned(12881,16),
    to_unsigned(12900,16),
    to_unsigned(12919,16),
    to_unsigned(12938,16),
    to_unsigned(12957,16),
    to_unsigned(12976,16),
    to_unsigned(12994,16),
    to_unsigned(13013,16),
    to_unsigned(13032,16),
    to_unsigned(13051,16),
    to_unsigned(13070,16),
    to_unsigned(13089,16),
    to_unsigned(13108,16),
    to_unsigned(13127,16),
    to_unsigned(13145,16),
    to_unsigned(13164,16),
    to_unsigned(13183,16),
    to_unsigned(13202,16),
    to_unsigned(13221,16),
    to_unsigned(13240,16),
    to_unsigned(13259,16),
    to_unsigned(13277,16),
    to_unsigned(13296,16),
    to_unsigned(13315,16),
    to_unsigned(13334,16),
    to_unsigned(13353,16),
    to_unsigned(13371,16),
    to_unsigned(13390,16),
    to_unsigned(13409,16),
    to_unsigned(13428,16),
    to_unsigned(13447,16),
    to_unsigned(13465,16),
    to_unsigned(13484,16),
    to_unsigned(13503,16),
    to_unsigned(13522,16),
    to_unsigned(13540,16),
    to_unsigned(13559,16),
    to_unsigned(13578,16),
    to_unsigned(13597,16),
    to_unsigned(13615,16),
    to_unsigned(13634,16),
    to_unsigned(13653,16),
    to_unsigned(13671,16),
    to_unsigned(13690,16),
    to_unsigned(13709,16),
    to_unsigned(13728,16),
    to_unsigned(13746,16),
    to_unsigned(13765,16),
    to_unsigned(13784,16),
    to_unsigned(13802,16),
    to_unsigned(13821,16),
    to_unsigned(13840,16),
    to_unsigned(13858,16),
    to_unsigned(13877,16),
    to_unsigned(13896,16),
    to_unsigned(13914,16),
    to_unsigned(13933,16),
    to_unsigned(13952,16),
    to_unsigned(13970,16),
    to_unsigned(13989,16),
    to_unsigned(14007,16),
    to_unsigned(14026,16),
    to_unsigned(14045,16),
    to_unsigned(14063,16),
    to_unsigned(14082,16),
    to_unsigned(14100,16),
    to_unsigned(14119,16),
    to_unsigned(14138,16),
    to_unsigned(14156,16),
    to_unsigned(14175,16),
    to_unsigned(14193,16),
    to_unsigned(14212,16),
    to_unsigned(14230,16),
    to_unsigned(14249,16),
    to_unsigned(14267,16),
    to_unsigned(14286,16),
    to_unsigned(14304,16),
    to_unsigned(14323,16),
    to_unsigned(14341,16),
    to_unsigned(14360,16),
    to_unsigned(14378,16),
    to_unsigned(14397,16),
    to_unsigned(14415,16),
    to_unsigned(14434,16),
    to_unsigned(14452,16),
    to_unsigned(14471,16),
    to_unsigned(14489,16),
    to_unsigned(14508,16),
    to_unsigned(14526,16),
    to_unsigned(14545,16),
    to_unsigned(14563,16),
    to_unsigned(14582,16),
    to_unsigned(14600,16),
    to_unsigned(14619,16),
    to_unsigned(14637,16),
    to_unsigned(14655,16),
    to_unsigned(14674,16),
    to_unsigned(14692,16),
    to_unsigned(14711,16),
    to_unsigned(14729,16),
    to_unsigned(14747,16),
    to_unsigned(14766,16),
    to_unsigned(14784,16),
    to_unsigned(14802,16),
    to_unsigned(14821,16),
    to_unsigned(14839,16),
    to_unsigned(14858,16),
    to_unsigned(14876,16),
    to_unsigned(14894,16),
    to_unsigned(14913,16),
    to_unsigned(14931,16),
    to_unsigned(14949,16),
    to_unsigned(14968,16),
    to_unsigned(14986,16),
    to_unsigned(15004,16),
    to_unsigned(15022,16),
    to_unsigned(15041,16),
    to_unsigned(15059,16),
    to_unsigned(15077,16),
    to_unsigned(15096,16),
    to_unsigned(15114,16),
    to_unsigned(15132,16),
    to_unsigned(15150,16),
    to_unsigned(15169,16),
    to_unsigned(15187,16),
    to_unsigned(15205,16),
    to_unsigned(15223,16),
    to_unsigned(15242,16),
    to_unsigned(15260,16),
    to_unsigned(15278,16),
    to_unsigned(15296,16),
    to_unsigned(15314,16),
    to_unsigned(15333,16),
    to_unsigned(15351,16),
    to_unsigned(15369,16),
    to_unsigned(15387,16),
    to_unsigned(15405,16),
    to_unsigned(15424,16),
    to_unsigned(15442,16),
    to_unsigned(15460,16),
    to_unsigned(15478,16),
    to_unsigned(15496,16),
    to_unsigned(15514,16),
    to_unsigned(15532,16),
    to_unsigned(15551,16),
    to_unsigned(15569,16),
    to_unsigned(15587,16),
    to_unsigned(15605,16),
    to_unsigned(15623,16),
    to_unsigned(15641,16),
    to_unsigned(15659,16),
    to_unsigned(15677,16),
    to_unsigned(15695,16),
    to_unsigned(15713,16),
    to_unsigned(15731,16),
    to_unsigned(15750,16),
    to_unsigned(15768,16),
    to_unsigned(15786,16),
    to_unsigned(15804,16),
    to_unsigned(15822,16),
    to_unsigned(15840,16),
    to_unsigned(15858,16),
    to_unsigned(15876,16),
    to_unsigned(15894,16),
    to_unsigned(15912,16),
    to_unsigned(15930,16),
    to_unsigned(15948,16),
    to_unsigned(15966,16),
    to_unsigned(15984,16),
    to_unsigned(16002,16),
    to_unsigned(16020,16),
    to_unsigned(16038,16),
    to_unsigned(16056,16),
    to_unsigned(16073,16),
    to_unsigned(16091,16),
    to_unsigned(16109,16),
    to_unsigned(16127,16),
    to_unsigned(16145,16),
    to_unsigned(16163,16),
    to_unsigned(16181,16),
    to_unsigned(16199,16),
    to_unsigned(16217,16),
    to_unsigned(16235,16),
    to_unsigned(16253,16),
    to_unsigned(16270,16),
    to_unsigned(16288,16),
    to_unsigned(16306,16),
    to_unsigned(16324,16),
    to_unsigned(16342,16),
    to_unsigned(16360,16),
    to_unsigned(16378,16),
    to_unsigned(16395,16),
    to_unsigned(16413,16),
    to_unsigned(16431,16),
    to_unsigned(16449,16),
    to_unsigned(16467,16),
    to_unsigned(16484,16),
    to_unsigned(16502,16),
    to_unsigned(16520,16),
    to_unsigned(16538,16),
    to_unsigned(16556,16),
    to_unsigned(16573,16),
    to_unsigned(16591,16),
    to_unsigned(16609,16),
    to_unsigned(16627,16),
    to_unsigned(16644,16),
    to_unsigned(16662,16),
    to_unsigned(16680,16),
    to_unsigned(16697,16),
    to_unsigned(16715,16),
    to_unsigned(16733,16),
    to_unsigned(16751,16),
    to_unsigned(16768,16),
    to_unsigned(16786,16),
    to_unsigned(16804,16),
    to_unsigned(16821,16),
    to_unsigned(16839,16),
    to_unsigned(16857,16),
    to_unsigned(16874,16),
    to_unsigned(16892,16),
    to_unsigned(16910,16),
    to_unsigned(16927,16),
    to_unsigned(16945,16),
    to_unsigned(16962,16),
    to_unsigned(16980,16),
    to_unsigned(16998,16),
    to_unsigned(17015,16),
    to_unsigned(17033,16),
    to_unsigned(17050,16),
    to_unsigned(17068,16),
    to_unsigned(17086,16),
    to_unsigned(17103,16),
    to_unsigned(17121,16),
    to_unsigned(17138,16),
    to_unsigned(17156,16),
    to_unsigned(17173,16),
    to_unsigned(17191,16),
    to_unsigned(17208,16),
    to_unsigned(17226,16),
    to_unsigned(17243,16),
    to_unsigned(17261,16),
    to_unsigned(17278,16),
    to_unsigned(17296,16),
    to_unsigned(17313,16),
    to_unsigned(17331,16),
    to_unsigned(17348,16),
    to_unsigned(17366,16),
    to_unsigned(17383,16),
    to_unsigned(17401,16),
    to_unsigned(17418,16),
    to_unsigned(17436,16),
    to_unsigned(17453,16),
    to_unsigned(17470,16),
    to_unsigned(17488,16),
    to_unsigned(17505,16),
    to_unsigned(17523,16),
    to_unsigned(17540,16),
    to_unsigned(17557,16),
    to_unsigned(17575,16),
    to_unsigned(17592,16),
    to_unsigned(17610,16),
    to_unsigned(17627,16),
    to_unsigned(17644,16),
    to_unsigned(17662,16),
    to_unsigned(17679,16),
    to_unsigned(17696,16),
    to_unsigned(17714,16),
    to_unsigned(17731,16),
    to_unsigned(17748,16),
    to_unsigned(17766,16),
    to_unsigned(17783,16),
    to_unsigned(17800,16),
    to_unsigned(17817,16),
    to_unsigned(17835,16),
    to_unsigned(17852,16),
    to_unsigned(17869,16),
    to_unsigned(17886,16),
    to_unsigned(17904,16),
    to_unsigned(17921,16),
    to_unsigned(17938,16),
    to_unsigned(17955,16),
    to_unsigned(17973,16),
    to_unsigned(17990,16),
    to_unsigned(18007,16),
    to_unsigned(18024,16),
    to_unsigned(18041,16),
    to_unsigned(18059,16),
    to_unsigned(18076,16),
    to_unsigned(18093,16),
    to_unsigned(18110,16),
    to_unsigned(18127,16),
    to_unsigned(18144,16),
    to_unsigned(18162,16),
    to_unsigned(18179,16),
    to_unsigned(18196,16),
    to_unsigned(18213,16),
    to_unsigned(18230,16),
    to_unsigned(18247,16),
    to_unsigned(18264,16),
    to_unsigned(18281,16),
    to_unsigned(18298,16),
    to_unsigned(18315,16),
    to_unsigned(18333,16),
    to_unsigned(18350,16),
    to_unsigned(18367,16),
    to_unsigned(18384,16),
    to_unsigned(18401,16),
    to_unsigned(18418,16),
    to_unsigned(18435,16),
    to_unsigned(18452,16),
    to_unsigned(18469,16),
    to_unsigned(18486,16),
    to_unsigned(18503,16),
    to_unsigned(18520,16),
    to_unsigned(18537,16),
    to_unsigned(18554,16),
    to_unsigned(18571,16),
    to_unsigned(18588,16),
    to_unsigned(18605,16),
    to_unsigned(18622,16),
    to_unsigned(18639,16),
    to_unsigned(18655,16),
    to_unsigned(18672,16),
    to_unsigned(18689,16),
    to_unsigned(18706,16),
    to_unsigned(18723,16),
    to_unsigned(18740,16),
    to_unsigned(18757,16),
    to_unsigned(18774,16),
    to_unsigned(18791,16),
    to_unsigned(18807,16),
    to_unsigned(18824,16),
    to_unsigned(18841,16),
    to_unsigned(18858,16),
    to_unsigned(18875,16),
    to_unsigned(18892,16),
    to_unsigned(18909,16),
    to_unsigned(18925,16),
    to_unsigned(18942,16),
    to_unsigned(18959,16),
    to_unsigned(18976,16),
    to_unsigned(18992,16),
    to_unsigned(19009,16),
    to_unsigned(19026,16),
    to_unsigned(19043,16),
    to_unsigned(19060,16),
    to_unsigned(19076,16),
    to_unsigned(19093,16),
    to_unsigned(19110,16),
    to_unsigned(19126,16),
    to_unsigned(19143,16),
    to_unsigned(19160,16),
    to_unsigned(19177,16),
    to_unsigned(19193,16),
    to_unsigned(19210,16),
    to_unsigned(19227,16),
    to_unsigned(19243,16),
    to_unsigned(19260,16),
    to_unsigned(19277,16),
    to_unsigned(19293,16),
    to_unsigned(19310,16),
    to_unsigned(19327,16),
    to_unsigned(19343,16),
    to_unsigned(19360,16),
    to_unsigned(19376,16),
    to_unsigned(19393,16),
    to_unsigned(19410,16),
    to_unsigned(19426,16),
    to_unsigned(19443,16),
    to_unsigned(19459,16),
    to_unsigned(19476,16),
    to_unsigned(19492,16),
    to_unsigned(19509,16),
    to_unsigned(19525,16),
    to_unsigned(19542,16),
    to_unsigned(19559,16),
    to_unsigned(19575,16),
    to_unsigned(19592,16),
    to_unsigned(19608,16),
    to_unsigned(19625,16),
    to_unsigned(19641,16),
    to_unsigned(19658,16),
    to_unsigned(19674,16),
    to_unsigned(19690,16),
    to_unsigned(19707,16),
    to_unsigned(19723,16),
    to_unsigned(19740,16),
    to_unsigned(19756,16),
    to_unsigned(19773,16),
    to_unsigned(19789,16),
    to_unsigned(19805,16),
    to_unsigned(19822,16),
    to_unsigned(19838,16),
    to_unsigned(19855,16),
    to_unsigned(19871,16),
    to_unsigned(19887,16),
    to_unsigned(19904,16),
    to_unsigned(19920,16),
    to_unsigned(19936,16),
    to_unsigned(19953,16),
    to_unsigned(19969,16),
    to_unsigned(19985,16),
    to_unsigned(20002,16),
    to_unsigned(20018,16),
    to_unsigned(20034,16),
    to_unsigned(20051,16),
    to_unsigned(20067,16),
    to_unsigned(20083,16),
    to_unsigned(20099,16),
    to_unsigned(20116,16),
    to_unsigned(20132,16),
    to_unsigned(20148,16),
    to_unsigned(20164,16),
    to_unsigned(20181,16),
    to_unsigned(20197,16),
    to_unsigned(20213,16),
    to_unsigned(20229,16),
    to_unsigned(20245,16),
    to_unsigned(20262,16),
    to_unsigned(20278,16),
    to_unsigned(20294,16),
    to_unsigned(20310,16),
    to_unsigned(20326,16),
    to_unsigned(20342,16),
    to_unsigned(20359,16),
    to_unsigned(20375,16),
    to_unsigned(20391,16),
    to_unsigned(20407,16),
    to_unsigned(20423,16),
    to_unsigned(20439,16),
    to_unsigned(20455,16),
    to_unsigned(20471,16),
    to_unsigned(20487,16),
    to_unsigned(20503,16),
    to_unsigned(20519,16),
    to_unsigned(20535,16),
    to_unsigned(20552,16),
    to_unsigned(20568,16),
    to_unsigned(20584,16),
    to_unsigned(20600,16),
    to_unsigned(20616,16),
    to_unsigned(20632,16),
    to_unsigned(20648,16),
    to_unsigned(20664,16),
    to_unsigned(20680,16),
    to_unsigned(20696,16),
    to_unsigned(20711,16),
    to_unsigned(20727,16),
    to_unsigned(20743,16),
    to_unsigned(20759,16),
    to_unsigned(20775,16),
    to_unsigned(20791,16),
    to_unsigned(20807,16),
    to_unsigned(20823,16),
    to_unsigned(20839,16),
    to_unsigned(20855,16),
    to_unsigned(20871,16),
    to_unsigned(20886,16),
    to_unsigned(20902,16),
    to_unsigned(20918,16),
    to_unsigned(20934,16),
    to_unsigned(20950,16),
    to_unsigned(20966,16),
    to_unsigned(20982,16),
    to_unsigned(20997,16),
    to_unsigned(21013,16),
    to_unsigned(21029,16),
    to_unsigned(21045,16),
    to_unsigned(21060,16),
    to_unsigned(21076,16),
    to_unsigned(21092,16),
    to_unsigned(21108,16),
    to_unsigned(21123,16),
    to_unsigned(21139,16),
    to_unsigned(21155,16),
    to_unsigned(21171,16),
    to_unsigned(21186,16),
    to_unsigned(21202,16),
    to_unsigned(21218,16),
    to_unsigned(21233,16),
    to_unsigned(21249,16),
    to_unsigned(21265,16),
    to_unsigned(21280,16),
    to_unsigned(21296,16),
    to_unsigned(21312,16),
    to_unsigned(21327,16),
    to_unsigned(21343,16),
    to_unsigned(21359,16),
    to_unsigned(21374,16),
    to_unsigned(21390,16),
    to_unsigned(21405,16),
    to_unsigned(21421,16),
    to_unsigned(21437,16),
    to_unsigned(21452,16),
    to_unsigned(21468,16),
    to_unsigned(21483,16),
    to_unsigned(21499,16),
    to_unsigned(21514,16),
    to_unsigned(21530,16),
    to_unsigned(21545,16),
    to_unsigned(21561,16),
    to_unsigned(21576,16),
    to_unsigned(21592,16),
    to_unsigned(21607,16),
    to_unsigned(21623,16),
    to_unsigned(21638,16),
    to_unsigned(21654,16),
    to_unsigned(21669,16),
    to_unsigned(21685,16),
    to_unsigned(21700,16),
    to_unsigned(21715,16),
    to_unsigned(21731,16),
    to_unsigned(21746,16),
    to_unsigned(21762,16),
    to_unsigned(21777,16),
    to_unsigned(21792,16),
    to_unsigned(21808,16),
    to_unsigned(21823,16),
    to_unsigned(21839,16),
    to_unsigned(21854,16),
    to_unsigned(21869,16),
    to_unsigned(21885,16),
    to_unsigned(21900,16),
    to_unsigned(21915,16),
    to_unsigned(21931,16),
    to_unsigned(21946,16),
    to_unsigned(21961,16),
    to_unsigned(21976,16),
    to_unsigned(21992,16),
    to_unsigned(22007,16),
    to_unsigned(22022,16),
    to_unsigned(22037,16),
    to_unsigned(22053,16),
    to_unsigned(22068,16),
    to_unsigned(22083,16),
    to_unsigned(22098,16),
    to_unsigned(22113,16),
    to_unsigned(22129,16),
    to_unsigned(22144,16),
    to_unsigned(22159,16),
    to_unsigned(22174,16),
    to_unsigned(22189,16),
    to_unsigned(22204,16),
    to_unsigned(22220,16),
    to_unsigned(22235,16),
    to_unsigned(22250,16),
    to_unsigned(22265,16),
    to_unsigned(22280,16),
    to_unsigned(22295,16),
    to_unsigned(22310,16),
    to_unsigned(22325,16),
    to_unsigned(22340,16),
    to_unsigned(22355,16),
    to_unsigned(22370,16),
    to_unsigned(22385,16),
    to_unsigned(22401,16),
    to_unsigned(22416,16),
    to_unsigned(22431,16),
    to_unsigned(22446,16),
    to_unsigned(22461,16),
    to_unsigned(22476,16),
    to_unsigned(22491,16),
    to_unsigned(22505,16),
    to_unsigned(22520,16),
    to_unsigned(22535,16),
    to_unsigned(22550,16),
    to_unsigned(22565,16),
    to_unsigned(22580,16),
    to_unsigned(22595,16),
    to_unsigned(22610,16),
    to_unsigned(22625,16),
    to_unsigned(22640,16),
    to_unsigned(22655,16),
    to_unsigned(22670,16),
    to_unsigned(22684,16),
    to_unsigned(22699,16),
    to_unsigned(22714,16),
    to_unsigned(22729,16),
    to_unsigned(22744,16),
    to_unsigned(22759,16),
    to_unsigned(22773,16),
    to_unsigned(22788,16),
    to_unsigned(22803,16),
    to_unsigned(22818,16),
    to_unsigned(22833,16),
    to_unsigned(22847,16),
    to_unsigned(22862,16),
    to_unsigned(22877,16),
    to_unsigned(22892,16),
    to_unsigned(22906,16),
    to_unsigned(22921,16),
    to_unsigned(22936,16),
    to_unsigned(22950,16),
    to_unsigned(22965,16),
    to_unsigned(22980,16),
    to_unsigned(22994,16),
    to_unsigned(23009,16),
    to_unsigned(23024,16),
    to_unsigned(23038,16),
    to_unsigned(23053,16),
    to_unsigned(23068,16),
    to_unsigned(23082,16),
    to_unsigned(23097,16),
    to_unsigned(23111,16),
    to_unsigned(23126,16),
    to_unsigned(23141,16),
    to_unsigned(23155,16),
    to_unsigned(23170,16),
    to_unsigned(23184,16),
    to_unsigned(23199,16),
    to_unsigned(23213,16),
    to_unsigned(23228,16),
    to_unsigned(23242,16),
    to_unsigned(23257,16),
    to_unsigned(23271,16),
    to_unsigned(23286,16),
    to_unsigned(23300,16),
    to_unsigned(23315,16),
    to_unsigned(23329,16),
    to_unsigned(23344,16),
    to_unsigned(23358,16),
    to_unsigned(23373,16),
    to_unsigned(23387,16),
    to_unsigned(23402,16),
    to_unsigned(23416,16),
    to_unsigned(23430,16),
    to_unsigned(23445,16),
    to_unsigned(23459,16),
    to_unsigned(23473,16),
    to_unsigned(23488,16),
    to_unsigned(23502,16),
    to_unsigned(23517,16),
    to_unsigned(23531,16),
    to_unsigned(23545,16),
    to_unsigned(23559,16),
    to_unsigned(23574,16),
    to_unsigned(23588,16),
    to_unsigned(23602,16),
    to_unsigned(23617,16),
    to_unsigned(23631,16),
    to_unsigned(23645,16),
    to_unsigned(23659,16),
    to_unsigned(23674,16),
    to_unsigned(23688,16),
    to_unsigned(23702,16),
    to_unsigned(23716,16),
    to_unsigned(23731,16),
    to_unsigned(23745,16),
    to_unsigned(23759,16),
    to_unsigned(23773,16),
    to_unsigned(23787,16),
    to_unsigned(23801,16),
    to_unsigned(23816,16),
    to_unsigned(23830,16),
    to_unsigned(23844,16),
    to_unsigned(23858,16),
    to_unsigned(23872,16),
    to_unsigned(23886,16),
    to_unsigned(23900,16),
    to_unsigned(23914,16),
    to_unsigned(23928,16),
    to_unsigned(23942,16),
    to_unsigned(23956,16),
    to_unsigned(23971,16),
    to_unsigned(23985,16),
    to_unsigned(23999,16),
    to_unsigned(24013,16),
    to_unsigned(24027,16),
    to_unsigned(24041,16),
    to_unsigned(24055,16),
    to_unsigned(24069,16),
    to_unsigned(24082,16),
    to_unsigned(24096,16),
    to_unsigned(24110,16),
    to_unsigned(24124,16),
    to_unsigned(24138,16),
    to_unsigned(24152,16),
    to_unsigned(24166,16),
    to_unsigned(24180,16),
    to_unsigned(24194,16),
    to_unsigned(24208,16),
    to_unsigned(24222,16),
    to_unsigned(24235,16),
    to_unsigned(24249,16),
    to_unsigned(24263,16),
    to_unsigned(24277,16),
    to_unsigned(24291,16),
    to_unsigned(24305,16),
    to_unsigned(24318,16),
    to_unsigned(24332,16),
    to_unsigned(24346,16),
    to_unsigned(24360,16),
    to_unsigned(24374,16),
    to_unsigned(24387,16),
    to_unsigned(24401,16),
    to_unsigned(24415,16),
    to_unsigned(24429,16),
    to_unsigned(24442,16),
    to_unsigned(24456,16),
    to_unsigned(24470,16),
    to_unsigned(24483,16),
    to_unsigned(24497,16),
    to_unsigned(24511,16),
    to_unsigned(24524,16),
    to_unsigned(24538,16),
    to_unsigned(24552,16),
    to_unsigned(24565,16),
    to_unsigned(24579,16),
    to_unsigned(24592,16),
    to_unsigned(24606,16),
    to_unsigned(24620,16),
    to_unsigned(24633,16),
    to_unsigned(24647,16),
    to_unsigned(24660,16),
    to_unsigned(24674,16),
    to_unsigned(24687,16),
    to_unsigned(24701,16),
    to_unsigned(24715,16),
    to_unsigned(24728,16),
    to_unsigned(24742,16),
    to_unsigned(24755,16),
    to_unsigned(24769,16),
    to_unsigned(24782,16),
    to_unsigned(24795,16),
    to_unsigned(24809,16),
    to_unsigned(24822,16),
    to_unsigned(24836,16),
    to_unsigned(24849,16),
    to_unsigned(24863,16),
    to_unsigned(24876,16),
    to_unsigned(24889,16),
    to_unsigned(24903,16),
    to_unsigned(24916,16),
    to_unsigned(24930,16),
    to_unsigned(24943,16),
    to_unsigned(24956,16),
    to_unsigned(24970,16),
    to_unsigned(24983,16),
    to_unsigned(24996,16),
    to_unsigned(25010,16),
    to_unsigned(25023,16),
    to_unsigned(25036,16),
    to_unsigned(25049,16),
    to_unsigned(25063,16),
    to_unsigned(25076,16),
    to_unsigned(25089,16),
    to_unsigned(25102,16),
    to_unsigned(25116,16),
    to_unsigned(25129,16),
    to_unsigned(25142,16),
    to_unsigned(25155,16),
    to_unsigned(25168,16),
    to_unsigned(25182,16),
    to_unsigned(25195,16),
    to_unsigned(25208,16),
    to_unsigned(25221,16),
    to_unsigned(25234,16),
    to_unsigned(25247,16),
    to_unsigned(25261,16),
    to_unsigned(25274,16),
    to_unsigned(25287,16),
    to_unsigned(25300,16),
    to_unsigned(25313,16),
    to_unsigned(25326,16),
    to_unsigned(25339,16),
    to_unsigned(25352,16),
    to_unsigned(25365,16),
    to_unsigned(25378,16),
    to_unsigned(25391,16),
    to_unsigned(25404,16),
    to_unsigned(25417,16),
    to_unsigned(25430,16),
    to_unsigned(25443,16),
    to_unsigned(25456,16),
    to_unsigned(25469,16),
    to_unsigned(25482,16),
    to_unsigned(25495,16),
    to_unsigned(25508,16),
    to_unsigned(25521,16),
    to_unsigned(25534,16),
    to_unsigned(25547,16),
    to_unsigned(25559,16),
    to_unsigned(25572,16),
    to_unsigned(25585,16),
    to_unsigned(25598,16),
    to_unsigned(25611,16),
    to_unsigned(25624,16),
    to_unsigned(25637,16),
    to_unsigned(25649,16),
    to_unsigned(25662,16),
    to_unsigned(25675,16),
    to_unsigned(25688,16),
    to_unsigned(25701,16),
    to_unsigned(25713,16),
    to_unsigned(25726,16),
    to_unsigned(25739,16),
    to_unsigned(25752,16),
    to_unsigned(25764,16),
    to_unsigned(25777,16),
    to_unsigned(25790,16),
    to_unsigned(25802,16),
    to_unsigned(25815,16),
    to_unsigned(25828,16),
    to_unsigned(25840,16),
    to_unsigned(25853,16),
    to_unsigned(25866,16),
    to_unsigned(25878,16),
    to_unsigned(25891,16),
    to_unsigned(25904,16),
    to_unsigned(25916,16),
    to_unsigned(25929,16),
    to_unsigned(25941,16),
    to_unsigned(25954,16),
    to_unsigned(25967,16),
    to_unsigned(25979,16),
    to_unsigned(25992,16),
    to_unsigned(26004,16),
    to_unsigned(26017,16),
    to_unsigned(26029,16),
    to_unsigned(26042,16),
    to_unsigned(26054,16),
    to_unsigned(26067,16),
    to_unsigned(26079,16),
    to_unsigned(26092,16),
    to_unsigned(26104,16),
    to_unsigned(26116,16),
    to_unsigned(26129,16),
    to_unsigned(26141,16),
    to_unsigned(26154,16),
    to_unsigned(26166,16),
    to_unsigned(26179,16),
    to_unsigned(26191,16),
    to_unsigned(26203,16),
    to_unsigned(26216,16),
    to_unsigned(26228,16),
    to_unsigned(26240,16),
    to_unsigned(26253,16),
    to_unsigned(26265,16),
    to_unsigned(26277,16),
    to_unsigned(26290,16),
    to_unsigned(26302,16),
    to_unsigned(26314,16),
    to_unsigned(26326,16),
    to_unsigned(26339,16),
    to_unsigned(26351,16),
    to_unsigned(26363,16),
    to_unsigned(26375,16),
    to_unsigned(26388,16),
    to_unsigned(26400,16),
    to_unsigned(26412,16),
    to_unsigned(26424,16),
    to_unsigned(26436,16),
    to_unsigned(26448,16),
    to_unsigned(26461,16),
    to_unsigned(26473,16),
    to_unsigned(26485,16),
    to_unsigned(26497,16),
    to_unsigned(26509,16),
    to_unsigned(26521,16),
    to_unsigned(26533,16),
    to_unsigned(26545,16),
    to_unsigned(26557,16),
    to_unsigned(26569,16),
    to_unsigned(26581,16),
    to_unsigned(26594,16),
    to_unsigned(26606,16),
    to_unsigned(26618,16),
    to_unsigned(26630,16),
    to_unsigned(26642,16),
    to_unsigned(26654,16),
    to_unsigned(26665,16),
    to_unsigned(26677,16),
    to_unsigned(26689,16),
    to_unsigned(26701,16),
    to_unsigned(26713,16),
    to_unsigned(26725,16),
    to_unsigned(26737,16),
    to_unsigned(26749,16),
    to_unsigned(26761,16),
    to_unsigned(26773,16),
    to_unsigned(26785,16),
    to_unsigned(26796,16),
    to_unsigned(26808,16),
    to_unsigned(26820,16),
    to_unsigned(26832,16),
    to_unsigned(26844,16),
    to_unsigned(26856,16),
    to_unsigned(26867,16),
    to_unsigned(26879,16),
    to_unsigned(26891,16),
    to_unsigned(26903,16),
    to_unsigned(26914,16),
    to_unsigned(26926,16),
    to_unsigned(26938,16),
    to_unsigned(26950,16),
    to_unsigned(26961,16),
    to_unsigned(26973,16),
    to_unsigned(26985,16),
    to_unsigned(26996,16),
    to_unsigned(27008,16),
    to_unsigned(27020,16),
    to_unsigned(27031,16),
    to_unsigned(27043,16),
    to_unsigned(27055,16),
    to_unsigned(27066,16),
    to_unsigned(27078,16),
    to_unsigned(27089,16),
    to_unsigned(27101,16),
    to_unsigned(27113,16),
    to_unsigned(27124,16),
    to_unsigned(27136,16),
    to_unsigned(27147,16),
    to_unsigned(27159,16),
    to_unsigned(27170,16),
    to_unsigned(27182,16),
    to_unsigned(27193,16),
    to_unsigned(27205,16),
    to_unsigned(27216,16),
    to_unsigned(27228,16),
    to_unsigned(27239,16),
    to_unsigned(27250,16),
    to_unsigned(27262,16),
    to_unsigned(27273,16),
    to_unsigned(27285,16),
    to_unsigned(27296,16),
    to_unsigned(27308,16),
    to_unsigned(27319,16),
    to_unsigned(27330,16),
    to_unsigned(27342,16),
    to_unsigned(27353,16),
    to_unsigned(27364,16),
    to_unsigned(27376,16),
    to_unsigned(27387,16),
    to_unsigned(27398,16),
    to_unsigned(27409,16),
    to_unsigned(27421,16),
    to_unsigned(27432,16),
    to_unsigned(27443,16),
    to_unsigned(27455,16),
    to_unsigned(27466,16),
    to_unsigned(27477,16),
    to_unsigned(27488,16),
    to_unsigned(27499,16),
    to_unsigned(27511,16),
    to_unsigned(27522,16),
    to_unsigned(27533,16),
    to_unsigned(27544,16),
    to_unsigned(27555,16),
    to_unsigned(27566,16),
    to_unsigned(27577,16),
    to_unsigned(27589,16),
    to_unsigned(27600,16),
    to_unsigned(27611,16),
    to_unsigned(27622,16),
    to_unsigned(27633,16),
    to_unsigned(27644,16),
    to_unsigned(27655,16),
    to_unsigned(27666,16),
    to_unsigned(27677,16),
    to_unsigned(27688,16),
    to_unsigned(27699,16),
    to_unsigned(27710,16),
    to_unsigned(27721,16),
    to_unsigned(27732,16),
    to_unsigned(27743,16),
    to_unsigned(27754,16),
    to_unsigned(27765,16),
    to_unsigned(27776,16),
    to_unsigned(27787,16),
    to_unsigned(27798,16),
    to_unsigned(27809,16),
    to_unsigned(27819,16),
    to_unsigned(27830,16),
    to_unsigned(27841,16),
    to_unsigned(27852,16),
    to_unsigned(27863,16),
    to_unsigned(27874,16),
    to_unsigned(27885,16),
    to_unsigned(27895,16),
    to_unsigned(27906,16),
    to_unsigned(27917,16),
    to_unsigned(27928,16),
    to_unsigned(27938,16),
    to_unsigned(27949,16),
    to_unsigned(27960,16),
    to_unsigned(27971,16),
    to_unsigned(27981,16),
    to_unsigned(27992,16),
    to_unsigned(28003,16),
    to_unsigned(28013,16),
    to_unsigned(28024,16),
    to_unsigned(28035,16),
    to_unsigned(28045,16),
    to_unsigned(28056,16),
    to_unsigned(28067,16),
    to_unsigned(28077,16),
    to_unsigned(28088,16),
    to_unsigned(28099,16),
    to_unsigned(28109,16),
    to_unsigned(28120,16),
    to_unsigned(28130,16),
    to_unsigned(28141,16),
    to_unsigned(28151,16),
    to_unsigned(28162,16),
    to_unsigned(28172,16),
    to_unsigned(28183,16),
    to_unsigned(28193,16),
    to_unsigned(28204,16),
    to_unsigned(28214,16),
    to_unsigned(28225,16),
    to_unsigned(28235,16),
    to_unsigned(28246,16),
    to_unsigned(28256,16),
    to_unsigned(28267,16),
    to_unsigned(28277,16),
    to_unsigned(28287,16),
    to_unsigned(28298,16),
    to_unsigned(28308,16),
    to_unsigned(28319,16),
    to_unsigned(28329,16),
    to_unsigned(28339,16),
    to_unsigned(28350,16),
    to_unsigned(28360,16),
    to_unsigned(28370,16),
    to_unsigned(28380,16),
    to_unsigned(28391,16),
    to_unsigned(28401,16),
    to_unsigned(28411,16),
    to_unsigned(28422,16),
    to_unsigned(28432,16),
    to_unsigned(28442,16),
    to_unsigned(28452,16),
    to_unsigned(28462,16),
    to_unsigned(28473,16),
    to_unsigned(28483,16),
    to_unsigned(28493,16),
    to_unsigned(28503,16),
    to_unsigned(28513,16),
    to_unsigned(28523,16),
    to_unsigned(28534,16),
    to_unsigned(28544,16),
    to_unsigned(28554,16),
    to_unsigned(28564,16),
    to_unsigned(28574,16),
    to_unsigned(28584,16),
    to_unsigned(28594,16),
    to_unsigned(28604,16),
    to_unsigned(28614,16),
    to_unsigned(28624,16),
    to_unsigned(28634,16),
    to_unsigned(28644,16),
    to_unsigned(28654,16),
    to_unsigned(28664,16),
    to_unsigned(28674,16),
    to_unsigned(28684,16),
    to_unsigned(28694,16),
    to_unsigned(28704,16),
    to_unsigned(28714,16),
    to_unsigned(28724,16),
    to_unsigned(28734,16),
    to_unsigned(28744,16),
    to_unsigned(28754,16),
    to_unsigned(28763,16),
    to_unsigned(28773,16),
    to_unsigned(28783,16),
    to_unsigned(28793,16),
    to_unsigned(28803,16),
    to_unsigned(28813,16),
    to_unsigned(28822,16),
    to_unsigned(28832,16),
    to_unsigned(28842,16),
    to_unsigned(28852,16),
    to_unsigned(28861,16),
    to_unsigned(28871,16),
    to_unsigned(28881,16),
    to_unsigned(28891,16),
    to_unsigned(28900,16),
    to_unsigned(28910,16),
    to_unsigned(28920,16),
    to_unsigned(28929,16),
    to_unsigned(28939,16),
    to_unsigned(28949,16),
    to_unsigned(28958,16),
    to_unsigned(28968,16),
    to_unsigned(28978,16),
    to_unsigned(28987,16),
    to_unsigned(28997,16),
    to_unsigned(29006,16),
    to_unsigned(29016,16),
    to_unsigned(29026,16),
    to_unsigned(29035,16),
    to_unsigned(29045,16),
    to_unsigned(29054,16),
    to_unsigned(29064,16),
    to_unsigned(29073,16),
    to_unsigned(29083,16),
    to_unsigned(29092,16),
    to_unsigned(29102,16),
    to_unsigned(29111,16),
    to_unsigned(29120,16),
    to_unsigned(29130,16),
    to_unsigned(29139,16),
    to_unsigned(29149,16),
    to_unsigned(29158,16),
    to_unsigned(29168,16),
    to_unsigned(29177,16),
    to_unsigned(29186,16),
    to_unsigned(29196,16),
    to_unsigned(29205,16),
    to_unsigned(29214,16),
    to_unsigned(29224,16),
    to_unsigned(29233,16),
    to_unsigned(29242,16),
    to_unsigned(29251,16),
    to_unsigned(29261,16),
    to_unsigned(29270,16),
    to_unsigned(29279,16),
    to_unsigned(29289,16),
    to_unsigned(29298,16),
    to_unsigned(29307,16),
    to_unsigned(29316,16),
    to_unsigned(29325,16),
    to_unsigned(29335,16),
    to_unsigned(29344,16),
    to_unsigned(29353,16),
    to_unsigned(29362,16),
    to_unsigned(29371,16),
    to_unsigned(29380,16),
    to_unsigned(29389,16),
    to_unsigned(29398,16),
    to_unsigned(29408,16),
    to_unsigned(29417,16),
    to_unsigned(29426,16),
    to_unsigned(29435,16),
    to_unsigned(29444,16),
    to_unsigned(29453,16),
    to_unsigned(29462,16),
    to_unsigned(29471,16),
    to_unsigned(29480,16),
    to_unsigned(29489,16),
    to_unsigned(29498,16),
    to_unsigned(29507,16),
    to_unsigned(29516,16),
    to_unsigned(29525,16),
    to_unsigned(29534,16),
    to_unsigned(29542,16),
    to_unsigned(29551,16),
    to_unsigned(29560,16),
    to_unsigned(29569,16),
    to_unsigned(29578,16),
    to_unsigned(29587,16),
    to_unsigned(29596,16),
    to_unsigned(29604,16),
    to_unsigned(29613,16),
    to_unsigned(29622,16),
    to_unsigned(29631,16),
    to_unsigned(29640,16),
    to_unsigned(29648,16),
    to_unsigned(29657,16),
    to_unsigned(29666,16),
    to_unsigned(29675,16),
    to_unsigned(29683,16),
    to_unsigned(29692,16),
    to_unsigned(29701,16),
    to_unsigned(29710,16),
    to_unsigned(29718,16),
    to_unsigned(29727,16),
    to_unsigned(29736,16),
    to_unsigned(29744,16),
    to_unsigned(29753,16),
    to_unsigned(29761,16),
    to_unsigned(29770,16),
    to_unsigned(29779,16),
    to_unsigned(29787,16),
    to_unsigned(29796,16),
    to_unsigned(29804,16),
    to_unsigned(29813,16),
    to_unsigned(29821,16),
    to_unsigned(29830,16),
    to_unsigned(29838,16),
    to_unsigned(29847,16),
    to_unsigned(29855,16),
    to_unsigned(29864,16),
    to_unsigned(29872,16),
    to_unsigned(29881,16),
    to_unsigned(29889,16),
    to_unsigned(29898,16),
    to_unsigned(29906,16),
    to_unsigned(29915,16),
    to_unsigned(29923,16),
    to_unsigned(29931,16),
    to_unsigned(29940,16),
    to_unsigned(29948,16),
    to_unsigned(29956,16),
    to_unsigned(29965,16),
    to_unsigned(29973,16),
    to_unsigned(29981,16),
    to_unsigned(29990,16),
    to_unsigned(29998,16),
    to_unsigned(30006,16),
    to_unsigned(30015,16),
    to_unsigned(30023,16),
    to_unsigned(30031,16),
    to_unsigned(30039,16),
    to_unsigned(30047,16),
    to_unsigned(30056,16),
    to_unsigned(30064,16),
    to_unsigned(30072,16),
    to_unsigned(30080,16),
    to_unsigned(30088,16),
    to_unsigned(30097,16),
    to_unsigned(30105,16),
    to_unsigned(30113,16),
    to_unsigned(30121,16),
    to_unsigned(30129,16),
    to_unsigned(30137,16),
    to_unsigned(30145,16),
    to_unsigned(30153,16),
    to_unsigned(30161,16),
    to_unsigned(30169,16),
    to_unsigned(30177,16),
    to_unsigned(30185,16),
    to_unsigned(30193,16),
    to_unsigned(30201,16),
    to_unsigned(30209,16),
    to_unsigned(30217,16),
    to_unsigned(30225,16),
    to_unsigned(30233,16),
    to_unsigned(30241,16),
    to_unsigned(30249,16),
    to_unsigned(30257,16),
    to_unsigned(30265,16),
    to_unsigned(30273,16),
    to_unsigned(30281,16),
    to_unsigned(30288,16),
    to_unsigned(30296,16),
    to_unsigned(30304,16),
    to_unsigned(30312,16),
    to_unsigned(30320,16),
    to_unsigned(30328,16),
    to_unsigned(30335,16),
    to_unsigned(30343,16),
    to_unsigned(30351,16),
    to_unsigned(30359,16),
    to_unsigned(30366,16),
    to_unsigned(30374,16),
    to_unsigned(30382,16),
    to_unsigned(30390,16),
    to_unsigned(30397,16),
    to_unsigned(30405,16),
    to_unsigned(30413,16),
    to_unsigned(30420,16),
    to_unsigned(30428,16),
    to_unsigned(30436,16),
    to_unsigned(30443,16),
    to_unsigned(30451,16),
    to_unsigned(30458,16),
    to_unsigned(30466,16),
    to_unsigned(30474,16),
    to_unsigned(30481,16),
    to_unsigned(30489,16),
    to_unsigned(30496,16),
    to_unsigned(30504,16),
    to_unsigned(30511,16),
    to_unsigned(30519,16),
    to_unsigned(30526,16),
    to_unsigned(30534,16),
    to_unsigned(30541,16),
    to_unsigned(30549,16),
    to_unsigned(30556,16),
    to_unsigned(30563,16),
    to_unsigned(30571,16),
    to_unsigned(30578,16),
    to_unsigned(30586,16),
    to_unsigned(30593,16),
    to_unsigned(30600,16),
    to_unsigned(30608,16),
    to_unsigned(30615,16),
    to_unsigned(30622,16),
    to_unsigned(30630,16),
    to_unsigned(30637,16),
    to_unsigned(30644,16),
    to_unsigned(30652,16),
    to_unsigned(30659,16),
    to_unsigned(30666,16),
    to_unsigned(30673,16),
    to_unsigned(30681,16),
    to_unsigned(30688,16),
    to_unsigned(30695,16),
    to_unsigned(30702,16),
    to_unsigned(30710,16),
    to_unsigned(30717,16),
    to_unsigned(30724,16),
    to_unsigned(30731,16),
    to_unsigned(30738,16),
    to_unsigned(30745,16),
    to_unsigned(30752,16),
    to_unsigned(30759,16),
    to_unsigned(30767,16),
    to_unsigned(30774,16),
    to_unsigned(30781,16),
    to_unsigned(30788,16),
    to_unsigned(30795,16),
    to_unsigned(30802,16),
    to_unsigned(30809,16),
    to_unsigned(30816,16),
    to_unsigned(30823,16),
    to_unsigned(30830,16),
    to_unsigned(30837,16),
    to_unsigned(30844,16),
    to_unsigned(30851,16),
    to_unsigned(30858,16),
    to_unsigned(30865,16),
    to_unsigned(30871,16),
    to_unsigned(30878,16),
    to_unsigned(30885,16),
    to_unsigned(30892,16),
    to_unsigned(30899,16),
    to_unsigned(30906,16),
    to_unsigned(30913,16),
    to_unsigned(30919,16),
    to_unsigned(30926,16),
    to_unsigned(30933,16),
    to_unsigned(30940,16),
    to_unsigned(30947,16),
    to_unsigned(30953,16),
    to_unsigned(30960,16),
    to_unsigned(30967,16),
    to_unsigned(30974,16),
    to_unsigned(30980,16),
    to_unsigned(30987,16),
    to_unsigned(30994,16),
    to_unsigned(31000,16),
    to_unsigned(31007,16),
    to_unsigned(31014,16),
    to_unsigned(31020,16),
    to_unsigned(31027,16),
    to_unsigned(31034,16),
    to_unsigned(31040,16),
    to_unsigned(31047,16),
    to_unsigned(31053,16),
    to_unsigned(31060,16),
    to_unsigned(31066,16),
    to_unsigned(31073,16),
    to_unsigned(31080,16),
    to_unsigned(31086,16),
    to_unsigned(31093,16),
    to_unsigned(31099,16),
    to_unsigned(31106,16),
    to_unsigned(31112,16),
    to_unsigned(31118,16),
    to_unsigned(31125,16),
    to_unsigned(31131,16),
    to_unsigned(31138,16),
    to_unsigned(31144,16),
    to_unsigned(31151,16),
    to_unsigned(31157,16),
    to_unsigned(31163,16),
    to_unsigned(31170,16),
    to_unsigned(31176,16),
    to_unsigned(31182,16),
    to_unsigned(31189,16),
    to_unsigned(31195,16),
    to_unsigned(31201,16),
    to_unsigned(31208,16),
    to_unsigned(31214,16),
    to_unsigned(31220,16),
    to_unsigned(31226,16),
    to_unsigned(31233,16),
    to_unsigned(31239,16),
    to_unsigned(31245,16),
    to_unsigned(31251,16),
    to_unsigned(31257,16),
    to_unsigned(31263,16),
    to_unsigned(31270,16),
    to_unsigned(31276,16),
    to_unsigned(31282,16),
    to_unsigned(31288,16),
    to_unsigned(31294,16),
    to_unsigned(31300,16),
    to_unsigned(31306,16),
    to_unsigned(31312,16),
    to_unsigned(31318,16),
    to_unsigned(31325,16),
    to_unsigned(31331,16),
    to_unsigned(31337,16),
    to_unsigned(31343,16),
    to_unsigned(31349,16),
    to_unsigned(31355,16),
    to_unsigned(31361,16),
    to_unsigned(31367,16),
    to_unsigned(31372,16),
    to_unsigned(31378,16),
    to_unsigned(31384,16),
    to_unsigned(31390,16),
    to_unsigned(31396,16),
    to_unsigned(31402,16),
    to_unsigned(31408,16),
    to_unsigned(31414,16),
    to_unsigned(31420,16),
    to_unsigned(31425,16),
    to_unsigned(31431,16),
    to_unsigned(31437,16),
    to_unsigned(31443,16),
    to_unsigned(31449,16),
    to_unsigned(31454,16),
    to_unsigned(31460,16),
    to_unsigned(31466,16),
    to_unsigned(31472,16),
    to_unsigned(31477,16),
    to_unsigned(31483,16),
    to_unsigned(31489,16),
    to_unsigned(31495,16),
    to_unsigned(31500,16),
    to_unsigned(31506,16),
    to_unsigned(31511,16),
    to_unsigned(31517,16),
    to_unsigned(31523,16),
    to_unsigned(31528,16),
    to_unsigned(31534,16),
    to_unsigned(31540,16),
    to_unsigned(31545,16),
    to_unsigned(31551,16),
    to_unsigned(31556,16),
    to_unsigned(31562,16),
    to_unsigned(31567,16),
    to_unsigned(31573,16),
    to_unsigned(31578,16),
    to_unsigned(31584,16),
    to_unsigned(31589,16),
    to_unsigned(31595,16),
    to_unsigned(31600,16),
    to_unsigned(31606,16),
    to_unsigned(31611,16),
    to_unsigned(31616,16),
    to_unsigned(31622,16),
    to_unsigned(31627,16),
    to_unsigned(31633,16),
    to_unsigned(31638,16),
    to_unsigned(31643,16),
    to_unsigned(31649,16),
    to_unsigned(31654,16),
    to_unsigned(31659,16),
    to_unsigned(31665,16),
    to_unsigned(31670,16),
    to_unsigned(31675,16),
    to_unsigned(31680,16),
    to_unsigned(31686,16),
    to_unsigned(31691,16),
    to_unsigned(31696,16),
    to_unsigned(31701,16),
    to_unsigned(31707,16),
    to_unsigned(31712,16),
    to_unsigned(31717,16),
    to_unsigned(31722,16),
    to_unsigned(31727,16),
    to_unsigned(31732,16),
    to_unsigned(31738,16),
    to_unsigned(31743,16),
    to_unsigned(31748,16),
    to_unsigned(31753,16),
    to_unsigned(31758,16),
    to_unsigned(31763,16),
    to_unsigned(31768,16),
    to_unsigned(31773,16),
    to_unsigned(31778,16),
    to_unsigned(31783,16),
    to_unsigned(31788,16),
    to_unsigned(31793,16),
    to_unsigned(31798,16),
    to_unsigned(31803,16),
    to_unsigned(31808,16),
    to_unsigned(31813,16),
    to_unsigned(31818,16),
    to_unsigned(31823,16),
    to_unsigned(31828,16),
    to_unsigned(31833,16),
    to_unsigned(31837,16),
    to_unsigned(31842,16),
    to_unsigned(31847,16),
    to_unsigned(31852,16),
    to_unsigned(31857,16),
    to_unsigned(31862,16),
    to_unsigned(31866,16),
    to_unsigned(31871,16),
    to_unsigned(31876,16),
    to_unsigned(31881,16),
    to_unsigned(31886,16),
    to_unsigned(31890,16),
    to_unsigned(31895,16),
    to_unsigned(31900,16),
    to_unsigned(31904,16),
    to_unsigned(31909,16),
    to_unsigned(31914,16),
    to_unsigned(31918,16),
    to_unsigned(31923,16),
    to_unsigned(31928,16),
    to_unsigned(31932,16),
    to_unsigned(31937,16),
    to_unsigned(31942,16),
    to_unsigned(31946,16),
    to_unsigned(31951,16),
    to_unsigned(31955,16),
    to_unsigned(31960,16),
    to_unsigned(31964,16),
    to_unsigned(31969,16),
    to_unsigned(31973,16),
    to_unsigned(31978,16),
    to_unsigned(31982,16),
    to_unsigned(31987,16),
    to_unsigned(31991,16),
    to_unsigned(31996,16),
    to_unsigned(32000,16),
    to_unsigned(32005,16),
    to_unsigned(32009,16),
    to_unsigned(32013,16),
    to_unsigned(32018,16),
    to_unsigned(32022,16),
    to_unsigned(32027,16),
    to_unsigned(32031,16),
    to_unsigned(32035,16),
    to_unsigned(32040,16),
    to_unsigned(32044,16),
    to_unsigned(32048,16),
    to_unsigned(32052,16),
    to_unsigned(32057,16),
    to_unsigned(32061,16),
    to_unsigned(32065,16),
    to_unsigned(32069,16),
    to_unsigned(32074,16),
    to_unsigned(32078,16),
    to_unsigned(32082,16),
    to_unsigned(32086,16),
    to_unsigned(32090,16),
    to_unsigned(32095,16),
    to_unsigned(32099,16),
    to_unsigned(32103,16),
    to_unsigned(32107,16),
    to_unsigned(32111,16),
    to_unsigned(32115,16),
    to_unsigned(32119,16),
    to_unsigned(32123,16),
    to_unsigned(32127,16),
    to_unsigned(32131,16),
    to_unsigned(32135,16),
    to_unsigned(32139,16),
    to_unsigned(32143,16),
    to_unsigned(32147,16),
    to_unsigned(32151,16),
    to_unsigned(32155,16),
    to_unsigned(32159,16),
    to_unsigned(32163,16),
    to_unsigned(32167,16),
    to_unsigned(32171,16),
    to_unsigned(32175,16),
    to_unsigned(32179,16),
    to_unsigned(32183,16),
    to_unsigned(32187,16),
    to_unsigned(32190,16),
    to_unsigned(32194,16),
    to_unsigned(32198,16),
    to_unsigned(32202,16),
    to_unsigned(32206,16),
    to_unsigned(32210,16),
    to_unsigned(32213,16),
    to_unsigned(32217,16),
    to_unsigned(32221,16),
    to_unsigned(32225,16),
    to_unsigned(32228,16),
    to_unsigned(32232,16),
    to_unsigned(32236,16),
    to_unsigned(32239,16),
    to_unsigned(32243,16),
    to_unsigned(32247,16),
    to_unsigned(32250,16),
    to_unsigned(32254,16),
    to_unsigned(32258,16),
    to_unsigned(32261,16),
    to_unsigned(32265,16),
    to_unsigned(32268,16),
    to_unsigned(32272,16),
    to_unsigned(32276,16),
    to_unsigned(32279,16),
    to_unsigned(32283,16),
    to_unsigned(32286,16),
    to_unsigned(32290,16),
    to_unsigned(32293,16),
    to_unsigned(32297,16),
    to_unsigned(32300,16),
    to_unsigned(32304,16),
    to_unsigned(32307,16),
    to_unsigned(32310,16),
    to_unsigned(32314,16),
    to_unsigned(32317,16),
    to_unsigned(32321,16),
    to_unsigned(32324,16),
    to_unsigned(32327,16),
    to_unsigned(32331,16),
    to_unsigned(32334,16),
    to_unsigned(32337,16),
    to_unsigned(32341,16),
    to_unsigned(32344,16),
    to_unsigned(32347,16),
    to_unsigned(32351,16),
    to_unsigned(32354,16),
    to_unsigned(32357,16),
    to_unsigned(32360,16),
    to_unsigned(32364,16),
    to_unsigned(32367,16),
    to_unsigned(32370,16),
    to_unsigned(32373,16),
    to_unsigned(32376,16),
    to_unsigned(32380,16),
    to_unsigned(32383,16),
    to_unsigned(32386,16),
    to_unsigned(32389,16),
    to_unsigned(32392,16),
    to_unsigned(32395,16),
    to_unsigned(32398,16),
    to_unsigned(32401,16),
    to_unsigned(32404,16),
    to_unsigned(32407,16),
    to_unsigned(32410,16),
    to_unsigned(32413,16),
    to_unsigned(32416,16),
    to_unsigned(32419,16),
    to_unsigned(32422,16),
    to_unsigned(32425,16),
    to_unsigned(32428,16),
    to_unsigned(32431,16),
    to_unsigned(32434,16),
    to_unsigned(32437,16),
    to_unsigned(32440,16),
    to_unsigned(32443,16),
    to_unsigned(32446,16),
    to_unsigned(32449,16),
    to_unsigned(32452,16),
    to_unsigned(32454,16),
    to_unsigned(32457,16),
    to_unsigned(32460,16),
    to_unsigned(32463,16),
    to_unsigned(32466,16),
    to_unsigned(32468,16),
    to_unsigned(32471,16),
    to_unsigned(32474,16),
    to_unsigned(32477,16),
    to_unsigned(32479,16),
    to_unsigned(32482,16),
    to_unsigned(32485,16),
    to_unsigned(32488,16),
    to_unsigned(32490,16),
    to_unsigned(32493,16),
    to_unsigned(32496,16),
    to_unsigned(32498,16),
    to_unsigned(32501,16),
    to_unsigned(32503,16),
    to_unsigned(32506,16),
    to_unsigned(32509,16),
    to_unsigned(32511,16),
    to_unsigned(32514,16),
    to_unsigned(32516,16),
    to_unsigned(32519,16),
    to_unsigned(32521,16),
    to_unsigned(32524,16),
    to_unsigned(32526,16),
    to_unsigned(32529,16),
    to_unsigned(32531,16),
    to_unsigned(32534,16),
    to_unsigned(32536,16),
    to_unsigned(32539,16),
    to_unsigned(32541,16),
    to_unsigned(32543,16),
    to_unsigned(32546,16),
    to_unsigned(32548,16),
    to_unsigned(32551,16),
    to_unsigned(32553,16),
    to_unsigned(32555,16),
    to_unsigned(32558,16),
    to_unsigned(32560,16),
    to_unsigned(32562,16),
    to_unsigned(32565,16),
    to_unsigned(32567,16),
    to_unsigned(32569,16),
    to_unsigned(32571,16),
    to_unsigned(32574,16),
    to_unsigned(32576,16),
    to_unsigned(32578,16),
    to_unsigned(32580,16),
    to_unsigned(32582,16),
    to_unsigned(32585,16),
    to_unsigned(32587,16),
    to_unsigned(32589,16),
    to_unsigned(32591,16),
    to_unsigned(32593,16),
    to_unsigned(32595,16),
    to_unsigned(32597,16),
    to_unsigned(32599,16),
    to_unsigned(32602,16),
    to_unsigned(32604,16),
    to_unsigned(32606,16),
    to_unsigned(32608,16),
    to_unsigned(32610,16),
    to_unsigned(32612,16),
    to_unsigned(32614,16),
    to_unsigned(32616,16),
    to_unsigned(32618,16),
    to_unsigned(32620,16),
    to_unsigned(32622,16),
    to_unsigned(32624,16),
    to_unsigned(32625,16),
    to_unsigned(32627,16),
    to_unsigned(32629,16),
    to_unsigned(32631,16),
    to_unsigned(32633,16),
    to_unsigned(32635,16),
    to_unsigned(32637,16),
    to_unsigned(32638,16),
    to_unsigned(32640,16),
    to_unsigned(32642,16),
    to_unsigned(32644,16),
    to_unsigned(32646,16),
    to_unsigned(32647,16),
    to_unsigned(32649,16),
    to_unsigned(32651,16),
    to_unsigned(32653,16),
    to_unsigned(32654,16),
    to_unsigned(32656,16),
    to_unsigned(32658,16),
    to_unsigned(32659,16),
    to_unsigned(32661,16),
    to_unsigned(32663,16),
    to_unsigned(32664,16),
    to_unsigned(32666,16),
    to_unsigned(32668,16),
    to_unsigned(32669,16),
    to_unsigned(32671,16),
    to_unsigned(32672,16),
    to_unsigned(32674,16),
    to_unsigned(32675,16),
    to_unsigned(32677,16),
    to_unsigned(32679,16),
    to_unsigned(32680,16),
    to_unsigned(32681,16),
    to_unsigned(32683,16),
    to_unsigned(32684,16),
    to_unsigned(32686,16),
    to_unsigned(32687,16),
    to_unsigned(32689,16),
    to_unsigned(32690,16),
    to_unsigned(32692,16),
    to_unsigned(32693,16),
    to_unsigned(32694,16),
    to_unsigned(32696,16),
    to_unsigned(32697,16),
    to_unsigned(32698,16),
    to_unsigned(32700,16),
    to_unsigned(32701,16),
    to_unsigned(32702,16),
    to_unsigned(32704,16),
    to_unsigned(32705,16),
    to_unsigned(32706,16),
    to_unsigned(32707,16),
    to_unsigned(32709,16),
    to_unsigned(32710,16),
    to_unsigned(32711,16),
    to_unsigned(32712,16),
    to_unsigned(32713,16),
    to_unsigned(32715,16),
    to_unsigned(32716,16),
    to_unsigned(32717,16),
    to_unsigned(32718,16),
    to_unsigned(32719,16),
    to_unsigned(32720,16),
    to_unsigned(32721,16),
    to_unsigned(32722,16),
    to_unsigned(32724,16),
    to_unsigned(32725,16),
    to_unsigned(32726,16),
    to_unsigned(32727,16),
    to_unsigned(32728,16),
    to_unsigned(32729,16),
    to_unsigned(32730,16),
    to_unsigned(32731,16),
    to_unsigned(32732,16),
    to_unsigned(32733,16),
    to_unsigned(32733,16),
    to_unsigned(32734,16),
    to_unsigned(32735,16),
    to_unsigned(32736,16),
    to_unsigned(32737,16),
    to_unsigned(32738,16),
    to_unsigned(32739,16),
    to_unsigned(32740,16),
    to_unsigned(32741,16),
    to_unsigned(32741,16),
    to_unsigned(32742,16),
    to_unsigned(32743,16),
    to_unsigned(32744,16),
    to_unsigned(32744,16),
    to_unsigned(32745,16),
    to_unsigned(32746,16),
    to_unsigned(32747,16),
    to_unsigned(32747,16),
    to_unsigned(32748,16),
    to_unsigned(32749,16),
    to_unsigned(32750,16),
    to_unsigned(32750,16),
    to_unsigned(32751,16),
    to_unsigned(32751,16),
    to_unsigned(32752,16),
    to_unsigned(32753,16),
    to_unsigned(32753,16),
    to_unsigned(32754,16),
    to_unsigned(32754,16),
    to_unsigned(32755,16),
    to_unsigned(32756,16),
    to_unsigned(32756,16),
    to_unsigned(32757,16),
    to_unsigned(32757,16),
    to_unsigned(32758,16),
    to_unsigned(32758,16),
    to_unsigned(32759,16),
    to_unsigned(32759,16),
    to_unsigned(32760,16),
    to_unsigned(32760,16),
    to_unsigned(32760,16),
    to_unsigned(32761,16),
    to_unsigned(32761,16),
    to_unsigned(32762,16),
    to_unsigned(32762,16),
    to_unsigned(32762,16),
    to_unsigned(32763,16),
    to_unsigned(32763,16),
    to_unsigned(32763,16),
    to_unsigned(32764,16),
    to_unsigned(32764,16),
    to_unsigned(32764,16),
    to_unsigned(32764,16),
    to_unsigned(32765,16),
    to_unsigned(32765,16),
    to_unsigned(32765,16),
    to_unsigned(32765,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32766,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16),
    to_unsigned(32767,16)
	);


-- Quarter sine lookup table
type lut_65536_x_32_type is array(0 to 16383) of unsigned(31 downto 0);

constant sine_lut_65536_x_32 : lut_65536_x_32_type := (
    to_unsigned(0,32),
    to_unsigned(205887,32),
    to_unsigned(411775,32),
    to_unsigned(617662,32),
    to_unsigned(823550,32),
    to_unsigned(1029437,32),
    to_unsigned(1235324,32),
    to_unsigned(1441212,32),
    to_unsigned(1647099,32),
    to_unsigned(1852987,32),
    to_unsigned(2058874,32),
    to_unsigned(2264761,32),
    to_unsigned(2470648,32),
    to_unsigned(2676536,32),
    to_unsigned(2882423,32),
    to_unsigned(3088310,32),
    to_unsigned(3294197,32),
    to_unsigned(3500085,32),
    to_unsigned(3705972,32),
    to_unsigned(3911859,32),
    to_unsigned(4117746,32),
    to_unsigned(4323633,32),
    to_unsigned(4529520,32),
    to_unsigned(4735407,32),
    to_unsigned(4941294,32),
    to_unsigned(5147180,32),
    to_unsigned(5353067,32),
    to_unsigned(5558954,32),
    to_unsigned(5764841,32),
    to_unsigned(5970727,32),
    to_unsigned(6176614,32),
    to_unsigned(6382501,32),
    to_unsigned(6588387,32),
    to_unsigned(6794273,32),
    to_unsigned(7000160,32),
    to_unsigned(7206046,32),
    to_unsigned(7411932,32),
    to_unsigned(7617818,32),
    to_unsigned(7823705,32),
    to_unsigned(8029591,32),
    to_unsigned(8235476,32),
    to_unsigned(8441362,32),
    to_unsigned(8647248,32),
    to_unsigned(8853134,32),
    to_unsigned(9059019,32),
    to_unsigned(9264905,32),
    to_unsigned(9470790,32),
    to_unsigned(9676676,32),
    to_unsigned(9882561,32),
    to_unsigned(10088446,32),
    to_unsigned(10294331,32),
    to_unsigned(10500216,32),
    to_unsigned(10706101,32),
    to_unsigned(10911986,32),
    to_unsigned(11117871,32),
    to_unsigned(11323755,32),
    to_unsigned(11529640,32),
    to_unsigned(11735524,32),
    to_unsigned(11941409,32),
    to_unsigned(12147293,32),
    to_unsigned(12353177,32),
    to_unsigned(12559061,32),
    to_unsigned(12764945,32),
    to_unsigned(12970828,32),
    to_unsigned(13176712,32),
    to_unsigned(13382595,32),
    to_unsigned(13588479,32),
    to_unsigned(13794362,32),
    to_unsigned(14000245,32),
    to_unsigned(14206128,32),
    to_unsigned(14412011,32),
    to_unsigned(14617894,32),
    to_unsigned(14823776,32),
    to_unsigned(15029659,32),
    to_unsigned(15235541,32),
    to_unsigned(15441423,32),
    to_unsigned(15647305,32),
    to_unsigned(15853187,32),
    to_unsigned(16059069,32),
    to_unsigned(16264950,32),
    to_unsigned(16470832,32),
    to_unsigned(16676713,32),
    to_unsigned(16882594,32),
    to_unsigned(17088475,32),
    to_unsigned(17294356,32),
    to_unsigned(17500237,32),
    to_unsigned(17706117,32),
    to_unsigned(17911997,32),
    to_unsigned(18117878,32),
    to_unsigned(18323758,32),
    to_unsigned(18529638,32),
    to_unsigned(18735517,32),
    to_unsigned(18941397,32),
    to_unsigned(19147276,32),
    to_unsigned(19353155,32),
    to_unsigned(19559034,32),
    to_unsigned(19764913,32),
    to_unsigned(19970791,32),
    to_unsigned(20176670,32),
    to_unsigned(20382548,32),
    to_unsigned(20588426,32),
    to_unsigned(20794304,32),
    to_unsigned(21000182,32),
    to_unsigned(21206059,32),
    to_unsigned(21411936,32),
    to_unsigned(21617814,32),
    to_unsigned(21823690,32),
    to_unsigned(22029567,32),
    to_unsigned(22235444,32),
    to_unsigned(22441320,32),
    to_unsigned(22647196,32),
    to_unsigned(22853072,32),
    to_unsigned(23058947,32),
    to_unsigned(23264823,32),
    to_unsigned(23470698,32),
    to_unsigned(23676573,32),
    to_unsigned(23882448,32),
    to_unsigned(24088323,32),
    to_unsigned(24294197,32),
    to_unsigned(24500071,32),
    to_unsigned(24705945,32),
    to_unsigned(24911819,32),
    to_unsigned(25117692,32),
    to_unsigned(25323565,32),
    to_unsigned(25529438,32),
    to_unsigned(25735311,32),
    to_unsigned(25941183,32),
    to_unsigned(26147056,32),
    to_unsigned(26352928,32),
    to_unsigned(26558800,32),
    to_unsigned(26764671,32),
    to_unsigned(26970542,32),
    to_unsigned(27176413,32),
    to_unsigned(27382284,32),
    to_unsigned(27588155,32),
    to_unsigned(27794025,32),
    to_unsigned(27999895,32),
    to_unsigned(28205765,32),
    to_unsigned(28411634,32),
    to_unsigned(28617504,32),
    to_unsigned(28823373,32),
    to_unsigned(29029242,32),
    to_unsigned(29235110,32),
    to_unsigned(29440978,32),
    to_unsigned(29646846,32),
    to_unsigned(29852714,32),
    to_unsigned(30058581,32),
    to_unsigned(30264448,32),
    to_unsigned(30470315,32),
    to_unsigned(30676182,32),
    to_unsigned(30882048,32),
    to_unsigned(31087914,32),
    to_unsigned(31293780,32),
    to_unsigned(31499645,32),
    to_unsigned(31705510,32),
    to_unsigned(31911375,32),
    to_unsigned(32117239,32),
    to_unsigned(32323104,32),
    to_unsigned(32528968,32),
    to_unsigned(32734831,32),
    to_unsigned(32940695,32),
    to_unsigned(33146558,32),
    to_unsigned(33352420,32),
    to_unsigned(33558283,32),
    to_unsigned(33764145,32),
    to_unsigned(33970007,32),
    to_unsigned(34175868,32),
    to_unsigned(34381729,32),
    to_unsigned(34587590,32),
    to_unsigned(34793451,32),
    to_unsigned(34999311,32),
    to_unsigned(35205171,32),
    to_unsigned(35411031,32),
    to_unsigned(35616890,32),
    to_unsigned(35822749,32),
    to_unsigned(36028607,32),
    to_unsigned(36234466,32),
    to_unsigned(36440324,32),
    to_unsigned(36646181,32),
    to_unsigned(36852039,32),
    to_unsigned(37057895,32),
    to_unsigned(37263752,32),
    to_unsigned(37469608,32),
    to_unsigned(37675464,32),
    to_unsigned(37881320,32),
    to_unsigned(38087175,32),
    to_unsigned(38293030,32),
    to_unsigned(38498884,32),
    to_unsigned(38704738,32),
    to_unsigned(38910592,32),
    to_unsigned(39116446,32),
    to_unsigned(39322299,32),
    to_unsigned(39528151,32),
    to_unsigned(39734004,32),
    to_unsigned(39939856,32),
    to_unsigned(40145707,32),
    to_unsigned(40351559,32),
    to_unsigned(40557410,32),
    to_unsigned(40763260,32),
    to_unsigned(40969110,32),
    to_unsigned(41174960,32),
    to_unsigned(41380809,32),
    to_unsigned(41586658,32),
    to_unsigned(41792507,32),
    to_unsigned(41998355,32),
    to_unsigned(42204203,32),
    to_unsigned(42410050,32),
    to_unsigned(42615898,32),
    to_unsigned(42821744,32),
    to_unsigned(43027591,32),
    to_unsigned(43233436,32),
    to_unsigned(43439282,32),
    to_unsigned(43645127,32),
    to_unsigned(43850972,32),
    to_unsigned(44056816,32),
    to_unsigned(44262660,32),
    to_unsigned(44468503,32),
    to_unsigned(44674346,32),
    to_unsigned(44880189,32),
    to_unsigned(45086031,32),
    to_unsigned(45291873,32),
    to_unsigned(45497715,32),
    to_unsigned(45703556,32),
    to_unsigned(45909396,32),
    to_unsigned(46115236,32),
    to_unsigned(46321076,32),
    to_unsigned(46526915,32),
    to_unsigned(46732754,32),
    to_unsigned(46938593,32),
    to_unsigned(47144431,32),
    to_unsigned(47350268,32),
    to_unsigned(47556105,32),
    to_unsigned(47761942,32),
    to_unsigned(47967778,32),
    to_unsigned(48173614,32),
    to_unsigned(48379449,32),
    to_unsigned(48585284,32),
    to_unsigned(48791119,32),
    to_unsigned(48996953,32),
    to_unsigned(49202787,32),
    to_unsigned(49408620,32),
    to_unsigned(49614452,32),
    to_unsigned(49820285,32),
    to_unsigned(50026116,32),
    to_unsigned(50231948,32),
    to_unsigned(50437779,32),
    to_unsigned(50643609,32),
    to_unsigned(50849439,32),
    to_unsigned(51055268,32),
    to_unsigned(51261097,32),
    to_unsigned(51466926,32),
    to_unsigned(51672754,32),
    to_unsigned(51878581,32),
    to_unsigned(52084409,32),
    to_unsigned(52290235,32),
    to_unsigned(52496061,32),
    to_unsigned(52701887,32),
    to_unsigned(52907712,32),
    to_unsigned(53113537,32),
    to_unsigned(53319361,32),
    to_unsigned(53525185,32),
    to_unsigned(53731008,32),
    to_unsigned(53936831,32),
    to_unsigned(54142653,32),
    to_unsigned(54348475,32),
    to_unsigned(54554296,32),
    to_unsigned(54760116,32),
    to_unsigned(54965937,32),
    to_unsigned(55171756,32),
    to_unsigned(55377576,32),
    to_unsigned(55583394,32),
    to_unsigned(55789212,32),
    to_unsigned(55995030,32),
    to_unsigned(56200847,32),
    to_unsigned(56406664,32),
    to_unsigned(56612480,32),
    to_unsigned(56818296,32),
    to_unsigned(57024111,32),
    to_unsigned(57229925,32),
    to_unsigned(57435739,32),
    to_unsigned(57641553,32),
    to_unsigned(57847366,32),
    to_unsigned(58053178,32),
    to_unsigned(58258990,32),
    to_unsigned(58464801,32),
    to_unsigned(58670612,32),
    to_unsigned(58876423,32),
    to_unsigned(59082232,32),
    to_unsigned(59288042,32),
    to_unsigned(59493850,32),
    to_unsigned(59699658,32),
    to_unsigned(59905466,32),
    to_unsigned(60111273,32),
    to_unsigned(60317079,32),
    to_unsigned(60522885,32),
    to_unsigned(60728691,32),
    to_unsigned(60934495,32),
    to_unsigned(61140300,32),
    to_unsigned(61346103,32),
    to_unsigned(61551906,32),
    to_unsigned(61757709,32),
    to_unsigned(61963511,32),
    to_unsigned(62169312,32),
    to_unsigned(62375113,32),
    to_unsigned(62580914,32),
    to_unsigned(62786713,32),
    to_unsigned(62992512,32),
    to_unsigned(63198311,32),
    to_unsigned(63404109,32),
    to_unsigned(63609906,32),
    to_unsigned(63815703,32),
    to_unsigned(64021499,32),
    to_unsigned(64227295,32),
    to_unsigned(64433090,32),
    to_unsigned(64638884,32),
    to_unsigned(64844678,32),
    to_unsigned(65050471,32),
    to_unsigned(65256264,32),
    to_unsigned(65462056,32),
    to_unsigned(65667847,32),
    to_unsigned(65873638,32),
    to_unsigned(66079428,32),
    to_unsigned(66285218,32),
    to_unsigned(66491007,32),
    to_unsigned(66696795,32),
    to_unsigned(66902583,32),
    to_unsigned(67108370,32),
    to_unsigned(67314157,32),
    to_unsigned(67519943,32),
    to_unsigned(67725728,32),
    to_unsigned(67931513,32),
    to_unsigned(68137297,32),
    to_unsigned(68343080,32),
    to_unsigned(68548863,32),
    to_unsigned(68754645,32),
    to_unsigned(68960427,32),
    to_unsigned(69166208,32),
    to_unsigned(69371988,32),
    to_unsigned(69577768,32),
    to_unsigned(69783547,32),
    to_unsigned(69989325,32),
    to_unsigned(70195103,32),
    to_unsigned(70400880,32),
    to_unsigned(70606656,32),
    to_unsigned(70812432,32),
    to_unsigned(71018207,32),
    to_unsigned(71223982,32),
    to_unsigned(71429756,32),
    to_unsigned(71635529,32),
    to_unsigned(71841301,32),
    to_unsigned(72047073,32),
    to_unsigned(72252844,32),
    to_unsigned(72458615,32),
    to_unsigned(72664385,32),
    to_unsigned(72870154,32),
    to_unsigned(73075922,32),
    to_unsigned(73281690,32),
    to_unsigned(73487457,32),
    to_unsigned(73693224,32),
    to_unsigned(73898990,32),
    to_unsigned(74104755,32),
    to_unsigned(74310519,32),
    to_unsigned(74516283,32),
    to_unsigned(74722046,32),
    to_unsigned(74927808,32),
    to_unsigned(75133570,32),
    to_unsigned(75339331,32),
    to_unsigned(75545092,32),
    to_unsigned(75750851,32),
    to_unsigned(75956610,32),
    to_unsigned(76162368,32),
    to_unsigned(76368126,32),
    to_unsigned(76573883,32),
    to_unsigned(76779639,32),
    to_unsigned(76985394,32),
    to_unsigned(77191149,32),
    to_unsigned(77396903,32),
    to_unsigned(77602656,32),
    to_unsigned(77808409,32),
    to_unsigned(78014161,32),
    to_unsigned(78219912,32),
    to_unsigned(78425662,32),
    to_unsigned(78631412,32),
    to_unsigned(78837161,32),
    to_unsigned(79042909,32),
    to_unsigned(79248657,32),
    to_unsigned(79454404,32),
    to_unsigned(79660150,32),
    to_unsigned(79865895,32),
    to_unsigned(80071640,32),
    to_unsigned(80277384,32),
    to_unsigned(80483127,32),
    to_unsigned(80688869,32),
    to_unsigned(80894611,32),
    to_unsigned(81100352,32),
    to_unsigned(81306092,32),
    to_unsigned(81511831,32),
    to_unsigned(81717570,32),
    to_unsigned(81923308,32),
    to_unsigned(82129045,32),
    to_unsigned(82334782,32),
    to_unsigned(82540517,32),
    to_unsigned(82746252,32),
    to_unsigned(82951986,32),
    to_unsigned(83157720,32),
    to_unsigned(83363452,32),
    to_unsigned(83569184,32),
    to_unsigned(83774915,32),
    to_unsigned(83980645,32),
    to_unsigned(84186375,32),
    to_unsigned(84392104,32),
    to_unsigned(84597832,32),
    to_unsigned(84803559,32),
    to_unsigned(85009285,32),
    to_unsigned(85215011,32),
    to_unsigned(85420736,32),
    to_unsigned(85626460,32),
    to_unsigned(85832183,32),
    to_unsigned(86037906,32),
    to_unsigned(86243627,32),
    to_unsigned(86449348,32),
    to_unsigned(86655069,32),
    to_unsigned(86860788,32),
    to_unsigned(87066506,32),
    to_unsigned(87272224,32),
    to_unsigned(87477941,32),
    to_unsigned(87683657,32),
    to_unsigned(87889372,32),
    to_unsigned(88095087,32),
    to_unsigned(88300801,32),
    to_unsigned(88506514,32),
    to_unsigned(88712226,32),
    to_unsigned(88917937,32),
    to_unsigned(89123647,32),
    to_unsigned(89329357,32),
    to_unsigned(89535066,32),
    to_unsigned(89740774,32),
    to_unsigned(89946481,32),
    to_unsigned(90152187,32),
    to_unsigned(90357893,32),
    to_unsigned(90563597,32),
    to_unsigned(90769301,32),
    to_unsigned(90975004,32),
    to_unsigned(91180706,32),
    to_unsigned(91386408,32),
    to_unsigned(91592108,32),
    to_unsigned(91797808,32),
    to_unsigned(92003507,32),
    to_unsigned(92209205,32),
    to_unsigned(92414902,32),
    to_unsigned(92620598,32),
    to_unsigned(92826293,32),
    to_unsigned(93031988,32),
    to_unsigned(93237682,32),
    to_unsigned(93443374,32),
    to_unsigned(93649066,32),
    to_unsigned(93854758,32),
    to_unsigned(94060448,32),
    to_unsigned(94266137,32),
    to_unsigned(94471826,32),
    to_unsigned(94677513,32),
    to_unsigned(94883200,32),
    to_unsigned(95088886,32),
    to_unsigned(95294571,32),
    to_unsigned(95500255,32),
    to_unsigned(95705939,32),
    to_unsigned(95911621,32),
    to_unsigned(96117303,32),
    to_unsigned(96322983,32),
    to_unsigned(96528663,32),
    to_unsigned(96734342,32),
    to_unsigned(96940020,32),
    to_unsigned(97145697,32),
    to_unsigned(97351373,32),
    to_unsigned(97557048,32),
    to_unsigned(97762723,32),
    to_unsigned(97968396,32),
    to_unsigned(98174069,32),
    to_unsigned(98379741,32),
    to_unsigned(98585411,32),
    to_unsigned(98791081,32),
    to_unsigned(98996750,32),
    to_unsigned(99202418,32),
    to_unsigned(99408086,32),
    to_unsigned(99613752,32),
    to_unsigned(99819417,32),
    to_unsigned(100025082,32),
    to_unsigned(100230745,32),
    to_unsigned(100436408,32),
    to_unsigned(100642069,32),
    to_unsigned(100847730,32),
    to_unsigned(101053390,32),
    to_unsigned(101259049,32),
    to_unsigned(101464707,32),
    to_unsigned(101670364,32),
    to_unsigned(101876020,32),
    to_unsigned(102081675,32),
    to_unsigned(102287329,32),
    to_unsigned(102492982,32),
    to_unsigned(102698635,32),
    to_unsigned(102904286,32),
    to_unsigned(103109936,32),
    to_unsigned(103315586,32),
    to_unsigned(103521234,32),
    to_unsigned(103726882,32),
    to_unsigned(103932529,32),
    to_unsigned(104138174,32),
    to_unsigned(104343819,32),
    to_unsigned(104549463,32),
    to_unsigned(104755106,32),
    to_unsigned(104960747,32),
    to_unsigned(105166388,32),
    to_unsigned(105372028,32),
    to_unsigned(105577667,32),
    to_unsigned(105783305,32),
    to_unsigned(105988942,32),
    to_unsigned(106194578,32),
    to_unsigned(106400213,32),
    to_unsigned(106605847,32),
    to_unsigned(106811480,32),
    to_unsigned(107017112,32),
    to_unsigned(107222743,32),
    to_unsigned(107428374,32),
    to_unsigned(107634003,32),
    to_unsigned(107839631,32),
    to_unsigned(108045258,32),
    to_unsigned(108250884,32),
    to_unsigned(108456509,32),
    to_unsigned(108662134,32),
    to_unsigned(108867757,32),
    to_unsigned(109073379,32),
    to_unsigned(109279000,32),
    to_unsigned(109484620,32),
    to_unsigned(109690239,32),
    to_unsigned(109895858,32),
    to_unsigned(110101475,32),
    to_unsigned(110307091,32),
    to_unsigned(110512706,32),
    to_unsigned(110718320,32),
    to_unsigned(110923933,32),
    to_unsigned(111129545,32),
    to_unsigned(111335156,32),
    to_unsigned(111540766,32),
    to_unsigned(111746375,32),
    to_unsigned(111951983,32),
    to_unsigned(112157590,32),
    to_unsigned(112363196,32),
    to_unsigned(112568801,32),
    to_unsigned(112774405,32),
    to_unsigned(112980008,32),
    to_unsigned(113185609,32),
    to_unsigned(113391210,32),
    to_unsigned(113596810,32),
    to_unsigned(113802408,32),
    to_unsigned(114008006,32),
    to_unsigned(114213603,32),
    to_unsigned(114419198,32),
    to_unsigned(114624793,32),
    to_unsigned(114830386,32),
    to_unsigned(115035978,32),
    to_unsigned(115241570,32),
    to_unsigned(115447160,32),
    to_unsigned(115652749,32),
    to_unsigned(115858337,32),
    to_unsigned(116063924,32),
    to_unsigned(116269510,32),
    to_unsigned(116475095,32),
    to_unsigned(116680679,32),
    to_unsigned(116886261,32),
    to_unsigned(117091843,32),
    to_unsigned(117297424,32),
    to_unsigned(117503003,32),
    to_unsigned(117708582,32),
    to_unsigned(117914159,32),
    to_unsigned(118119735,32),
    to_unsigned(118325311,32),
    to_unsigned(118530885,32),
    to_unsigned(118736458,32),
    to_unsigned(118942030,32),
    to_unsigned(119147600,32),
    to_unsigned(119353170,32),
    to_unsigned(119558739,32),
    to_unsigned(119764306,32),
    to_unsigned(119969873,32),
    to_unsigned(120175438,32),
    to_unsigned(120381002,32),
    to_unsigned(120586565,32),
    to_unsigned(120792127,32),
    to_unsigned(120997688,32),
    to_unsigned(121203248,32),
    to_unsigned(121408807,32),
    to_unsigned(121614364,32),
    to_unsigned(121819921,32),
    to_unsigned(122025476,32),
    to_unsigned(122231030,32),
    to_unsigned(122436583,32),
    to_unsigned(122642135,32),
    to_unsigned(122847686,32),
    to_unsigned(123053236,32),
    to_unsigned(123258784,32),
    to_unsigned(123464332,32),
    to_unsigned(123669878,32),
    to_unsigned(123875423,32),
    to_unsigned(124080967,32),
    to_unsigned(124286510,32),
    to_unsigned(124492052,32),
    to_unsigned(124697593,32),
    to_unsigned(124903132,32),
    to_unsigned(125108670,32),
    to_unsigned(125314207,32),
    to_unsigned(125519743,32),
    to_unsigned(125725278,32),
    to_unsigned(125930812,32),
    to_unsigned(126136345,32),
    to_unsigned(126341876,32),
    to_unsigned(126547406,32),
    to_unsigned(126752935,32),
    to_unsigned(126958463,32),
    to_unsigned(127163990,32),
    to_unsigned(127369515,32),
    to_unsigned(127575040,32),
    to_unsigned(127780563,32),
    to_unsigned(127986085,32),
    to_unsigned(128191606,32),
    to_unsigned(128397125,32),
    to_unsigned(128602644,32),
    to_unsigned(128808161,32),
    to_unsigned(129013677,32),
    to_unsigned(129219192,32),
    to_unsigned(129424706,32),
    to_unsigned(129630219,32),
    to_unsigned(129835730,32),
    to_unsigned(130041240,32),
    to_unsigned(130246749,32),
    to_unsigned(130452257,32),
    to_unsigned(130657764,32),
    to_unsigned(130863269,32),
    to_unsigned(131068773,32),
    to_unsigned(131274276,32),
    to_unsigned(131479778,32),
    to_unsigned(131685278,32),
    to_unsigned(131890778,32),
    to_unsigned(132096276,32),
    to_unsigned(132301773,32),
    to_unsigned(132507269,32),
    to_unsigned(132712763,32),
    to_unsigned(132918256,32),
    to_unsigned(133123748,32),
    to_unsigned(133329239,32),
    to_unsigned(133534729,32),
    to_unsigned(133740217,32),
    to_unsigned(133945704,32),
    to_unsigned(134151190,32),
    to_unsigned(134356675,32),
    to_unsigned(134562158,32),
    to_unsigned(134767641,32),
    to_unsigned(134973122,32),
    to_unsigned(135178601,32),
    to_unsigned(135384080,32),
    to_unsigned(135589557,32),
    to_unsigned(135795033,32),
    to_unsigned(136000508,32),
    to_unsigned(136205981,32),
    to_unsigned(136411454,32),
    to_unsigned(136616924,32),
    to_unsigned(136822394,32),
    to_unsigned(137027863,32),
    to_unsigned(137233330,32),
    to_unsigned(137438796,32),
    to_unsigned(137644261,32),
    to_unsigned(137849724,32),
    to_unsigned(138055186,32),
    to_unsigned(138260647,32),
    to_unsigned(138466107,32),
    to_unsigned(138671565,32),
    to_unsigned(138877022,32),
    to_unsigned(139082478,32),
    to_unsigned(139287932,32),
    to_unsigned(139493386,32),
    to_unsigned(139698838,32),
    to_unsigned(139904288,32),
    to_unsigned(140109738,32),
    to_unsigned(140315186,32),
    to_unsigned(140520633,32),
    to_unsigned(140726078,32),
    to_unsigned(140931522,32),
    to_unsigned(141136965,32),
    to_unsigned(141342407,32),
    to_unsigned(141547847,32),
    to_unsigned(141753286,32),
    to_unsigned(141958724,32),
    to_unsigned(142164160,32),
    to_unsigned(142369596,32),
    to_unsigned(142575029,32),
    to_unsigned(142780462,32),
    to_unsigned(142985893,32),
    to_unsigned(143191323,32),
    to_unsigned(143396751,32),
    to_unsigned(143602179,32),
    to_unsigned(143807605,32),
    to_unsigned(144013029,32),
    to_unsigned(144218452,32),
    to_unsigned(144423874,32),
    to_unsigned(144629295,32),
    to_unsigned(144834714,32),
    to_unsigned(145040132,32),
    to_unsigned(145245549,32),
    to_unsigned(145450964,32),
    to_unsigned(145656378,32),
    to_unsigned(145861791,32),
    to_unsigned(146067202,32),
    to_unsigned(146272612,32),
    to_unsigned(146478021,32),
    to_unsigned(146683428,32),
    to_unsigned(146888834,32),
    to_unsigned(147094238,32),
    to_unsigned(147299641,32),
    to_unsigned(147505043,32),
    to_unsigned(147710444,32),
    to_unsigned(147915843,32),
    to_unsigned(148121241,32),
    to_unsigned(148326637,32),
    to_unsigned(148532032,32),
    to_unsigned(148737426,32),
    to_unsigned(148942818,32),
    to_unsigned(149148209,32),
    to_unsigned(149353599,32),
    to_unsigned(149558987,32),
    to_unsigned(149764374,32),
    to_unsigned(149969759,32),
    to_unsigned(150175143,32),
    to_unsigned(150380526,32),
    to_unsigned(150585907,32),
    to_unsigned(150791287,32),
    to_unsigned(150996665,32),
    to_unsigned(151202043,32),
    to_unsigned(151407418,32),
    to_unsigned(151612793,32),
    to_unsigned(151818166,32),
    to_unsigned(152023537,32),
    to_unsigned(152228907,32),
    to_unsigned(152434276,32),
    to_unsigned(152639644,32),
    to_unsigned(152845010,32),
    to_unsigned(153050374,32),
    to_unsigned(153255737,32),
    to_unsigned(153461099,32),
    to_unsigned(153666459,32),
    to_unsigned(153871818,32),
    to_unsigned(154077176,32),
    to_unsigned(154282532,32),
    to_unsigned(154487887,32),
    to_unsigned(154693240,32),
    to_unsigned(154898592,32),
    to_unsigned(155103942,32),
    to_unsigned(155309291,32),
    to_unsigned(155514639,32),
    to_unsigned(155719985,32),
    to_unsigned(155925329,32),
    to_unsigned(156130673,32),
    to_unsigned(156336015,32),
    to_unsigned(156541355,32),
    to_unsigned(156746694,32),
    to_unsigned(156952031,32),
    to_unsigned(157157368,32),
    to_unsigned(157362702,32),
    to_unsigned(157568035,32),
    to_unsigned(157773367,32),
    to_unsigned(157978697,32),
    to_unsigned(158184026,32),
    to_unsigned(158389354,32),
    to_unsigned(158594679,32),
    to_unsigned(158800004,32),
    to_unsigned(159005327,32),
    to_unsigned(159210648,32),
    to_unsigned(159415969,32),
    to_unsigned(159621287,32),
    to_unsigned(159826604,32),
    to_unsigned(160031920,32),
    to_unsigned(160237234,32),
    to_unsigned(160442547,32),
    to_unsigned(160647858,32),
    to_unsigned(160853168,32),
    to_unsigned(161058476,32),
    to_unsigned(161263783,32),
    to_unsigned(161469088,32),
    to_unsigned(161674392,32),
    to_unsigned(161879695,32),
    to_unsigned(162084995,32),
    to_unsigned(162290295,32),
    to_unsigned(162495593,32),
    to_unsigned(162700889,32),
    to_unsigned(162906184,32),
    to_unsigned(163111478,32),
    to_unsigned(163316769,32),
    to_unsigned(163522060,32),
    to_unsigned(163727349,32),
    to_unsigned(163932636,32),
    to_unsigned(164137922,32),
    to_unsigned(164343206,32),
    to_unsigned(164548489,32),
    to_unsigned(164753771,32),
    to_unsigned(164959051,32),
    to_unsigned(165164329,32),
    to_unsigned(165369606,32),
    to_unsigned(165574881,32),
    to_unsigned(165780155,32),
    to_unsigned(165985427,32),
    to_unsigned(166190698,32),
    to_unsigned(166395967,32),
    to_unsigned(166601235,32),
    to_unsigned(166806501,32),
    to_unsigned(167011765,32),
    to_unsigned(167217028,32),
    to_unsigned(167422290,32),
    to_unsigned(167627550,32),
    to_unsigned(167832808,32),
    to_unsigned(168038065,32),
    to_unsigned(168243321,32),
    to_unsigned(168448574,32),
    to_unsigned(168653827,32),
    to_unsigned(168859077,32),
    to_unsigned(169064327,32),
    to_unsigned(169269574,32),
    to_unsigned(169474820,32),
    to_unsigned(169680065,32),
    to_unsigned(169885308,32),
    to_unsigned(170090549,32),
    to_unsigned(170295789,32),
    to_unsigned(170501027,32),
    to_unsigned(170706264,32),
    to_unsigned(170911499,32),
    to_unsigned(171116732,32),
    to_unsigned(171321964,32),
    to_unsigned(171527195,32),
    to_unsigned(171732424,32),
    to_unsigned(171937651,32),
    to_unsigned(172142877,32),
    to_unsigned(172348101,32),
    to_unsigned(172553323,32),
    to_unsigned(172758544,32),
    to_unsigned(172963763,32),
    to_unsigned(173168981,32),
    to_unsigned(173374197,32),
    to_unsigned(173579412,32),
    to_unsigned(173784625,32),
    to_unsigned(173989836,32),
    to_unsigned(174195046,32),
    to_unsigned(174400254,32),
    to_unsigned(174605461,32),
    to_unsigned(174810665,32),
    to_unsigned(175015869,32),
    to_unsigned(175221071,32),
    to_unsigned(175426271,32),
    to_unsigned(175631469,32),
    to_unsigned(175836666,32),
    to_unsigned(176041861,32),
    to_unsigned(176247055,32),
    to_unsigned(176452247,32),
    to_unsigned(176657437,32),
    to_unsigned(176862626,32),
    to_unsigned(177067813,32),
    to_unsigned(177272999,32),
    to_unsigned(177478183,32),
    to_unsigned(177683365,32),
    to_unsigned(177888546,32),
    to_unsigned(178093725,32),
    to_unsigned(178298902,32),
    to_unsigned(178504078,32),
    to_unsigned(178709252,32),
    to_unsigned(178914424,32),
    to_unsigned(179119595,32),
    to_unsigned(179324764,32),
    to_unsigned(179529932,32),
    to_unsigned(179735098,32),
    to_unsigned(179940262,32),
    to_unsigned(180145424,32),
    to_unsigned(180350585,32),
    to_unsigned(180555745,32),
    to_unsigned(180760902,32),
    to_unsigned(180966058,32),
    to_unsigned(181171212,32),
    to_unsigned(181376365,32),
    to_unsigned(181581516,32),
    to_unsigned(181786665,32),
    to_unsigned(181991813,32),
    to_unsigned(182196959,32),
    to_unsigned(182402103,32),
    to_unsigned(182607245,32),
    to_unsigned(182812386,32),
    to_unsigned(183017525,32),
    to_unsigned(183222663,32),
    to_unsigned(183427799,32),
    to_unsigned(183632933,32),
    to_unsigned(183838065,32),
    to_unsigned(184043196,32),
    to_unsigned(184248325,32),
    to_unsigned(184453453,32),
    to_unsigned(184658578,32),
    to_unsigned(184863702,32),
    to_unsigned(185068825,32),
    to_unsigned(185273945,32),
    to_unsigned(185479064,32),
    to_unsigned(185684181,32),
    to_unsigned(185889297,32),
    to_unsigned(186094410,32),
    to_unsigned(186299523,32),
    to_unsigned(186504633,32),
    to_unsigned(186709741,32),
    to_unsigned(186914848,32),
    to_unsigned(187119954,32),
    to_unsigned(187325057,32),
    to_unsigned(187530159,32),
    to_unsigned(187735259,32),
    to_unsigned(187940357,32),
    to_unsigned(188145454,32),
    to_unsigned(188350549,32),
    to_unsigned(188555642,32),
    to_unsigned(188760733,32),
    to_unsigned(188965823,32),
    to_unsigned(189170911,32),
    to_unsigned(189375997,32),
    to_unsigned(189581081,32),
    to_unsigned(189786164,32),
    to_unsigned(189991245,32),
    to_unsigned(190196324,32),
    to_unsigned(190401402,32),
    to_unsigned(190606477,32),
    to_unsigned(190811551,32),
    to_unsigned(191016623,32),
    to_unsigned(191221694,32),
    to_unsigned(191426762,32),
    to_unsigned(191631829,32),
    to_unsigned(191836895,32),
    to_unsigned(192041958,32),
    to_unsigned(192247020,32),
    to_unsigned(192452079,32),
    to_unsigned(192657138,32),
    to_unsigned(192862194,32),
    to_unsigned(193067248,32),
    to_unsigned(193272301,32),
    to_unsigned(193477352,32),
    to_unsigned(193682401,32),
    to_unsigned(193887449,32),
    to_unsigned(194092494,32),
    to_unsigned(194297538,32),
    to_unsigned(194502580,32),
    to_unsigned(194707621,32),
    to_unsigned(194912659,32),
    to_unsigned(195117696,32),
    to_unsigned(195322731,32),
    to_unsigned(195527764,32),
    to_unsigned(195732795,32),
    to_unsigned(195937825,32),
    to_unsigned(196142853,32),
    to_unsigned(196347879,32),
    to_unsigned(196552903,32),
    to_unsigned(196757925,32),
    to_unsigned(196962946,32),
    to_unsigned(197167964,32),
    to_unsigned(197372981,32),
    to_unsigned(197577996,32),
    to_unsigned(197783009,32),
    to_unsigned(197988021,32),
    to_unsigned(198193030,32),
    to_unsigned(198398038,32),
    to_unsigned(198603044,32),
    to_unsigned(198808048,32),
    to_unsigned(199013051,32),
    to_unsigned(199218051,32),
    to_unsigned(199423050,32),
    to_unsigned(199628047,32),
    to_unsigned(199833042,32),
    to_unsigned(200038035,32),
    to_unsigned(200243026,32),
    to_unsigned(200448016,32),
    to_unsigned(200653003,32),
    to_unsigned(200857989,32),
    to_unsigned(201062973,32),
    to_unsigned(201267955,32),
    to_unsigned(201472935,32),
    to_unsigned(201677914,32),
    to_unsigned(201882890,32),
    to_unsigned(202087865,32),
    to_unsigned(202292838,32),
    to_unsigned(202497809,32),
    to_unsigned(202702778,32),
    to_unsigned(202907745,32),
    to_unsigned(203112710,32),
    to_unsigned(203317674,32),
    to_unsigned(203522636,32),
    to_unsigned(203727595,32),
    to_unsigned(203932553,32),
    to_unsigned(204137509,32),
    to_unsigned(204342463,32),
    to_unsigned(204547416,32),
    to_unsigned(204752366,32),
    to_unsigned(204957315,32),
    to_unsigned(205162261,32),
    to_unsigned(205367206,32),
    to_unsigned(205572149,32),
    to_unsigned(205777090,32),
    to_unsigned(205982029,32),
    to_unsigned(206186966,32),
    to_unsigned(206391901,32),
    to_unsigned(206596835,32),
    to_unsigned(206801766,32),
    to_unsigned(207006696,32),
    to_unsigned(207211623,32),
    to_unsigned(207416549,32),
    to_unsigned(207621473,32),
    to_unsigned(207826395,32),
    to_unsigned(208031315,32),
    to_unsigned(208236233,32),
    to_unsigned(208441149,32),
    to_unsigned(208646064,32),
    to_unsigned(208850976,32),
    to_unsigned(209055887,32),
    to_unsigned(209260795,32),
    to_unsigned(209465702,32),
    to_unsigned(209670606,32),
    to_unsigned(209875509,32),
    to_unsigned(210080410,32),
    to_unsigned(210285309,32),
    to_unsigned(210490206,32),
    to_unsigned(210695101,32),
    to_unsigned(210899994,32),
    to_unsigned(211104885,32),
    to_unsigned(211309775,32),
    to_unsigned(211514662,32),
    to_unsigned(211719547,32),
    to_unsigned(211924431,32),
    to_unsigned(212129312,32),
    to_unsigned(212334192,32),
    to_unsigned(212539069,32),
    to_unsigned(212743945,32),
    to_unsigned(212948818,32),
    to_unsigned(213153690,32),
    to_unsigned(213358560,32),
    to_unsigned(213563427,32),
    to_unsigned(213768293,32),
    to_unsigned(213973157,32),
    to_unsigned(214178019,32),
    to_unsigned(214382879,32),
    to_unsigned(214587737,32),
    to_unsigned(214792593,32),
    to_unsigned(214997447,32),
    to_unsigned(215202299,32),
    to_unsigned(215407149,32),
    to_unsigned(215611997,32),
    to_unsigned(215816843,32),
    to_unsigned(216021687,32),
    to_unsigned(216226529,32),
    to_unsigned(216431369,32),
    to_unsigned(216636207,32),
    to_unsigned(216841043,32),
    to_unsigned(217045877,32),
    to_unsigned(217250710,32),
    to_unsigned(217455540,32),
    to_unsigned(217660368,32),
    to_unsigned(217865194,32),
    to_unsigned(218070018,32),
    to_unsigned(218274840,32),
    to_unsigned(218479660,32),
    to_unsigned(218684479,32),
    to_unsigned(218889295,32),
    to_unsigned(219094109,32),
    to_unsigned(219298921,32),
    to_unsigned(219503731,32),
    to_unsigned(219708539,32),
    to_unsigned(219913345,32),
    to_unsigned(220118149,32),
    to_unsigned(220322951,32),
    to_unsigned(220527751,32),
    to_unsigned(220732549,32),
    to_unsigned(220937345,32),
    to_unsigned(221142139,32),
    to_unsigned(221346930,32),
    to_unsigned(221551720,32),
    to_unsigned(221756508,32),
    to_unsigned(221961294,32),
    to_unsigned(222166077,32),
    to_unsigned(222370859,32),
    to_unsigned(222575639,32),
    to_unsigned(222780416,32),
    to_unsigned(222985192,32),
    to_unsigned(223189965,32),
    to_unsigned(223394737,32),
    to_unsigned(223599506,32),
    to_unsigned(223804273,32),
    to_unsigned(224009039,32),
    to_unsigned(224213802,32),
    to_unsigned(224418563,32),
    to_unsigned(224623322,32),
    to_unsigned(224828079,32),
    to_unsigned(225032834,32),
    to_unsigned(225237587,32),
    to_unsigned(225442338,32),
    to_unsigned(225647086,32),
    to_unsigned(225851833,32),
    to_unsigned(226056577,32),
    to_unsigned(226261320,32),
    to_unsigned(226466060,32),
    to_unsigned(226670799,32),
    to_unsigned(226875535,32),
    to_unsigned(227080269,32),
    to_unsigned(227285001,32),
    to_unsigned(227489731,32),
    to_unsigned(227694459,32),
    to_unsigned(227899185,32),
    to_unsigned(228103909,32),
    to_unsigned(228308630,32),
    to_unsigned(228513350,32),
    to_unsigned(228718067,32),
    to_unsigned(228922782,32),
    to_unsigned(229127496,32),
    to_unsigned(229332207,32),
    to_unsigned(229536916,32),
    to_unsigned(229741623,32),
    to_unsigned(229946327,32),
    to_unsigned(230151030,32),
    to_unsigned(230355731,32),
    to_unsigned(230560429,32),
    to_unsigned(230765125,32),
    to_unsigned(230969819,32),
    to_unsigned(231174512,32),
    to_unsigned(231379201,32),
    to_unsigned(231583889,32),
    to_unsigned(231788575,32),
    to_unsigned(231993258,32),
    to_unsigned(232197940,32),
    to_unsigned(232402619,32),
    to_unsigned(232607296,32),
    to_unsigned(232811971,32),
    to_unsigned(233016644,32),
    to_unsigned(233221315,32),
    to_unsigned(233425983,32),
    to_unsigned(233630650,32),
    to_unsigned(233835314,32),
    to_unsigned(234039976,32),
    to_unsigned(234244636,32),
    to_unsigned(234449294,32),
    to_unsigned(234653950,32),
    to_unsigned(234858603,32),
    to_unsigned(235063255,32),
    to_unsigned(235267904,32),
    to_unsigned(235472551,32),
    to_unsigned(235677196,32),
    to_unsigned(235881839,32),
    to_unsigned(236086479,32),
    to_unsigned(236291117,32),
    to_unsigned(236495754,32),
    to_unsigned(236700388,32),
    to_unsigned(236905020,32),
    to_unsigned(237109649,32),
    to_unsigned(237314277,32),
    to_unsigned(237518902,32),
    to_unsigned(237723525,32),
    to_unsigned(237928146,32),
    to_unsigned(238132765,32),
    to_unsigned(238337381,32),
    to_unsigned(238541996,32),
    to_unsigned(238746608,32),
    to_unsigned(238951218,32),
    to_unsigned(239155826,32),
    to_unsigned(239360431,32),
    to_unsigned(239565035,32),
    to_unsigned(239769636,32),
    to_unsigned(239974235,32),
    to_unsigned(240178832,32),
    to_unsigned(240383426,32),
    to_unsigned(240588019,32),
    to_unsigned(240792609,32),
    to_unsigned(240997197,32),
    to_unsigned(241201782,32),
    to_unsigned(241406366,32),
    to_unsigned(241610947,32),
    to_unsigned(241815526,32),
    to_unsigned(242020103,32),
    to_unsigned(242224678,32),
    to_unsigned(242429250,32),
    to_unsigned(242633820,32),
    to_unsigned(242838388,32),
    to_unsigned(243042954,32),
    to_unsigned(243247517,32),
    to_unsigned(243452079,32),
    to_unsigned(243656638,32),
    to_unsigned(243861194,32),
    to_unsigned(244065749,32),
    to_unsigned(244270301,32),
    to_unsigned(244474851,32),
    to_unsigned(244679399,32),
    to_unsigned(244883945,32),
    to_unsigned(245088488,32),
    to_unsigned(245293029,32),
    to_unsigned(245497568,32),
    to_unsigned(245702104,32),
    to_unsigned(245906638,32),
    to_unsigned(246111170,32),
    to_unsigned(246315700,32),
    to_unsigned(246520228,32),
    to_unsigned(246724753,32),
    to_unsigned(246929276,32),
    to_unsigned(247133796,32),
    to_unsigned(247338315,32),
    to_unsigned(247542831,32),
    to_unsigned(247747345,32),
    to_unsigned(247951856,32),
    to_unsigned(248156366,32),
    to_unsigned(248360873,32),
    to_unsigned(248565377,32),
    to_unsigned(248769880,32),
    to_unsigned(248974380,32),
    to_unsigned(249178878,32),
    to_unsigned(249383373,32),
    to_unsigned(249587867,32),
    to_unsigned(249792358,32),
    to_unsigned(249996846,32),
    to_unsigned(250201333,32),
    to_unsigned(250405817,32),
    to_unsigned(250610299,32),
    to_unsigned(250814778,32),
    to_unsigned(251019255,32),
    to_unsigned(251223730,32),
    to_unsigned(251428203,32),
    to_unsigned(251632673,32),
    to_unsigned(251837141,32),
    to_unsigned(252041607,32),
    to_unsigned(252246070,32),
    to_unsigned(252450531,32),
    to_unsigned(252654990,32),
    to_unsigned(252859446,32),
    to_unsigned(253063900,32),
    to_unsigned(253268352,32),
    to_unsigned(253472801,32),
    to_unsigned(253677248,32),
    to_unsigned(253881693,32),
    to_unsigned(254086135,32),
    to_unsigned(254290575,32),
    to_unsigned(254495013,32),
    to_unsigned(254699448,32),
    to_unsigned(254903881,32),
    to_unsigned(255108312,32),
    to_unsigned(255312740,32),
    to_unsigned(255517166,32),
    to_unsigned(255721590,32),
    to_unsigned(255926011,32),
    to_unsigned(256130430,32),
    to_unsigned(256334847,32),
    to_unsigned(256539261,32),
    to_unsigned(256743673,32),
    to_unsigned(256948082,32),
    to_unsigned(257152490,32),
    to_unsigned(257356894,32),
    to_unsigned(257561297,32),
    to_unsigned(257765697,32),
    to_unsigned(257970095,32),
    to_unsigned(258174490,32),
    to_unsigned(258378883,32),
    to_unsigned(258583273,32),
    to_unsigned(258787662,32),
    to_unsigned(258992047,32),
    to_unsigned(259196431,32),
    to_unsigned(259400812,32),
    to_unsigned(259605190,32),
    to_unsigned(259809567,32),
    to_unsigned(260013941,32),
    to_unsigned(260218312,32),
    to_unsigned(260422681,32),
    to_unsigned(260627048,32),
    to_unsigned(260831412,32),
    to_unsigned(261035774,32),
    to_unsigned(261240134,32),
    to_unsigned(261444491,32),
    to_unsigned(261648846,32),
    to_unsigned(261853198,32),
    to_unsigned(262057548,32),
    to_unsigned(262261895,32),
    to_unsigned(262466240,32),
    to_unsigned(262670583,32),
    to_unsigned(262874923,32),
    to_unsigned(263079261,32),
    to_unsigned(263283596,32),
    to_unsigned(263487929,32),
    to_unsigned(263692260,32),
    to_unsigned(263896588,32),
    to_unsigned(264100914,32),
    to_unsigned(264305237,32),
    to_unsigned(264509558,32),
    to_unsigned(264713877,32),
    to_unsigned(264918193,32),
    to_unsigned(265122506,32),
    to_unsigned(265326817,32),
    to_unsigned(265531126,32),
    to_unsigned(265735432,32),
    to_unsigned(265939736,32),
    to_unsigned(266144037,32),
    to_unsigned(266348336,32),
    to_unsigned(266552633,32),
    to_unsigned(266756927,32),
    to_unsigned(266961218,32),
    to_unsigned(267165508,32),
    to_unsigned(267369794,32),
    to_unsigned(267574078,32),
    to_unsigned(267778360,32),
    to_unsigned(267982639,32),
    to_unsigned(268186916,32),
    to_unsigned(268391191,32),
    to_unsigned(268595462,32),
    to_unsigned(268799732,32),
    to_unsigned(269003999,32),
    to_unsigned(269208263,32),
    to_unsigned(269412525,32),
    to_unsigned(269616785,32),
    to_unsigned(269821042,32),
    to_unsigned(270025296,32),
    to_unsigned(270229549,32),
    to_unsigned(270433798,32),
    to_unsigned(270638045,32),
    to_unsigned(270842290,32),
    to_unsigned(271046532,32),
    to_unsigned(271250772,32),
    to_unsigned(271455009,32),
    to_unsigned(271659243,32),
    to_unsigned(271863476,32),
    to_unsigned(272067705,32),
    to_unsigned(272271932,32),
    to_unsigned(272476157,32),
    to_unsigned(272680379,32),
    to_unsigned(272884599,32),
    to_unsigned(273088816,32),
    to_unsigned(273293031,32),
    to_unsigned(273497243,32),
    to_unsigned(273701452,32),
    to_unsigned(273905660,32),
    to_unsigned(274109864,32),
    to_unsigned(274314066,32),
    to_unsigned(274518266,32),
    to_unsigned(274722463,32),
    to_unsigned(274926657,32),
    to_unsigned(275130849,32),
    to_unsigned(275335039,32),
    to_unsigned(275539225,32),
    to_unsigned(275743410,32),
    to_unsigned(275947592,32),
    to_unsigned(276151771,32),
    to_unsigned(276355948,32),
    to_unsigned(276560122,32),
    to_unsigned(276764294,32),
    to_unsigned(276968463,32),
    to_unsigned(277172629,32),
    to_unsigned(277376793,32),
    to_unsigned(277580955,32),
    to_unsigned(277785114,32),
    to_unsigned(277989270,32),
    to_unsigned(278193424,32),
    to_unsigned(278397575,32),
    to_unsigned(278601724,32),
    to_unsigned(278805870,32),
    to_unsigned(279010014,32),
    to_unsigned(279214155,32),
    to_unsigned(279418293,32),
    to_unsigned(279622429,32),
    to_unsigned(279826562,32),
    to_unsigned(280030693,32),
    to_unsigned(280234821,32),
    to_unsigned(280438947,32),
    to_unsigned(280643070,32),
    to_unsigned(280847190,32),
    to_unsigned(281051308,32),
    to_unsigned(281255423,32),
    to_unsigned(281459536,32),
    to_unsigned(281663646,32),
    to_unsigned(281867754,32),
    to_unsigned(282071859,32),
    to_unsigned(282275961,32),
    to_unsigned(282480061,32),
    to_unsigned(282684158,32),
    to_unsigned(282888252,32),
    to_unsigned(283092344,32),
    to_unsigned(283296433,32),
    to_unsigned(283500520,32),
    to_unsigned(283704604,32),
    to_unsigned(283908686,32),
    to_unsigned(284112765,32),
    to_unsigned(284316841,32),
    to_unsigned(284520915,32),
    to_unsigned(284724986,32),
    to_unsigned(284929054,32),
    to_unsigned(285133120,32),
    to_unsigned(285337183,32),
    to_unsigned(285541244,32),
    to_unsigned(285745302,32),
    to_unsigned(285949357,32),
    to_unsigned(286153410,32),
    to_unsigned(286357460,32),
    to_unsigned(286561507,32),
    to_unsigned(286765552,32),
    to_unsigned(286969594,32),
    to_unsigned(287173634,32),
    to_unsigned(287377671,32),
    to_unsigned(287581705,32),
    to_unsigned(287785737,32),
    to_unsigned(287989766,32),
    to_unsigned(288193792,32),
    to_unsigned(288397816,32),
    to_unsigned(288601837,32),
    to_unsigned(288805855,32),
    to_unsigned(289009871,32),
    to_unsigned(289213884,32),
    to_unsigned(289417894,32),
    to_unsigned(289621902,32),
    to_unsigned(289825907,32),
    to_unsigned(290029909,32),
    to_unsigned(290233909,32),
    to_unsigned(290437906,32),
    to_unsigned(290641901,32),
    to_unsigned(290845892,32),
    to_unsigned(291049881,32),
    to_unsigned(291253868,32),
    to_unsigned(291457852,32),
    to_unsigned(291661833,32),
    to_unsigned(291865811,32),
    to_unsigned(292069787,32),
    to_unsigned(292273760,32),
    to_unsigned(292477730,32),
    to_unsigned(292681697,32),
    to_unsigned(292885662,32),
    to_unsigned(293089625,32),
    to_unsigned(293293584,32),
    to_unsigned(293497541,32),
    to_unsigned(293701495,32),
    to_unsigned(293905447,32),
    to_unsigned(294109395,32),
    to_unsigned(294313341,32),
    to_unsigned(294517285,32),
    to_unsigned(294721225,32),
    to_unsigned(294925163,32),
    to_unsigned(295129098,32),
    to_unsigned(295333031,32),
    to_unsigned(295536961,32),
    to_unsigned(295740888,32),
    to_unsigned(295944812,32),
    to_unsigned(296148734,32),
    to_unsigned(296352653,32),
    to_unsigned(296556569,32),
    to_unsigned(296760482,32),
    to_unsigned(296964393,32),
    to_unsigned(297168301,32),
    to_unsigned(297372206,32),
    to_unsigned(297576109,32),
    to_unsigned(297780008,32),
    to_unsigned(297983905,32),
    to_unsigned(298187800,32),
    to_unsigned(298391691,32),
    to_unsigned(298595580,32),
    to_unsigned(298799466,32),
    to_unsigned(299003350,32),
    to_unsigned(299207230,32),
    to_unsigned(299411108,32),
    to_unsigned(299614983,32),
    to_unsigned(299818855,32),
    to_unsigned(300022725,32),
    to_unsigned(300226592,32),
    to_unsigned(300430456,32),
    to_unsigned(300634317,32),
    to_unsigned(300838176,32),
    to_unsigned(301042031,32),
    to_unsigned(301245884,32),
    to_unsigned(301449735,32),
    to_unsigned(301653582,32),
    to_unsigned(301857427,32),
    to_unsigned(302061269,32),
    to_unsigned(302265108,32),
    to_unsigned(302468944,32),
    to_unsigned(302672778,32),
    to_unsigned(302876609,32),
    to_unsigned(303080437,32),
    to_unsigned(303284262,32),
    to_unsigned(303488084,32),
    to_unsigned(303691904,32),
    to_unsigned(303895721,32),
    to_unsigned(304099535,32),
    to_unsigned(304303346,32),
    to_unsigned(304507155,32),
    to_unsigned(304710960,32),
    to_unsigned(304914763,32),
    to_unsigned(305118563,32),
    to_unsigned(305322361,32),
    to_unsigned(305526155,32),
    to_unsigned(305729947,32),
    to_unsigned(305933735,32),
    to_unsigned(306137522,32),
    to_unsigned(306341305,32),
    to_unsigned(306545085,32),
    to_unsigned(306748863,32),
    to_unsigned(306952637,32),
    to_unsigned(307156409,32),
    to_unsigned(307360179,32),
    to_unsigned(307563945,32),
    to_unsigned(307767708,32),
    to_unsigned(307971469,32),
    to_unsigned(308175227,32),
    to_unsigned(308378982,32),
    to_unsigned(308582734,32),
    to_unsigned(308786483,32),
    to_unsigned(308990230,32),
    to_unsigned(309193973,32),
    to_unsigned(309397714,32),
    to_unsigned(309601452,32),
    to_unsigned(309805187,32),
    to_unsigned(310008919,32),
    to_unsigned(310212649,32),
    to_unsigned(310416375,32),
    to_unsigned(310620099,32),
    to_unsigned(310823820,32),
    to_unsigned(311027538,32),
    to_unsigned(311231253,32),
    to_unsigned(311434965,32),
    to_unsigned(311638674,32),
    to_unsigned(311842381,32),
    to_unsigned(312046085,32),
    to_unsigned(312249785,32),
    to_unsigned(312453483,32),
    to_unsigned(312657178,32),
    to_unsigned(312860871,32),
    to_unsigned(313064560,32),
    to_unsigned(313268246,32),
    to_unsigned(313471930,32),
    to_unsigned(313675611,32),
    to_unsigned(313879288,32),
    to_unsigned(314082963,32),
    to_unsigned(314286635,32),
    to_unsigned(314490304,32),
    to_unsigned(314693971,32),
    to_unsigned(314897634,32),
    to_unsigned(315101294,32),
    to_unsigned(315304952,32),
    to_unsigned(315508607,32),
    to_unsigned(315712258,32),
    to_unsigned(315915907,32),
    to_unsigned(316119553,32),
    to_unsigned(316323196,32),
    to_unsigned(316526836,32),
    to_unsigned(316730474,32),
    to_unsigned(316934108,32),
    to_unsigned(317137739,32),
    to_unsigned(317341368,32),
    to_unsigned(317544993,32),
    to_unsigned(317748616,32),
    to_unsigned(317952236,32),
    to_unsigned(318155852,32),
    to_unsigned(318359466,32),
    to_unsigned(318563077,32),
    to_unsigned(318766685,32),
    to_unsigned(318970290,32),
    to_unsigned(319173893,32),
    to_unsigned(319377492,32),
    to_unsigned(319581088,32),
    to_unsigned(319784681,32),
    to_unsigned(319988272,32),
    to_unsigned(320191859,32),
    to_unsigned(320395444,32),
    to_unsigned(320599025,32),
    to_unsigned(320802604,32),
    to_unsigned(321006180,32),
    to_unsigned(321209753,32),
    to_unsigned(321413322,32),
    to_unsigned(321616889,32),
    to_unsigned(321820453,32),
    to_unsigned(322024014,32),
    to_unsigned(322227572,32),
    to_unsigned(322431127,32),
    to_unsigned(322634679,32),
    to_unsigned(322838228,32),
    to_unsigned(323041774,32),
    to_unsigned(323245317,32),
    to_unsigned(323448857,32),
    to_unsigned(323652395,32),
    to_unsigned(323855929,32),
    to_unsigned(324059460,32),
    to_unsigned(324262988,32),
    to_unsigned(324466514,32),
    to_unsigned(324670036,32),
    to_unsigned(324873555,32),
    to_unsigned(325077071,32),
    to_unsigned(325280585,32),
    to_unsigned(325484095,32),
    to_unsigned(325687602,32),
    to_unsigned(325891107,32),
    to_unsigned(326094608,32),
    to_unsigned(326298107,32),
    to_unsigned(326501602,32),
    to_unsigned(326705094,32),
    to_unsigned(326908584,32),
    to_unsigned(327112070,32),
    to_unsigned(327315553,32),
    to_unsigned(327519034,32),
    to_unsigned(327722511,32),
    to_unsigned(327925985,32),
    to_unsigned(328129457,32),
    to_unsigned(328332925,32),
    to_unsigned(328536390,32),
    to_unsigned(328739852,32),
    to_unsigned(328943312,32),
    to_unsigned(329146768,32),
    to_unsigned(329350221,32),
    to_unsigned(329553671,32),
    to_unsigned(329757118,32),
    to_unsigned(329960562,32),
    to_unsigned(330164004,32),
    to_unsigned(330367442,32),
    to_unsigned(330570877,32),
    to_unsigned(330774308,32),
    to_unsigned(330977737,32),
    to_unsigned(331181163,32),
    to_unsigned(331384586,32),
    to_unsigned(331588006,32),
    to_unsigned(331791423,32),
    to_unsigned(331994836,32),
    to_unsigned(332198247,32),
    to_unsigned(332401654,32),
    to_unsigned(332605059,32),
    to_unsigned(332808460,32),
    to_unsigned(333011859,32),
    to_unsigned(333215254,32),
    to_unsigned(333418646,32),
    to_unsigned(333622036,32),
    to_unsigned(333825422,32),
    to_unsigned(334028805,32),
    to_unsigned(334232185,32),
    to_unsigned(334435562,32),
    to_unsigned(334638936,32),
    to_unsigned(334842306,32),
    to_unsigned(335045674,32),
    to_unsigned(335249039,32),
    to_unsigned(335452400,32),
    to_unsigned(335655759,32),
    to_unsigned(335859114,32),
    to_unsigned(336062467,32),
    to_unsigned(336265816,32),
    to_unsigned(336469162,32),
    to_unsigned(336672505,32),
    to_unsigned(336875845,32),
    to_unsigned(337079182,32),
    to_unsigned(337282515,32),
    to_unsigned(337485846,32),
    to_unsigned(337689173,32),
    to_unsigned(337892498,32),
    to_unsigned(338095819,32),
    to_unsigned(338299137,32),
    to_unsigned(338502453,32),
    to_unsigned(338705765,32),
    to_unsigned(338909073,32),
    to_unsigned(339112379,32),
    to_unsigned(339315682,32),
    to_unsigned(339518981,32),
    to_unsigned(339722278,32),
    to_unsigned(339925571,32),
    to_unsigned(340128861,32),
    to_unsigned(340332148,32),
    to_unsigned(340535432,32),
    to_unsigned(340738713,32),
    to_unsigned(340941990,32),
    to_unsigned(341145265,32),
    to_unsigned(341348536,32),
    to_unsigned(341551805,32),
    to_unsigned(341755070,32),
    to_unsigned(341958332,32),
    to_unsigned(342161590,32),
    to_unsigned(342364846,32),
    to_unsigned(342568099,32),
    to_unsigned(342771348,32),
    to_unsigned(342974594,32),
    to_unsigned(343177837,32),
    to_unsigned(343381077,32),
    to_unsigned(343584314,32),
    to_unsigned(343787548,32),
    to_unsigned(343990778,32),
    to_unsigned(344194005,32),
    to_unsigned(344397229,32),
    to_unsigned(344600450,32),
    to_unsigned(344803668,32),
    to_unsigned(345006883,32),
    to_unsigned(345210094,32),
    to_unsigned(345413302,32),
    to_unsigned(345616507,32),
    to_unsigned(345819709,32),
    to_unsigned(346022908,32),
    to_unsigned(346226104,32),
    to_unsigned(346429296,32),
    to_unsigned(346632485,32),
    to_unsigned(346835671,32),
    to_unsigned(347038854,32),
    to_unsigned(347242034,32),
    to_unsigned(347445210,32),
    to_unsigned(347648383,32),
    to_unsigned(347851553,32),
    to_unsigned(348054720,32),
    to_unsigned(348257884,32),
    to_unsigned(348461044,32),
    to_unsigned(348664202,32),
    to_unsigned(348867356,32),
    to_unsigned(349070506,32),
    to_unsigned(349273654,32),
    to_unsigned(349476798,32),
    to_unsigned(349679940,32),
    to_unsigned(349883078,32),
    to_unsigned(350086212,32),
    to_unsigned(350289344,32),
    to_unsigned(350492472,32),
    to_unsigned(350695597,32),
    to_unsigned(350898719,32),
    to_unsigned(351101838,32),
    to_unsigned(351304953,32),
    to_unsigned(351508066,32),
    to_unsigned(351711174,32),
    to_unsigned(351914280,32),
    to_unsigned(352117383,32),
    to_unsigned(352320482,32),
    to_unsigned(352523578,32),
    to_unsigned(352726671,32),
    to_unsigned(352929760,32),
    to_unsigned(353132847,32),
    to_unsigned(353335930,32),
    to_unsigned(353539010,32),
    to_unsigned(353742086,32),
    to_unsigned(353945159,32),
    to_unsigned(354148229,32),
    to_unsigned(354351296,32),
    to_unsigned(354554360,32),
    to_unsigned(354757420,32),
    to_unsigned(354960477,32),
    to_unsigned(355163531,32),
    to_unsigned(355366581,32),
    to_unsigned(355569629,32),
    to_unsigned(355772673,32),
    to_unsigned(355975713,32),
    to_unsigned(356178751,32),
    to_unsigned(356381785,32),
    to_unsigned(356584816,32),
    to_unsigned(356787843,32),
    to_unsigned(356990868,32),
    to_unsigned(357193889,32),
    to_unsigned(357396906,32),
    to_unsigned(357599921,32),
    to_unsigned(357802932,32),
    to_unsigned(358005940,32),
    to_unsigned(358208944,32),
    to_unsigned(358411946,32),
    to_unsigned(358614944,32),
    to_unsigned(358817938,32),
    to_unsigned(359020930,32),
    to_unsigned(359223918,32),
    to_unsigned(359426903,32),
    to_unsigned(359629884,32),
    to_unsigned(359832862,32),
    to_unsigned(360035837,32),
    to_unsigned(360238809,32),
    to_unsigned(360441777,32),
    to_unsigned(360644742,32),
    to_unsigned(360847704,32),
    to_unsigned(361050662,32),
    to_unsigned(361253617,32),
    to_unsigned(361456569,32),
    to_unsigned(361659517,32),
    to_unsigned(361862462,32),
    to_unsigned(362065404,32),
    to_unsigned(362268342,32),
    to_unsigned(362471277,32),
    to_unsigned(362674209,32),
    to_unsigned(362877138,32),
    to_unsigned(363080063,32),
    to_unsigned(363282984,32),
    to_unsigned(363485903,32),
    to_unsigned(363688818,32),
    to_unsigned(363891729,32),
    to_unsigned(364094638,32),
    to_unsigned(364297543,32),
    to_unsigned(364500444,32),
    to_unsigned(364703343,32),
    to_unsigned(364906238,32),
    to_unsigned(365109129,32),
    to_unsigned(365312018,32),
    to_unsigned(365514902,32),
    to_unsigned(365717784,32),
    to_unsigned(365920662,32),
    to_unsigned(366123537,32),
    to_unsigned(366326408,32),
    to_unsigned(366529276,32),
    to_unsigned(366732141,32),
    to_unsigned(366935002,32),
    to_unsigned(367137860,32),
    to_unsigned(367340715,32),
    to_unsigned(367543566,32),
    to_unsigned(367746414,32),
    to_unsigned(367949258,32),
    to_unsigned(368152099,32),
    to_unsigned(368354937,32),
    to_unsigned(368557771,32),
    to_unsigned(368760602,32),
    to_unsigned(368963430,32),
    to_unsigned(369166254,32),
    to_unsigned(369369075,32),
    to_unsigned(369571892,32),
    to_unsigned(369774706,32),
    to_unsigned(369977517,32),
    to_unsigned(370180324,32),
    to_unsigned(370383127,32),
    to_unsigned(370585928,32),
    to_unsigned(370788725,32),
    to_unsigned(370991518,32),
    to_unsigned(371194308,32),
    to_unsigned(371397095,32),
    to_unsigned(371599878,32),
    to_unsigned(371802658,32),
    to_unsigned(372005435,32),
    to_unsigned(372208208,32),
    to_unsigned(372410977,32),
    to_unsigned(372613743,32),
    to_unsigned(372816506,32),
    to_unsigned(373019266,32),
    to_unsigned(373222021,32),
    to_unsigned(373424774,32),
    to_unsigned(373627523,32),
    to_unsigned(373830269,32),
    to_unsigned(374033011,32),
    to_unsigned(374235749,32),
    to_unsigned(374438485,32),
    to_unsigned(374641217,32),
    to_unsigned(374843945,32),
    to_unsigned(375046670,32),
    to_unsigned(375249391,32),
    to_unsigned(375452110,32),
    to_unsigned(375654824,32),
    to_unsigned(375857535,32),
    to_unsigned(376060243,32),
    to_unsigned(376262947,32),
    to_unsigned(376465648,32),
    to_unsigned(376668345,32),
    to_unsigned(376871039,32),
    to_unsigned(377073730,32),
    to_unsigned(377276417,32),
    to_unsigned(377479100,32),
    to_unsigned(377681780,32),
    to_unsigned(377884457,32),
    to_unsigned(378087130,32),
    to_unsigned(378289799,32),
    to_unsigned(378492465,32),
    to_unsigned(378695128,32),
    to_unsigned(378897787,32),
    to_unsigned(379100443,32),
    to_unsigned(379303095,32),
    to_unsigned(379505744,32),
    to_unsigned(379708389,32),
    to_unsigned(379911031,32),
    to_unsigned(380113669,32),
    to_unsigned(380316304,32),
    to_unsigned(380518935,32),
    to_unsigned(380721562,32),
    to_unsigned(380924187,32),
    to_unsigned(381126807,32),
    to_unsigned(381329425,32),
    to_unsigned(381532038,32),
    to_unsigned(381734649,32),
    to_unsigned(381937255,32),
    to_unsigned(382139859,32),
    to_unsigned(382342458,32),
    to_unsigned(382545054,32),
    to_unsigned(382747647,32),
    to_unsigned(382950236,32),
    to_unsigned(383152822,32),
    to_unsigned(383355404,32),
    to_unsigned(383557982,32),
    to_unsigned(383760557,32),
    to_unsigned(383963129,32),
    to_unsigned(384165697,32),
    to_unsigned(384368261,32),
    to_unsigned(384570822,32),
    to_unsigned(384773380,32),
    to_unsigned(384975934,32),
    to_unsigned(385178484,32),
    to_unsigned(385381031,32),
    to_unsigned(385583574,32),
    to_unsigned(385786114,32),
    to_unsigned(385988650,32),
    to_unsigned(386191182,32),
    to_unsigned(386393711,32),
    to_unsigned(386596237,32),
    to_unsigned(386798759,32),
    to_unsigned(387001277,32),
    to_unsigned(387203792,32),
    to_unsigned(387406303,32),
    to_unsigned(387608811,32),
    to_unsigned(387811315,32),
    to_unsigned(388013816,32),
    to_unsigned(388216313,32),
    to_unsigned(388418806,32),
    to_unsigned(388621296,32),
    to_unsigned(388823782,32),
    to_unsigned(389026265,32),
    to_unsigned(389228744,32),
    to_unsigned(389431220,32),
    to_unsigned(389633692,32),
    to_unsigned(389836160,32),
    to_unsigned(390038625,32),
    to_unsigned(390241086,32),
    to_unsigned(390443544,32),
    to_unsigned(390645998,32),
    to_unsigned(390848448,32),
    to_unsigned(391050895,32),
    to_unsigned(391253339,32),
    to_unsigned(391455778,32),
    to_unsigned(391658214,32),
    to_unsigned(391860647,32),
    to_unsigned(392063076,32),
    to_unsigned(392265501,32),
    to_unsigned(392467923,32),
    to_unsigned(392670341,32),
    to_unsigned(392872755,32),
    to_unsigned(393075166,32),
    to_unsigned(393277573,32),
    to_unsigned(393479977,32),
    to_unsigned(393682377,32),
    to_unsigned(393884773,32),
    to_unsigned(394087166,32),
    to_unsigned(394289555,32),
    to_unsigned(394491941,32),
    to_unsigned(394694323,32),
    to_unsigned(394896701,32),
    to_unsigned(395099076,32),
    to_unsigned(395301447,32),
    to_unsigned(395503814,32),
    to_unsigned(395706178,32),
    to_unsigned(395908538,32),
    to_unsigned(396110894,32),
    to_unsigned(396313247,32),
    to_unsigned(396515596,32),
    to_unsigned(396717942,32),
    to_unsigned(396920284,32),
    to_unsigned(397122622,32),
    to_unsigned(397324957,32),
    to_unsigned(397527288,32),
    to_unsigned(397729615,32),
    to_unsigned(397931938,32),
    to_unsigned(398134258,32),
    to_unsigned(398336575,32),
    to_unsigned(398538887,32),
    to_unsigned(398741196,32),
    to_unsigned(398943502,32),
    to_unsigned(399145803,32),
    to_unsigned(399348101,32),
    to_unsigned(399550396,32),
    to_unsigned(399752686,32),
    to_unsigned(399954973,32),
    to_unsigned(400157257,32),
    to_unsigned(400359536,32),
    to_unsigned(400561812,32),
    to_unsigned(400764084,32),
    to_unsigned(400966353,32),
    to_unsigned(401168618,32),
    to_unsigned(401370879,32),
    to_unsigned(401573136,32),
    to_unsigned(401775390,32),
    to_unsigned(401977640,32),
    to_unsigned(402179887,32),
    to_unsigned(402382130,32),
    to_unsigned(402584369,32),
    to_unsigned(402786604,32),
    to_unsigned(402988836,32),
    to_unsigned(403191063,32),
    to_unsigned(403393288,32),
    to_unsigned(403595508,32),
    to_unsigned(403797725,32),
    to_unsigned(403999938,32),
    to_unsigned(404202147,32),
    to_unsigned(404404353,32),
    to_unsigned(404606555,32),
    to_unsigned(404808753,32),
    to_unsigned(405010948,32),
    to_unsigned(405213139,32),
    to_unsigned(405415326,32),
    to_unsigned(405617509,32),
    to_unsigned(405819689,32),
    to_unsigned(406021864,32),
    to_unsigned(406224037,32),
    to_unsigned(406426205,32),
    to_unsigned(406628370,32),
    to_unsigned(406830531,32),
    to_unsigned(407032688,32),
    to_unsigned(407234841,32),
    to_unsigned(407436991,32),
    to_unsigned(407639137,32),
    to_unsigned(407841279,32),
    to_unsigned(408043418,32),
    to_unsigned(408245552,32),
    to_unsigned(408447683,32),
    to_unsigned(408649810,32),
    to_unsigned(408851934,32),
    to_unsigned(409054054,32),
    to_unsigned(409256170,32),
    to_unsigned(409458282,32),
    to_unsigned(409660390,32),
    to_unsigned(409862495,32),
    to_unsigned(410064596,32),
    to_unsigned(410266693,32),
    to_unsigned(410468786,32),
    to_unsigned(410670876,32),
    to_unsigned(410872961,32),
    to_unsigned(411075043,32),
    to_unsigned(411277122,32),
    to_unsigned(411479196,32),
    to_unsigned(411681267,32),
    to_unsigned(411883334,32),
    to_unsigned(412085397,32),
    to_unsigned(412287456,32),
    to_unsigned(412489512,32),
    to_unsigned(412691563,32),
    to_unsigned(412893611,32),
    to_unsigned(413095655,32),
    to_unsigned(413297696,32),
    to_unsigned(413499732,32),
    to_unsigned(413701765,32),
    to_unsigned(413903794,32),
    to_unsigned(414105819,32),
    to_unsigned(414307840,32),
    to_unsigned(414509858,32),
    to_unsigned(414711872,32),
    to_unsigned(414913882,32),
    to_unsigned(415115888,32),
    to_unsigned(415317890,32),
    to_unsigned(415519888,32),
    to_unsigned(415721883,32),
    to_unsigned(415923874,32),
    to_unsigned(416125861,32),
    to_unsigned(416327844,32),
    to_unsigned(416529823,32),
    to_unsigned(416731799,32),
    to_unsigned(416933771,32),
    to_unsigned(417135738,32),
    to_unsigned(417337702,32),
    to_unsigned(417539663,32),
    to_unsigned(417741619,32),
    to_unsigned(417943571,32),
    to_unsigned(418145520,32),
    to_unsigned(418347465,32),
    to_unsigned(418549406,32),
    to_unsigned(418751343,32),
    to_unsigned(418953276,32),
    to_unsigned(419155206,32),
    to_unsigned(419357131,32),
    to_unsigned(419559053,32),
    to_unsigned(419760971,32),
    to_unsigned(419962885,32),
    to_unsigned(420164795,32),
    to_unsigned(420366701,32),
    to_unsigned(420568604,32),
    to_unsigned(420770502,32),
    to_unsigned(420972397,32),
    to_unsigned(421174288,32),
    to_unsigned(421376175,32),
    to_unsigned(421578058,32),
    to_unsigned(421779937,32),
    to_unsigned(421981812,32),
    to_unsigned(422183684,32),
    to_unsigned(422385551,32),
    to_unsigned(422587415,32),
    to_unsigned(422789275,32),
    to_unsigned(422991130,32),
    to_unsigned(423192983,32),
    to_unsigned(423394831,32),
    to_unsigned(423596675,32),
    to_unsigned(423798515,32),
    to_unsigned(424000352,32),
    to_unsigned(424202184,32),
    to_unsigned(424404013,32),
    to_unsigned(424605838,32),
    to_unsigned(424807658,32),
    to_unsigned(425009475,32),
    to_unsigned(425211288,32),
    to_unsigned(425413098,32),
    to_unsigned(425614903,32),
    to_unsigned(425816704,32),
    to_unsigned(426018501,32),
    to_unsigned(426220295,32),
    to_unsigned(426422084,32),
    to_unsigned(426623870,32),
    to_unsigned(426825652,32),
    to_unsigned(427027430,32),
    to_unsigned(427229203,32),
    to_unsigned(427430973,32),
    to_unsigned(427632739,32),
    to_unsigned(427834501,32),
    to_unsigned(428036260,32),
    to_unsigned(428238014,32),
    to_unsigned(428439764,32),
    to_unsigned(428641510,32),
    to_unsigned(428843253,32),
    to_unsigned(429044991,32),
    to_unsigned(429246726,32),
    to_unsigned(429448456,32),
    to_unsigned(429650183,32),
    to_unsigned(429851906,32),
    to_unsigned(430053624,32),
    to_unsigned(430255339,32),
    to_unsigned(430457050,32),
    to_unsigned(430658757,32),
    to_unsigned(430860460,32),
    to_unsigned(431062159,32),
    to_unsigned(431263854,32),
    to_unsigned(431465545,32),
    to_unsigned(431667232,32),
    to_unsigned(431868915,32),
    to_unsigned(432070594,32),
    to_unsigned(432272269,32),
    to_unsigned(432473940,32),
    to_unsigned(432675607,32),
    to_unsigned(432877270,32),
    to_unsigned(433078930,32),
    to_unsigned(433280585,32),
    to_unsigned(433482236,32),
    to_unsigned(433683883,32),
    to_unsigned(433885527,32),
    to_unsigned(434087166,32),
    to_unsigned(434288801,32),
    to_unsigned(434490433,32),
    to_unsigned(434692060,32),
    to_unsigned(434893683,32),
    to_unsigned(435095303,32),
    to_unsigned(435296918,32),
    to_unsigned(435498529,32),
    to_unsigned(435700137,32),
    to_unsigned(435901740,32),
    to_unsigned(436103339,32),
    to_unsigned(436304935,32),
    to_unsigned(436506526,32),
    to_unsigned(436708113,32),
    to_unsigned(436909697,32),
    to_unsigned(437111276,32),
    to_unsigned(437312851,32),
    to_unsigned(437514422,32),
    to_unsigned(437715989,32),
    to_unsigned(437917553,32),
    to_unsigned(438119112,32),
    to_unsigned(438320667,32),
    to_unsigned(438522218,32),
    to_unsigned(438723765,32),
    to_unsigned(438925308,32),
    to_unsigned(439126847,32),
    to_unsigned(439328382,32),
    to_unsigned(439529913,32),
    to_unsigned(439731440,32),
    to_unsigned(439932963,32),
    to_unsigned(440134481,32),
    to_unsigned(440335996,32),
    to_unsigned(440537507,32),
    to_unsigned(440739014,32),
    to_unsigned(440940516,32),
    to_unsigned(441142015,32),
    to_unsigned(441343509,32),
    to_unsigned(441545000,32),
    to_unsigned(441746486,32),
    to_unsigned(441947968,32),
    to_unsigned(442149447,32),
    to_unsigned(442350921,32),
    to_unsigned(442552391,32),
    to_unsigned(442753857,32),
    to_unsigned(442955319,32),
    to_unsigned(443156777,32),
    to_unsigned(443358231,32),
    to_unsigned(443559681,32),
    to_unsigned(443761126,32),
    to_unsigned(443962568,32),
    to_unsigned(444164005,32),
    to_unsigned(444365439,32),
    to_unsigned(444566868,32),
    to_unsigned(444768293,32),
    to_unsigned(444969715,32),
    to_unsigned(445171132,32),
    to_unsigned(445372545,32),
    to_unsigned(445573954,32),
    to_unsigned(445775359,32),
    to_unsigned(445976759,32),
    to_unsigned(446178156,32),
    to_unsigned(446379548,32),
    to_unsigned(446580937,32),
    to_unsigned(446782321,32),
    to_unsigned(446983701,32),
    to_unsigned(447185077,32),
    to_unsigned(447386449,32),
    to_unsigned(447587817,32),
    to_unsigned(447789181,32),
    to_unsigned(447990541,32),
    to_unsigned(448191896,32),
    to_unsigned(448393248,32),
    to_unsigned(448594595,32),
    to_unsigned(448795938,32),
    to_unsigned(448997277,32),
    to_unsigned(449198612,32),
    to_unsigned(449399943,32),
    to_unsigned(449601269,32),
    to_unsigned(449802592,32),
    to_unsigned(450003910,32),
    to_unsigned(450205225,32),
    to_unsigned(450406535,32),
    to_unsigned(450607841,32),
    to_unsigned(450809143,32),
    to_unsigned(451010440,32),
    to_unsigned(451211734,32),
    to_unsigned(451413023,32),
    to_unsigned(451614308,32),
    to_unsigned(451815589,32),
    to_unsigned(452016866,32),
    to_unsigned(452218139,32),
    to_unsigned(452419408,32),
    to_unsigned(452620672,32),
    to_unsigned(452821933,32),
    to_unsigned(453023189,32),
    to_unsigned(453224441,32),
    to_unsigned(453425689,32),
    to_unsigned(453626932,32),
    to_unsigned(453828172,32),
    to_unsigned(454029407,32),
    to_unsigned(454230638,32),
    to_unsigned(454431865,32),
    to_unsigned(454633088,32),
    to_unsigned(454834306,32),
    to_unsigned(455035521,32),
    to_unsigned(455236731,32),
    to_unsigned(455437937,32),
    to_unsigned(455639139,32),
    to_unsigned(455840337,32),
    to_unsigned(456041530,32),
    to_unsigned(456242719,32),
    to_unsigned(456443905,32),
    to_unsigned(456645085,32),
    to_unsigned(456846262,32),
    to_unsigned(457047435,32),
    to_unsigned(457248603,32),
    to_unsigned(457449767,32),
    to_unsigned(457650927,32),
    to_unsigned(457852083,32),
    to_unsigned(458053234,32),
    to_unsigned(458254381,32),
    to_unsigned(458455525,32),
    to_unsigned(458656663,32),
    to_unsigned(458857798,32),
    to_unsigned(459058928,32),
    to_unsigned(459260055,32),
    to_unsigned(459461177,32),
    to_unsigned(459662294,32),
    to_unsigned(459863408,32),
    to_unsigned(460064517,32),
    to_unsigned(460265622,32),
    to_unsigned(460466723,32),
    to_unsigned(460667820,32),
    to_unsigned(460868912,32),
    to_unsigned(461070000,32),
    to_unsigned(461271084,32),
    to_unsigned(461472164,32),
    to_unsigned(461673239,32),
    to_unsigned(461874310,32),
    to_unsigned(462075377,32),
    to_unsigned(462276440,32),
    to_unsigned(462477498,32),
    to_unsigned(462678553,32),
    to_unsigned(462879603,32),
    to_unsigned(463080648,32),
    to_unsigned(463281690,32),
    to_unsigned(463482727,32),
    to_unsigned(463683760,32),
    to_unsigned(463884788,32),
    to_unsigned(464085813,32),
    to_unsigned(464286833,32),
    to_unsigned(464487849,32),
    to_unsigned(464688860,32),
    to_unsigned(464889868,32),
    to_unsigned(465090871,32),
    to_unsigned(465291869,32),
    to_unsigned(465492864,32),
    to_unsigned(465693854,32),
    to_unsigned(465894840,32),
    to_unsigned(466095822,32),
    to_unsigned(466296799,32),
    to_unsigned(466497772,32),
    to_unsigned(466698741,32),
    to_unsigned(466899705,32),
    to_unsigned(467100665,32),
    to_unsigned(467301621,32),
    to_unsigned(467502573,32),
    to_unsigned(467703520,32),
    to_unsigned(467904463,32),
    to_unsigned(468105402,32),
    to_unsigned(468306336,32),
    to_unsigned(468507266,32),
    to_unsigned(468708192,32),
    to_unsigned(468909114,32),
    to_unsigned(469110031,32),
    to_unsigned(469310944,32),
    to_unsigned(469511852,32),
    to_unsigned(469712757,32),
    to_unsigned(469913656,32),
    to_unsigned(470114552,32),
    to_unsigned(470315443,32),
    to_unsigned(470516330,32),
    to_unsigned(470717213,32),
    to_unsigned(470918091,32),
    to_unsigned(471118965,32),
    to_unsigned(471319835,32),
    to_unsigned(471520700,32),
    to_unsigned(471721561,32),
    to_unsigned(471922418,32),
    to_unsigned(472123270,32),
    to_unsigned(472324118,32),
    to_unsigned(472524962,32),
    to_unsigned(472725801,32),
    to_unsigned(472926636,32),
    to_unsigned(473127466,32),
    to_unsigned(473328293,32),
    to_unsigned(473529115,32),
    to_unsigned(473729932,32),
    to_unsigned(473930745,32),
    to_unsigned(474131554,32),
    to_unsigned(474332359,32),
    to_unsigned(474533159,32),
    to_unsigned(474733954,32),
    to_unsigned(474934746,32),
    to_unsigned(475135533,32),
    to_unsigned(475336315,32),
    to_unsigned(475537094,32),
    to_unsigned(475737868,32),
    to_unsigned(475938637,32),
    to_unsigned(476139402,32),
    to_unsigned(476340163,32),
    to_unsigned(476540919,32),
    to_unsigned(476741672,32),
    to_unsigned(476942419,32),
    to_unsigned(477143162,32),
    to_unsigned(477343901,32),
    to_unsigned(477544636,32),
    to_unsigned(477745366,32),
    to_unsigned(477946092,32),
    to_unsigned(478146813,32),
    to_unsigned(478347530,32),
    to_unsigned(478548242,32),
    to_unsigned(478748950,32),
    to_unsigned(478949654,32),
    to_unsigned(479150353,32),
    to_unsigned(479351048,32),
    to_unsigned(479551739,32),
    to_unsigned(479752425,32),
    to_unsigned(479953107,32),
    to_unsigned(480153784,32),
    to_unsigned(480354457,32),
    to_unsigned(480555125,32),
    to_unsigned(480755789,32),
    to_unsigned(480956449,32),
    to_unsigned(481157104,32),
    to_unsigned(481357755,32),
    to_unsigned(481558401,32),
    to_unsigned(481759043,32),
    to_unsigned(481959681,32),
    to_unsigned(482160314,32),
    to_unsigned(482360942,32),
    to_unsigned(482561566,32),
    to_unsigned(482762186,32),
    to_unsigned(482962802,32),
    to_unsigned(483163412,32),
    to_unsigned(483364019,32),
    to_unsigned(483564621,32),
    to_unsigned(483765218,32),
    to_unsigned(483965811,32),
    to_unsigned(484166400,32),
    to_unsigned(484366984,32),
    to_unsigned(484567564,32),
    to_unsigned(484768139,32),
    to_unsigned(484968710,32),
    to_unsigned(485169277,32),
    to_unsigned(485369839,32),
    to_unsigned(485570396,32),
    to_unsigned(485770949,32),
    to_unsigned(485971498,32),
    to_unsigned(486172042,32),
    to_unsigned(486372581,32),
    to_unsigned(486573116,32),
    to_unsigned(486773647,32),
    to_unsigned(486974173,32),
    to_unsigned(487174695,32),
    to_unsigned(487375212,32),
    to_unsigned(487575725,32),
    to_unsigned(487776233,32),
    to_unsigned(487976737,32),
    to_unsigned(488177236,32),
    to_unsigned(488377731,32),
    to_unsigned(488578221,32),
    to_unsigned(488778707,32),
    to_unsigned(488979189,32),
    to_unsigned(489179665,32),
    to_unsigned(489380138,32),
    to_unsigned(489580606,32),
    to_unsigned(489781069,32),
    to_unsigned(489981528,32),
    to_unsigned(490181982,32),
    to_unsigned(490382432,32),
    to_unsigned(490582877,32),
    to_unsigned(490783318,32),
    to_unsigned(490983754,32),
    to_unsigned(491184186,32),
    to_unsigned(491384614,32),
    to_unsigned(491585036,32),
    to_unsigned(491785455,32),
    to_unsigned(491985868,32),
    to_unsigned(492186277,32),
    to_unsigned(492386682,32),
    to_unsigned(492587082,32),
    to_unsigned(492787478,32),
    to_unsigned(492987869,32),
    to_unsigned(493188256,32),
    to_unsigned(493388638,32),
    to_unsigned(493589015,32),
    to_unsigned(493789388,32),
    to_unsigned(493989756,32),
    to_unsigned(494190120,32),
    to_unsigned(494390480,32),
    to_unsigned(494590835,32),
    to_unsigned(494791185,32),
    to_unsigned(494991530,32),
    to_unsigned(495191872,32),
    to_unsigned(495392208,32),
    to_unsigned(495592540,32),
    to_unsigned(495792868,32),
    to_unsigned(495993191,32),
    to_unsigned(496193509,32),
    to_unsigned(496393823,32),
    to_unsigned(496594132,32),
    to_unsigned(496794437,32),
    to_unsigned(496994737,32),
    to_unsigned(497195032,32),
    to_unsigned(497395323,32),
    to_unsigned(497595610,32),
    to_unsigned(497795892,32),
    to_unsigned(497996169,32),
    to_unsigned(498196442,32),
    to_unsigned(498396710,32),
    to_unsigned(498596973,32),
    to_unsigned(498797232,32),
    to_unsigned(498997487,32),
    to_unsigned(499197736,32),
    to_unsigned(499397981,32),
    to_unsigned(499598222,32),
    to_unsigned(499798458,32),
    to_unsigned(499998689,32),
    to_unsigned(500198916,32),
    to_unsigned(500399138,32),
    to_unsigned(500599356,32),
    to_unsigned(500799569,32),
    to_unsigned(500999777,32),
    to_unsigned(501199981,32),
    to_unsigned(501400180,32),
    to_unsigned(501600375,32),
    to_unsigned(501800565,32),
    to_unsigned(502000750,32),
    to_unsigned(502200931,32),
    to_unsigned(502401107,32),
    to_unsigned(502601279,32),
    to_unsigned(502801446,32),
    to_unsigned(503001608,32),
    to_unsigned(503201766,32),
    to_unsigned(503401919,32),
    to_unsigned(503602067,32),
    to_unsigned(503802211,32),
    to_unsigned(504002350,32),
    to_unsigned(504202484,32),
    to_unsigned(504402614,32),
    to_unsigned(504602739,32),
    to_unsigned(504802860,32),
    to_unsigned(505002976,32),
    to_unsigned(505203087,32),
    to_unsigned(505403194,32),
    to_unsigned(505603296,32),
    to_unsigned(505803393,32),
    to_unsigned(506003486,32),
    to_unsigned(506203574,32),
    to_unsigned(506403658,32),
    to_unsigned(506603736,32),
    to_unsigned(506803810,32),
    to_unsigned(507003880,32),
    to_unsigned(507203945,32),
    to_unsigned(507404005,32),
    to_unsigned(507604060,32),
    to_unsigned(507804111,32),
    to_unsigned(508004157,32),
    to_unsigned(508204199,32),
    to_unsigned(508404236,32),
    to_unsigned(508604268,32),
    to_unsigned(508804295,32),
    to_unsigned(509004318,32),
    to_unsigned(509204336,32),
    to_unsigned(509404349,32),
    to_unsigned(509604358,32),
    to_unsigned(509804362,32),
    to_unsigned(510004361,32),
    to_unsigned(510204356,32),
    to_unsigned(510404346,32),
    to_unsigned(510604331,32),
    to_unsigned(510804312,32),
    to_unsigned(511004288,32),
    to_unsigned(511204259,32),
    to_unsigned(511404226,32),
    to_unsigned(511604187,32),
    to_unsigned(511804144,32),
    to_unsigned(512004097,32),
    to_unsigned(512204045,32),
    to_unsigned(512403987,32),
    to_unsigned(512603926,32),
    to_unsigned(512803859,32),
    to_unsigned(513003788,32),
    to_unsigned(513203712,32),
    to_unsigned(513403632,32),
    to_unsigned(513603546,32),
    to_unsigned(513803456,32),
    to_unsigned(514003362,32),
    to_unsigned(514203262,32),
    to_unsigned(514403158,32),
    to_unsigned(514603049,32),
    to_unsigned(514802935,32),
    to_unsigned(515002817,32),
    to_unsigned(515202694,32),
    to_unsigned(515402566,32),
    to_unsigned(515602433,32),
    to_unsigned(515802296,32),
    to_unsigned(516002154,32),
    to_unsigned(516202007,32),
    to_unsigned(516401856,32),
    to_unsigned(516601699,32),
    to_unsigned(516801538,32),
    to_unsigned(517001372,32),
    to_unsigned(517201202,32),
    to_unsigned(517401026,32),
    to_unsigned(517600846,32),
    to_unsigned(517800662,32),
    to_unsigned(518000472,32),
    to_unsigned(518200278,32),
    to_unsigned(518400078,32),
    to_unsigned(518599875,32),
    to_unsigned(518799666,32),
    to_unsigned(518999453,32),
    to_unsigned(519199234,32),
    to_unsigned(519399011,32),
    to_unsigned(519598784,32),
    to_unsigned(519798551,32),
    to_unsigned(519998314,32),
    to_unsigned(520198072,32),
    to_unsigned(520397825,32),
    to_unsigned(520597573,32),
    to_unsigned(520797317,32),
    to_unsigned(520997056,32),
    to_unsigned(521196790,32),
    to_unsigned(521396519,32),
    to_unsigned(521596243,32),
    to_unsigned(521795963,32),
    to_unsigned(521995678,32),
    to_unsigned(522195388,32),
    to_unsigned(522395093,32),
    to_unsigned(522594793,32),
    to_unsigned(522794489,32),
    to_unsigned(522994180,32),
    to_unsigned(523193866,32),
    to_unsigned(523393547,32),
    to_unsigned(523593223,32),
    to_unsigned(523792895,32),
    to_unsigned(523992562,32),
    to_unsigned(524192224,32),
    to_unsigned(524391881,32),
    to_unsigned(524591533,32),
    to_unsigned(524791181,32),
    to_unsigned(524990823,32),
    to_unsigned(525190461,32),
    to_unsigned(525390094,32),
    to_unsigned(525589722,32),
    to_unsigned(525789346,32),
    to_unsigned(525988964,32),
    to_unsigned(526188578,32),
    to_unsigned(526388187,32),
    to_unsigned(526587791,32),
    to_unsigned(526787390,32),
    to_unsigned(526986984,32),
    to_unsigned(527186574,32),
    to_unsigned(527386158,32),
    to_unsigned(527585738,32),
    to_unsigned(527785313,32),
    to_unsigned(527984883,32),
    to_unsigned(528184448,32),
    to_unsigned(528384009,32),
    to_unsigned(528583564,32),
    to_unsigned(528783115,32),
    to_unsigned(528982661,32),
    to_unsigned(529182202,32),
    to_unsigned(529381738,32),
    to_unsigned(529581269,32),
    to_unsigned(529780795,32),
    to_unsigned(529980317,32),
    to_unsigned(530179834,32),
    to_unsigned(530379345,32),
    to_unsigned(530578852,32),
    to_unsigned(530778354,32),
    to_unsigned(530977851,32),
    to_unsigned(531177343,32),
    to_unsigned(531376831,32),
    to_unsigned(531576313,32),
    to_unsigned(531775791,32),
    to_unsigned(531975263,32),
    to_unsigned(532174731,32),
    to_unsigned(532374194,32),
    to_unsigned(532573652,32),
    to_unsigned(532773105,32),
    to_unsigned(532972553,32),
    to_unsigned(533171997,32),
    to_unsigned(533371435,32),
    to_unsigned(533570869,32),
    to_unsigned(533770297,32),
    to_unsigned(533969721,32),
    to_unsigned(534169140,32),
    to_unsigned(534368554,32),
    to_unsigned(534567963,32),
    to_unsigned(534767367,32),
    to_unsigned(534966766,32),
    to_unsigned(535166160,32),
    to_unsigned(535365549,32),
    to_unsigned(535564934,32),
    to_unsigned(535764313,32),
    to_unsigned(535963688,32),
    to_unsigned(536163057,32),
    to_unsigned(536362422,32),
    to_unsigned(536561782,32),
    to_unsigned(536761137,32),
    to_unsigned(536960486,32),
    to_unsigned(537159831,32),
    to_unsigned(537359171,32),
    to_unsigned(537558506,32),
    to_unsigned(537757837,32),
    to_unsigned(537957162,32),
    to_unsigned(538156482,32),
    to_unsigned(538355797,32),
    to_unsigned(538555108,32),
    to_unsigned(538754413,32),
    to_unsigned(538953714,32),
    to_unsigned(539153009,32),
    to_unsigned(539352300,32),
    to_unsigned(539551585,32),
    to_unsigned(539750866,32),
    to_unsigned(539950141,32),
    to_unsigned(540149412,32),
    to_unsigned(540348678,32),
    to_unsigned(540547939,32),
    to_unsigned(540747194,32),
    to_unsigned(540946445,32),
    to_unsigned(541145691,32),
    to_unsigned(541344932,32),
    to_unsigned(541544168,32),
    to_unsigned(541743399,32),
    to_unsigned(541942625,32),
    to_unsigned(542141846,32),
    to_unsigned(542341062,32),
    to_unsigned(542540273,32),
    to_unsigned(542739479,32),
    to_unsigned(542938680,32),
    to_unsigned(543137876,32),
    to_unsigned(543337067,32),
    to_unsigned(543536253,32),
    to_unsigned(543735434,32),
    to_unsigned(543934610,32),
    to_unsigned(544133781,32),
    to_unsigned(544332947,32),
    to_unsigned(544532108,32),
    to_unsigned(544731264,32),
    to_unsigned(544930415,32),
    to_unsigned(545129561,32),
    to_unsigned(545328702,32),
    to_unsigned(545527838,32),
    to_unsigned(545726969,32),
    to_unsigned(545926095,32),
    to_unsigned(546125216,32),
    to_unsigned(546324332,32),
    to_unsigned(546523443,32),
    to_unsigned(546722549,32),
    to_unsigned(546921650,32),
    to_unsigned(547120745,32),
    to_unsigned(547319836,32),
    to_unsigned(547518922,32),
    to_unsigned(547718003,32),
    to_unsigned(547917078,32),
    to_unsigned(548116149,32),
    to_unsigned(548315215,32),
    to_unsigned(548514275,32),
    to_unsigned(548713331,32),
    to_unsigned(548912381,32),
    to_unsigned(549111427,32),
    to_unsigned(549310467,32),
    to_unsigned(549509503,32),
    to_unsigned(549708533,32),
    to_unsigned(549907558,32),
    to_unsigned(550106578,32),
    to_unsigned(550305593,32),
    to_unsigned(550504604,32),
    to_unsigned(550703609,32),
    to_unsigned(550902609,32),
    to_unsigned(551101603,32),
    to_unsigned(551300593,32),
    to_unsigned(551499578,32),
    to_unsigned(551698558,32),
    to_unsigned(551897532,32),
    to_unsigned(552096502,32),
    to_unsigned(552295466,32),
    to_unsigned(552494426,32),
    to_unsigned(552693380,32),
    to_unsigned(552892329,32),
    to_unsigned(553091274,32),
    to_unsigned(553290213,32),
    to_unsigned(553489147,32),
    to_unsigned(553688076,32),
    to_unsigned(553886999,32),
    to_unsigned(554085918,32),
    to_unsigned(554284832,32),
    to_unsigned(554483740,32),
    to_unsigned(554682644,32),
    to_unsigned(554881542,32),
    to_unsigned(555080435,32),
    to_unsigned(555279323,32),
    to_unsigned(555478207,32),
    to_unsigned(555677084,32),
    to_unsigned(555875957,32),
    to_unsigned(556074825,32),
    to_unsigned(556273688,32),
    to_unsigned(556472545,32),
    to_unsigned(556671397,32),
    to_unsigned(556870245,32),
    to_unsigned(557069087,32),
    to_unsigned(557267924,32),
    to_unsigned(557466756,32),
    to_unsigned(557665583,32),
    to_unsigned(557864404,32),
    to_unsigned(558063221,32),
    to_unsigned(558262032,32),
    to_unsigned(558460838,32),
    to_unsigned(558659639,32),
    to_unsigned(558858435,32),
    to_unsigned(559057226,32),
    to_unsigned(559256012,32),
    to_unsigned(559454793,32),
    to_unsigned(559653568,32),
    to_unsigned(559852338,32),
    to_unsigned(560051103,32),
    to_unsigned(560249863,32),
    to_unsigned(560448618,32),
    to_unsigned(560647368,32),
    to_unsigned(560846113,32),
    to_unsigned(561044852,32),
    to_unsigned(561243586,32),
    to_unsigned(561442315,32),
    to_unsigned(561641039,32),
    to_unsigned(561839758,32),
    to_unsigned(562038471,32),
    to_unsigned(562237180,32),
    to_unsigned(562435883,32),
    to_unsigned(562634581,32),
    to_unsigned(562833274,32),
    to_unsigned(563031962,32),
    to_unsigned(563230644,32),
    to_unsigned(563429322,32),
    to_unsigned(563627994,32),
    to_unsigned(563826661,32),
    to_unsigned(564025323,32),
    to_unsigned(564223979,32),
    to_unsigned(564422631,32),
    to_unsigned(564621277,32),
    to_unsigned(564819918,32),
    to_unsigned(565018554,32),
    to_unsigned(565217185,32),
    to_unsigned(565415810,32),
    to_unsigned(565614431,32),
    to_unsigned(565813046,32),
    to_unsigned(566011656,32),
    to_unsigned(566210260,32),
    to_unsigned(566408860,32),
    to_unsigned(566607454,32),
    to_unsigned(566806043,32),
    to_unsigned(567004627,32),
    to_unsigned(567203206,32),
    to_unsigned(567401779,32),
    to_unsigned(567600348,32),
    to_unsigned(567798911,32),
    to_unsigned(567997468,32),
    to_unsigned(568196021,32),
    to_unsigned(568394568,32),
    to_unsigned(568593110,32),
    to_unsigned(568791647,32),
    to_unsigned(568990179,32),
    to_unsigned(569188705,32),
    to_unsigned(569387227,32),
    to_unsigned(569585743,32),
    to_unsigned(569784253,32),
    to_unsigned(569982759,32),
    to_unsigned(570181259,32),
    to_unsigned(570379754,32),
    to_unsigned(570578244,32),
    to_unsigned(570776729,32),
    to_unsigned(570975208,32),
    to_unsigned(571173682,32),
    to_unsigned(571372151,32),
    to_unsigned(571570614,32),
    to_unsigned(571769073,32),
    to_unsigned(571967526,32),
    to_unsigned(572165973,32),
    to_unsigned(572364416,32),
    to_unsigned(572562853,32),
    to_unsigned(572761285,32),
    to_unsigned(572959712,32),
    to_unsigned(573158133,32),
    to_unsigned(573356550,32),
    to_unsigned(573554960,32),
    to_unsigned(573753366,32),
    to_unsigned(573951766,32),
    to_unsigned(574150162,32),
    to_unsigned(574348551,32),
    to_unsigned(574546936,32),
    to_unsigned(574745315,32),
    to_unsigned(574943689,32),
    to_unsigned(575142058,32),
    to_unsigned(575340421,32),
    to_unsigned(575538779,32),
    to_unsigned(575737132,32),
    to_unsigned(575935480,32),
    to_unsigned(576133822,32),
    to_unsigned(576332159,32),
    to_unsigned(576530491,32),
    to_unsigned(576728817,32),
    to_unsigned(576927138,32),
    to_unsigned(577125454,32),
    to_unsigned(577323764,32),
    to_unsigned(577522069,32),
    to_unsigned(577720369,32),
    to_unsigned(577918664,32),
    to_unsigned(578116953,32),
    to_unsigned(578315237,32),
    to_unsigned(578513515,32),
    to_unsigned(578711789,32),
    to_unsigned(578910057,32),
    to_unsigned(579108319,32),
    to_unsigned(579306577,32),
    to_unsigned(579504829,32),
    to_unsigned(579703075,32),
    to_unsigned(579901317,32),
    to_unsigned(580099553,32),
    to_unsigned(580297783,32),
    to_unsigned(580496008,32),
    to_unsigned(580694228,32),
    to_unsigned(580892443,32),
    to_unsigned(581090652,32),
    to_unsigned(581288856,32),
    to_unsigned(581487055,32),
    to_unsigned(581685248,32),
    to_unsigned(581883436,32),
    to_unsigned(582081619,32),
    to_unsigned(582279796,32),
    to_unsigned(582477968,32),
    to_unsigned(582676134,32),
    to_unsigned(582874296,32),
    to_unsigned(583072451,32),
    to_unsigned(583270602,32),
    to_unsigned(583468747,32),
    to_unsigned(583666887,32),
    to_unsigned(583865021,32),
    to_unsigned(584063150,32),
    to_unsigned(584261274,32),
    to_unsigned(584459392,32),
    to_unsigned(584657505,32),
    to_unsigned(584855612,32),
    to_unsigned(585053715,32),
    to_unsigned(585251811,32),
    to_unsigned(585449903,32),
    to_unsigned(585647989,32),
    to_unsigned(585846069,32),
    to_unsigned(586044144,32),
    to_unsigned(586242214,32),
    to_unsigned(586440279,32),
    to_unsigned(586638338,32),
    to_unsigned(586836392,32),
    to_unsigned(587034440,32),
    to_unsigned(587232483,32),
    to_unsigned(587430520,32),
    to_unsigned(587628552,32),
    to_unsigned(587826579,32),
    to_unsigned(588024600,32),
    to_unsigned(588222616,32),
    to_unsigned(588420627,32),
    to_unsigned(588618632,32),
    to_unsigned(588816631,32),
    to_unsigned(589014626,32),
    to_unsigned(589212614,32),
    to_unsigned(589410598,32),
    to_unsigned(589608576,32),
    to_unsigned(589806548,32),
    to_unsigned(590004515,32),
    to_unsigned(590202477,32),
    to_unsigned(590400433,32),
    to_unsigned(590598384,32),
    to_unsigned(590796330,32),
    to_unsigned(590994270,32),
    to_unsigned(591192204,32),
    to_unsigned(591390134,32),
    to_unsigned(591588057,32),
    to_unsigned(591785976,32),
    to_unsigned(591983888,32),
    to_unsigned(592181796,32),
    to_unsigned(592379698,32),
    to_unsigned(592577594,32),
    to_unsigned(592775485,32),
    to_unsigned(592973371,32),
    to_unsigned(593171251,32),
    to_unsigned(593369126,32),
    to_unsigned(593566995,32),
    to_unsigned(593764859,32),
    to_unsigned(593962717,32),
    to_unsigned(594160570,32),
    to_unsigned(594358417,32),
    to_unsigned(594556259,32),
    to_unsigned(594754096,32),
    to_unsigned(594951927,32),
    to_unsigned(595149752,32),
    to_unsigned(595347573,32),
    to_unsigned(595545387,32),
    to_unsigned(595743196,32),
    to_unsigned(595941000,32),
    to_unsigned(596138798,32),
    to_unsigned(596336591,32),
    to_unsigned(596534378,32),
    to_unsigned(596732160,32),
    to_unsigned(596929936,32),
    to_unsigned(597127707,32),
    to_unsigned(597325472,32),
    to_unsigned(597523232,32),
    to_unsigned(597720986,32),
    to_unsigned(597918735,32),
    to_unsigned(598116478,32),
    to_unsigned(598314216,32),
    to_unsigned(598511948,32),
    to_unsigned(598709675,32),
    to_unsigned(598907397,32),
    to_unsigned(599105112,32),
    to_unsigned(599302823,32),
    to_unsigned(599500527,32),
    to_unsigned(599698227,32),
    to_unsigned(599895920,32),
    to_unsigned(600093609,32),
    to_unsigned(600291291,32),
    to_unsigned(600488969,32),
    to_unsigned(600686640,32),
    to_unsigned(600884307,32),
    to_unsigned(601081967,32),
    to_unsigned(601279622,32),
    to_unsigned(601477272,32),
    to_unsigned(601674916,32),
    to_unsigned(601872554,32),
    to_unsigned(602070188,32),
    to_unsigned(602267815,32),
    to_unsigned(602465437,32),
    to_unsigned(602663053,32),
    to_unsigned(602860664,32),
    to_unsigned(603058269,32),
    to_unsigned(603255869,32),
    to_unsigned(603453463,32),
    to_unsigned(603651052,32),
    to_unsigned(603848635,32),
    to_unsigned(604046213,32),
    to_unsigned(604243785,32),
    to_unsigned(604441351,32),
    to_unsigned(604638912,32),
    to_unsigned(604836468,32),
    to_unsigned(605034017,32),
    to_unsigned(605231562,32),
    to_unsigned(605429100,32),
    to_unsigned(605626634,32),
    to_unsigned(605824161,32),
    to_unsigned(606021683,32),
    to_unsigned(606219199,32),
    to_unsigned(606416710,32),
    to_unsigned(606614216,32),
    to_unsigned(606811715,32),
    to_unsigned(607009209,32),
    to_unsigned(607206698,32),
    to_unsigned(607404181,32),
    to_unsigned(607601658,32),
    to_unsigned(607799130,32),
    to_unsigned(607996596,32),
    to_unsigned(608194057,32),
    to_unsigned(608391512,32),
    to_unsigned(608588961,32),
    to_unsigned(608786405,32),
    to_unsigned(608983843,32),
    to_unsigned(609181276,32),
    to_unsigned(609378703,32),
    to_unsigned(609576124,32),
    to_unsigned(609773540,32),
    to_unsigned(609970950,32),
    to_unsigned(610168355,32),
    to_unsigned(610365754,32),
    to_unsigned(610563147,32),
    to_unsigned(610760535,32),
    to_unsigned(610957917,32),
    to_unsigned(611155294,32),
    to_unsigned(611352665,32),
    to_unsigned(611550030,32),
    to_unsigned(611747390,32),
    to_unsigned(611944744,32),
    to_unsigned(612142092,32),
    to_unsigned(612339435,32),
    to_unsigned(612536772,32),
    to_unsigned(612734104,32),
    to_unsigned(612931430,32),
    to_unsigned(613128750,32),
    to_unsigned(613326065,32),
    to_unsigned(613523374,32),
    to_unsigned(613720677,32),
    to_unsigned(613917975,32),
    to_unsigned(614115267,32),
    to_unsigned(614312554,32),
    to_unsigned(614509834,32),
    to_unsigned(614707110,32),
    to_unsigned(614904379,32),
    to_unsigned(615101643,32),
    to_unsigned(615298901,32),
    to_unsigned(615496154,32),
    to_unsigned(615693401,32),
    to_unsigned(615890642,32),
    to_unsigned(616087877,32),
    to_unsigned(616285107,32),
    to_unsigned(616482332,32),
    to_unsigned(616679550,32),
    to_unsigned(616876763,32),
    to_unsigned(617073970,32),
    to_unsigned(617271172,32),
    to_unsigned(617468368,32),
    to_unsigned(617665558,32),
    to_unsigned(617862743,32),
    to_unsigned(618059921,32),
    to_unsigned(618257095,32),
    to_unsigned(618454262,32),
    to_unsigned(618651424,32),
    to_unsigned(618848580,32),
    to_unsigned(619045731,32),
    to_unsigned(619242875,32),
    to_unsigned(619440014,32),
    to_unsigned(619637148,32),
    to_unsigned(619834275,32),
    to_unsigned(620031397,32),
    to_unsigned(620228514,32),
    to_unsigned(620425624,32),
    to_unsigned(620622729,32),
    to_unsigned(620819828,32),
    to_unsigned(621016922,32),
    to_unsigned(621214009,32),
    to_unsigned(621411091,32),
    to_unsigned(621608168,32),
    to_unsigned(621805238,32),
    to_unsigned(622002303,32),
    to_unsigned(622199362,32),
    to_unsigned(622396416,32),
    to_unsigned(622593464,32),
    to_unsigned(622790506,32),
    to_unsigned(622987542,32),
    to_unsigned(623184573,32),
    to_unsigned(623381597,32),
    to_unsigned(623578616,32),
    to_unsigned(623775630,32),
    to_unsigned(623972638,32),
    to_unsigned(624169639,32),
    to_unsigned(624366636,32),
    to_unsigned(624563626,32),
    to_unsigned(624760611,32),
    to_unsigned(624957590,32),
    to_unsigned(625154563,32),
    to_unsigned(625351530,32),
    to_unsigned(625548492,32),
    to_unsigned(625745448,32),
    to_unsigned(625942398,32),
    to_unsigned(626139343,32),
    to_unsigned(626336281,32),
    to_unsigned(626533214,32),
    to_unsigned(626730141,32),
    to_unsigned(626927063,32),
    to_unsigned(627123979,32),
    to_unsigned(627320888,32),
    to_unsigned(627517793,32),
    to_unsigned(627714691,32),
    to_unsigned(627911584,32),
    to_unsigned(628108470,32),
    to_unsigned(628305351,32),
    to_unsigned(628502227,32),
    to_unsigned(628699096,32),
    to_unsigned(628895960,32),
    to_unsigned(629092818,32),
    to_unsigned(629289670,32),
    to_unsigned(629486516,32),
    to_unsigned(629683357,32),
    to_unsigned(629880192,32),
    to_unsigned(630077021,32),
    to_unsigned(630273844,32),
    to_unsigned(630470661,32),
    to_unsigned(630667473,32),
    to_unsigned(630864279,32),
    to_unsigned(631061079,32),
    to_unsigned(631257873,32),
    to_unsigned(631454661,32),
    to_unsigned(631651444,32),
    to_unsigned(631848221,32),
    to_unsigned(632044992,32),
    to_unsigned(632241757,32),
    to_unsigned(632438516,32),
    to_unsigned(632635270,32),
    to_unsigned(632832018,32),
    to_unsigned(633028760,32),
    to_unsigned(633225496,32),
    to_unsigned(633422226,32),
    to_unsigned(633618951,32),
    to_unsigned(633815669,32),
    to_unsigned(634012382,32),
    to_unsigned(634209089,32),
    to_unsigned(634405790,32),
    to_unsigned(634602486,32),
    to_unsigned(634799175,32),
    to_unsigned(634995859,32),
    to_unsigned(635192537,32),
    to_unsigned(635389209,32),
    to_unsigned(635585875,32),
    to_unsigned(635782535,32),
    to_unsigned(635979190,32),
    to_unsigned(636175838,32),
    to_unsigned(636372481,32),
    to_unsigned(636569118,32),
    to_unsigned(636765749,32),
    to_unsigned(636962374,32),
    to_unsigned(637158994,32),
    to_unsigned(637355607,32),
    to_unsigned(637552215,32),
    to_unsigned(637748816,32),
    to_unsigned(637945412,32),
    to_unsigned(638142002,32),
    to_unsigned(638338587,32),
    to_unsigned(638535165,32),
    to_unsigned(638731737,32),
    to_unsigned(638928304,32),
    to_unsigned(639124865,32),
    to_unsigned(639321420,32),
    to_unsigned(639517969,32),
    to_unsigned(639714512,32),
    to_unsigned(639911049,32),
    to_unsigned(640107580,32),
    to_unsigned(640304106,32),
    to_unsigned(640500625,32),
    to_unsigned(640697139,32),
    to_unsigned(640893647,32),
    to_unsigned(641090149,32),
    to_unsigned(641286645,32),
    to_unsigned(641483135,32),
    to_unsigned(641679619,32),
    to_unsigned(641876097,32),
    to_unsigned(642072570,32),
    to_unsigned(642269036,32),
    to_unsigned(642465497,32),
    to_unsigned(642661951,32),
    to_unsigned(642858400,32),
    to_unsigned(643054843,32),
    to_unsigned(643251280,32),
    to_unsigned(643447711,32),
    to_unsigned(643644136,32),
    to_unsigned(643840556,32),
    to_unsigned(644036969,32),
    to_unsigned(644233376,32),
    to_unsigned(644429778,32),
    to_unsigned(644626173,32),
    to_unsigned(644822563,32),
    to_unsigned(645018947,32),
    to_unsigned(645215324,32),
    to_unsigned(645411696,32),
    to_unsigned(645608062,32),
    to_unsigned(645804422,32),
    to_unsigned(646000776,32),
    to_unsigned(646197124,32),
    to_unsigned(646393466,32),
    to_unsigned(646589803,32),
    to_unsigned(646786133,32),
    to_unsigned(646982457,32),
    to_unsigned(647178775,32),
    to_unsigned(647375088,32),
    to_unsigned(647571394,32),
    to_unsigned(647767695,32),
    to_unsigned(647963989,32),
    to_unsigned(648160278,32),
    to_unsigned(648356561,32),
    to_unsigned(648552837,32),
    to_unsigned(648749108,32),
    to_unsigned(648945373,32),
    to_unsigned(649141632,32),
    to_unsigned(649337885,32),
    to_unsigned(649534131,32),
    to_unsigned(649730372,32),
    to_unsigned(649926607,32),
    to_unsigned(650122836,32),
    to_unsigned(650319059,32),
    to_unsigned(650515276,32),
    to_unsigned(650711487,32),
    to_unsigned(650907692,32),
    to_unsigned(651103891,32),
    to_unsigned(651300084,32),
    to_unsigned(651496272,32),
    to_unsigned(651692453,32),
    to_unsigned(651888628,32),
    to_unsigned(652084797,32),
    to_unsigned(652280960,32),
    to_unsigned(652477117,32),
    to_unsigned(652673268,32),
    to_unsigned(652869413,32),
    to_unsigned(653065553,32),
    to_unsigned(653261686,32),
    to_unsigned(653457813,32),
    to_unsigned(653653934,32),
    to_unsigned(653850049,32),
    to_unsigned(654046158,32),
    to_unsigned(654242261,32),
    to_unsigned(654438358,32),
    to_unsigned(654634449,32),
    to_unsigned(654830534,32),
    to_unsigned(655026613,32),
    to_unsigned(655222686,32),
    to_unsigned(655418753,32),
    to_unsigned(655614814,32),
    to_unsigned(655810869,32),
    to_unsigned(656006918,32),
    to_unsigned(656202961,32),
    to_unsigned(656398998,32),
    to_unsigned(656595029,32),
    to_unsigned(656791053,32),
    to_unsigned(656987072,32),
    to_unsigned(657183085,32),
    to_unsigned(657379091,32),
    to_unsigned(657575092,32),
    to_unsigned(657771087,32),
    to_unsigned(657967075,32),
    to_unsigned(658163058,32),
    to_unsigned(658359034,32),
    to_unsigned(658555004,32),
    to_unsigned(658750969,32),
    to_unsigned(658946927,32),
    to_unsigned(659142879,32),
    to_unsigned(659338825,32),
    to_unsigned(659534765,32),
    to_unsigned(659730699,32),
    to_unsigned(659926627,32),
    to_unsigned(660122549,32),
    to_unsigned(660318465,32),
    to_unsigned(660514375,32),
    to_unsigned(660710279,32),
    to_unsigned(660906176,32),
    to_unsigned(661102068,32),
    to_unsigned(661297953,32),
    to_unsigned(661493833,32),
    to_unsigned(661689706,32),
    to_unsigned(661885573,32),
    to_unsigned(662081434,32),
    to_unsigned(662277289,32),
    to_unsigned(662473138,32),
    to_unsigned(662668981,32),
    to_unsigned(662864818,32),
    to_unsigned(663060649,32),
    to_unsigned(663256473,32),
    to_unsigned(663452292,32),
    to_unsigned(663648104,32),
    to_unsigned(663843910,32),
    to_unsigned(664039711,32),
    to_unsigned(664235505,32),
    to_unsigned(664431293,32),
    to_unsigned(664627075,32),
    to_unsigned(664822850,32),
    to_unsigned(665018620,32),
    to_unsigned(665214383,32),
    to_unsigned(665410141,32),
    to_unsigned(665605892,32),
    to_unsigned(665801637,32),
    to_unsigned(665997377,32),
    to_unsigned(666193109,32),
    to_unsigned(666388836,32),
    to_unsigned(666584557,32),
    to_unsigned(666780272,32),
    to_unsigned(666975980,32),
    to_unsigned(667171682,32),
    to_unsigned(667367379,32),
    to_unsigned(667563069,32),
    to_unsigned(667758753,32),
    to_unsigned(667954430,32),
    to_unsigned(668150102,32),
    to_unsigned(668345767,32),
    to_unsigned(668541427,32),
    to_unsigned(668737080,32),
    to_unsigned(668932727,32),
    to_unsigned(669128368,32),
    to_unsigned(669324003,32),
    to_unsigned(669519631,32),
    to_unsigned(669715254,32),
    to_unsigned(669910870,32),
    to_unsigned(670106480,32),
    to_unsigned(670302084,32),
    to_unsigned(670497682,32),
    to_unsigned(670693274,32),
    to_unsigned(670888859,32),
    to_unsigned(671084439,32),
    to_unsigned(671280012,32),
    to_unsigned(671475579,32),
    to_unsigned(671671140,32),
    to_unsigned(671866694,32),
    to_unsigned(672062243,32),
    to_unsigned(672257785,32),
    to_unsigned(672453321,32),
    to_unsigned(672648851,32),
    to_unsigned(672844375,32),
    to_unsigned(673039892,32),
    to_unsigned(673235404,32),
    to_unsigned(673430909,32),
    to_unsigned(673626408,32),
    to_unsigned(673821901,32),
    to_unsigned(674017387,32),
    to_unsigned(674212868,32),
    to_unsigned(674408342,32),
    to_unsigned(674603810,32),
    to_unsigned(674799272,32),
    to_unsigned(674994727,32),
    to_unsigned(675190177,32),
    to_unsigned(675385620,32),
    to_unsigned(675581057,32),
    to_unsigned(675776488,32),
    to_unsigned(675971912,32),
    to_unsigned(676167331,32),
    to_unsigned(676362743,32),
    to_unsigned(676558149,32),
    to_unsigned(676753549,32),
    to_unsigned(676948942,32),
    to_unsigned(677144329,32),
    to_unsigned(677339710,32),
    to_unsigned(677535085,32),
    to_unsigned(677730454,32),
    to_unsigned(677925816,32),
    to_unsigned(678121172,32),
    to_unsigned(678316522,32),
    to_unsigned(678511866,32),
    to_unsigned(678707203,32),
    to_unsigned(678902534,32),
    to_unsigned(679097859,32),
    to_unsigned(679293178,32),
    to_unsigned(679488491,32),
    to_unsigned(679683797,32),
    to_unsigned(679879097,32),
    to_unsigned(680074390,32),
    to_unsigned(680269678,32),
    to_unsigned(680464959,32),
    to_unsigned(680660234,32),
    to_unsigned(680855503,32),
    to_unsigned(681050765,32),
    to_unsigned(681246021,32),
    to_unsigned(681441271,32),
    to_unsigned(681636515,32),
    to_unsigned(681831752,32),
    to_unsigned(682026984,32),
    to_unsigned(682222208,32),
    to_unsigned(682417427,32),
    to_unsigned(682612639,32),
    to_unsigned(682807845,32),
    to_unsigned(683003045,32),
    to_unsigned(683198239,32),
    to_unsigned(683393426,32),
    to_unsigned(683588607,32),
    to_unsigned(683783781,32),
    to_unsigned(683978950,32),
    to_unsigned(684174112,32),
    to_unsigned(684369268,32),
    to_unsigned(684564417,32),
    to_unsigned(684759560,32),
    to_unsigned(684954697,32),
    to_unsigned(685149828,32),
    to_unsigned(685344952,32),
    to_unsigned(685540070,32),
    to_unsigned(685735182,32),
    to_unsigned(685930287,32),
    to_unsigned(686125386,32),
    to_unsigned(686320479,32),
    to_unsigned(686515566,32),
    to_unsigned(686710646,32),
    to_unsigned(686905720,32),
    to_unsigned(687100787,32),
    to_unsigned(687295848,32),
    to_unsigned(687490903,32),
    to_unsigned(687685952,32),
    to_unsigned(687880994,32),
    to_unsigned(688076030,32),
    to_unsigned(688271060,32),
    to_unsigned(688466083,32),
    to_unsigned(688661100,32),
    to_unsigned(688856111,32),
    to_unsigned(689051115,32),
    to_unsigned(689246113,32),
    to_unsigned(689441105,32),
    to_unsigned(689636090,32),
    to_unsigned(689831069,32),
    to_unsigned(690026042,32),
    to_unsigned(690221008,32),
    to_unsigned(690415968,32),
    to_unsigned(690610921,32),
    to_unsigned(690805869,32),
    to_unsigned(691000810,32),
    to_unsigned(691195744,32),
    to_unsigned(691390672,32),
    to_unsigned(691585594,32),
    to_unsigned(691780510,32),
    to_unsigned(691975419,32),
    to_unsigned(692170321,32),
    to_unsigned(692365218,32),
    to_unsigned(692560108,32),
    to_unsigned(692754992,32),
    to_unsigned(692949869,32),
    to_unsigned(693144740,32),
    to_unsigned(693339604,32),
    to_unsigned(693534463,32),
    to_unsigned(693729314,32),
    to_unsigned(693924160,32),
    to_unsigned(694118999,32),
    to_unsigned(694313832,32),
    to_unsigned(694508658,32),
    to_unsigned(694703478,32),
    to_unsigned(694898291,32),
    to_unsigned(695093098,32),
    to_unsigned(695287899,32),
    to_unsigned(695482694,32),
    to_unsigned(695677481,32),
    to_unsigned(695872263,32),
    to_unsigned(696067038,32),
    to_unsigned(696261807,32),
    to_unsigned(696456569,32),
    to_unsigned(696651325,32),
    to_unsigned(696846075,32),
    to_unsigned(697040818,32),
    to_unsigned(697235555,32),
    to_unsigned(697430285,32),
    to_unsigned(697625009,32),
    to_unsigned(697819727,32),
    to_unsigned(698014438,32),
    to_unsigned(698209142,32),
    to_unsigned(698403841,32),
    to_unsigned(698598533,32),
    to_unsigned(698793218,32),
    to_unsigned(698987897,32),
    to_unsigned(699182570,32),
    to_unsigned(699377236,32),
    to_unsigned(699571896,32),
    to_unsigned(699766549,32),
    to_unsigned(699961196,32),
    to_unsigned(700155836,32),
    to_unsigned(700350470,32),
    to_unsigned(700545098,32),
    to_unsigned(700739719,32),
    to_unsigned(700934334,32),
    to_unsigned(701128942,32),
    to_unsigned(701323544,32),
    to_unsigned(701518139,32),
    to_unsigned(701712728,32),
    to_unsigned(701907310,32),
    to_unsigned(702101886,32),
    to_unsigned(702296456,32),
    to_unsigned(702491019,32),
    to_unsigned(702685576,32),
    to_unsigned(702880126,32),
    to_unsigned(703074669,32),
    to_unsigned(703269207,32),
    to_unsigned(703463738,32),
    to_unsigned(703658262,32),
    to_unsigned(703852780,32),
    to_unsigned(704047291,32),
    to_unsigned(704241796,32),
    to_unsigned(704436294,32),
    to_unsigned(704630786,32),
    to_unsigned(704825272,32),
    to_unsigned(705019751,32),
    to_unsigned(705214223,32),
    to_unsigned(705408689,32),
    to_unsigned(705603149,32),
    to_unsigned(705797602,32),
    to_unsigned(705992049,32),
    to_unsigned(706186489,32),
    to_unsigned(706380922,32),
    to_unsigned(706575350,32),
    to_unsigned(706769770,32),
    to_unsigned(706964184,32),
    to_unsigned(707158592,32),
    to_unsigned(707352993,32),
    to_unsigned(707547388,32),
    to_unsigned(707741776,32),
    to_unsigned(707936157,32),
    to_unsigned(708130532,32),
    to_unsigned(708324901,32),
    to_unsigned(708519263,32),
    to_unsigned(708713619,32),
    to_unsigned(708907968,32),
    to_unsigned(709102310,32),
    to_unsigned(709296646,32),
    to_unsigned(709490976,32),
    to_unsigned(709685299,32),
    to_unsigned(709879615,32),
    to_unsigned(710073925,32),
    to_unsigned(710268229,32),
    to_unsigned(710462526,32),
    to_unsigned(710656816,32),
    to_unsigned(710851100,32),
    to_unsigned(711045377,32),
    to_unsigned(711239648,32),
    to_unsigned(711433912,32),
    to_unsigned(711628170,32),
    to_unsigned(711822421,32),
    to_unsigned(712016665,32),
    to_unsigned(712210903,32),
    to_unsigned(712405135,32),
    to_unsigned(712599360,32),
    to_unsigned(712793578,32),
    to_unsigned(712987790,32),
    to_unsigned(713181995,32),
    to_unsigned(713376194,32),
    to_unsigned(713570386,32),
    to_unsigned(713764572,32),
    to_unsigned(713958751,32),
    to_unsigned(714152924,32),
    to_unsigned(714347089,32),
    to_unsigned(714541249,32),
    to_unsigned(714735402,32),
    to_unsigned(714929548,32),
    to_unsigned(715123688,32),
    to_unsigned(715317821,32),
    to_unsigned(715511947,32),
    to_unsigned(715706067,32),
    to_unsigned(715900180,32),
    to_unsigned(716094287,32),
    to_unsigned(716288387,32),
    to_unsigned(716482481,32),
    to_unsigned(716676568,32),
    to_unsigned(716870648,32),
    to_unsigned(717064722,32),
    to_unsigned(717258790,32),
    to_unsigned(717452850,32),
    to_unsigned(717646904,32),
    to_unsigned(717840952,32),
    to_unsigned(718034993,32),
    to_unsigned(718229027,32),
    to_unsigned(718423055,32),
    to_unsigned(718617076,32),
    to_unsigned(718811090,32),
    to_unsigned(719005098,32),
    to_unsigned(719199099,32),
    to_unsigned(719393094,32),
    to_unsigned(719587082,32),
    to_unsigned(719781063,32),
    to_unsigned(719975038,32),
    to_unsigned(720169006,32),
    to_unsigned(720362968,32),
    to_unsigned(720556923,32),
    to_unsigned(720750871,32),
    to_unsigned(720944813,32),
    to_unsigned(721138748,32),
    to_unsigned(721332676,32),
    to_unsigned(721526598,32),
    to_unsigned(721720513,32),
    to_unsigned(721914422,32),
    to_unsigned(722108324,32),
    to_unsigned(722302219,32),
    to_unsigned(722496108,32),
    to_unsigned(722689990,32),
    to_unsigned(722883865,32),
    to_unsigned(723077734,32),
    to_unsigned(723271596,32),
    to_unsigned(723465451,32),
    to_unsigned(723659300,32),
    to_unsigned(723853142,32),
    to_unsigned(724046977,32),
    to_unsigned(724240806,32),
    to_unsigned(724434628,32),
    to_unsigned(724628444,32),
    to_unsigned(724822252,32),
    to_unsigned(725016055,32),
    to_unsigned(725209850,32),
    to_unsigned(725403639,32),
    to_unsigned(725597421,32),
    to_unsigned(725791197,32),
    to_unsigned(725984965,32),
    to_unsigned(726178728,32),
    to_unsigned(726372483,32),
    to_unsigned(726566232,32),
    to_unsigned(726759974,32),
    to_unsigned(726953709,32),
    to_unsigned(727147438,32),
    to_unsigned(727341160,32),
    to_unsigned(727534876,32),
    to_unsigned(727728584,32),
    to_unsigned(727922286,32),
    to_unsigned(728115982,32),
    to_unsigned(728309670,32),
    to_unsigned(728503352,32),
    to_unsigned(728697027,32),
    to_unsigned(728890696,32),
    to_unsigned(729084358,32),
    to_unsigned(729278013,32),
    to_unsigned(729471661,32),
    to_unsigned(729665303,32),
    to_unsigned(729858938,32),
    to_unsigned(730052566,32),
    to_unsigned(730246188,32),
    to_unsigned(730439803,32),
    to_unsigned(730633411,32),
    to_unsigned(730827012,32),
    to_unsigned(731020607,32),
    to_unsigned(731214195,32),
    to_unsigned(731407776,32),
    to_unsigned(731601351,32),
    to_unsigned(731794919,32),
    to_unsigned(731988480,32),
    to_unsigned(732182034,32),
    to_unsigned(732375582,32),
    to_unsigned(732569123,32),
    to_unsigned(732762657,32),
    to_unsigned(732956184,32),
    to_unsigned(733149705,32),
    to_unsigned(733343219,32),
    to_unsigned(733536726,32),
    to_unsigned(733730227,32),
    to_unsigned(733923721,32),
    to_unsigned(734117208,32),
    to_unsigned(734310688,32),
    to_unsigned(734504161,32),
    to_unsigned(734697628,32),
    to_unsigned(734891088,32),
    to_unsigned(735084541,32),
    to_unsigned(735277988,32),
    to_unsigned(735471428,32),
    to_unsigned(735664861,32),
    to_unsigned(735858287,32),
    to_unsigned(736051706,32),
    to_unsigned(736245119,32),
    to_unsigned(736438525,32),
    to_unsigned(736631924,32),
    to_unsigned(736825316,32),
    to_unsigned(737018702,32),
    to_unsigned(737212081,32),
    to_unsigned(737405453,32),
    to_unsigned(737598818,32),
    to_unsigned(737792177,32),
    to_unsigned(737985528,32),
    to_unsigned(738178873,32),
    to_unsigned(738372212,32),
    to_unsigned(738565543,32),
    to_unsigned(738758867,32),
    to_unsigned(738952185,32),
    to_unsigned(739145496,32),
    to_unsigned(739338800,32),
    to_unsigned(739532098,32),
    to_unsigned(739725388,32),
    to_unsigned(739918672,32),
    to_unsigned(740111949,32),
    to_unsigned(740305219,32),
    to_unsigned(740498483,32),
    to_unsigned(740691739,32),
    to_unsigned(740884989,32),
    to_unsigned(741078232,32),
    to_unsigned(741271468,32),
    to_unsigned(741464698,32),
    to_unsigned(741657920,32),
    to_unsigned(741851136,32),
    to_unsigned(742044345,32),
    to_unsigned(742237547,32),
    to_unsigned(742430742,32),
    to_unsigned(742623930,32),
    to_unsigned(742817112,32),
    to_unsigned(743010287,32),
    to_unsigned(743203455,32),
    to_unsigned(743396616,32),
    to_unsigned(743589770,32),
    to_unsigned(743782918,32),
    to_unsigned(743976058,32),
    to_unsigned(744169192,32),
    to_unsigned(744362319,32),
    to_unsigned(744555439,32),
    to_unsigned(744748552,32),
    to_unsigned(744941659,32),
    to_unsigned(745134758,32),
    to_unsigned(745327851,32),
    to_unsigned(745520937,32),
    to_unsigned(745714016,32),
    to_unsigned(745907088,32),
    to_unsigned(746100153,32),
    to_unsigned(746293211,32),
    to_unsigned(746486263,32),
    to_unsigned(746679308,32),
    to_unsigned(746872346,32),
    to_unsigned(747065377,32),
    to_unsigned(747258401,32),
    to_unsigned(747451418,32),
    to_unsigned(747644428,32),
    to_unsigned(747837432,32),
    to_unsigned(748030428,32),
    to_unsigned(748223418,32),
    to_unsigned(748416401,32),
    to_unsigned(748609377,32),
    to_unsigned(748802346,32),
    to_unsigned(748995308,32),
    to_unsigned(749188264,32),
    to_unsigned(749381212,32),
    to_unsigned(749574154,32),
    to_unsigned(749767088,32),
    to_unsigned(749960016,32),
    to_unsigned(750152937,32),
    to_unsigned(750345851,32),
    to_unsigned(750538758,32),
    to_unsigned(750731658,32),
    to_unsigned(750924552,32),
    to_unsigned(751117438,32),
    to_unsigned(751310318,32),
    to_unsigned(751503190,32),
    to_unsigned(751696056,32),
    to_unsigned(751888915,32),
    to_unsigned(752081766,32),
    to_unsigned(752274611,32),
    to_unsigned(752467449,32),
    to_unsigned(752660281,32),
    to_unsigned(752853105,32),
    to_unsigned(753045922,32),
    to_unsigned(753238732,32),
    to_unsigned(753431536,32),
    to_unsigned(753624332,32),
    to_unsigned(753817122,32),
    to_unsigned(754009904,32),
    to_unsigned(754202680,32),
    to_unsigned(754395449,32),
    to_unsigned(754588211,32),
    to_unsigned(754780966,32),
    to_unsigned(754973714,32),
    to_unsigned(755166455,32),
    to_unsigned(755359189,32),
    to_unsigned(755551916,32),
    to_unsigned(755744636,32),
    to_unsigned(755937350,32),
    to_unsigned(756130056,32),
    to_unsigned(756322755,32),
    to_unsigned(756515448,32),
    to_unsigned(756708133,32),
    to_unsigned(756900812,32),
    to_unsigned(757093483,32),
    to_unsigned(757286148,32),
    to_unsigned(757478805,32),
    to_unsigned(757671456,32),
    to_unsigned(757864100,32),
    to_unsigned(758056736,32),
    to_unsigned(758249366,32),
    to_unsigned(758441989,32),
    to_unsigned(758634605,32),
    to_unsigned(758827214,32),
    to_unsigned(759019816,32),
    to_unsigned(759212410,32),
    to_unsigned(759404998,32),
    to_unsigned(759597579,32),
    to_unsigned(759790153,32),
    to_unsigned(759982720,32),
    to_unsigned(760175280,32),
    to_unsigned(760367833,32),
    to_unsigned(760560379,32),
    to_unsigned(760752918,32),
    to_unsigned(760945450,32),
    to_unsigned(761137975,32),
    to_unsigned(761330493,32),
    to_unsigned(761523004,32),
    to_unsigned(761715508,32),
    to_unsigned(761908005,32),
    to_unsigned(762100495,32),
    to_unsigned(762292979,32),
    to_unsigned(762485455,32),
    to_unsigned(762677924,32),
    to_unsigned(762870386,32),
    to_unsigned(763062841,32),
    to_unsigned(763255289,32),
    to_unsigned(763447729,32),
    to_unsigned(763640163,32),
    to_unsigned(763832590,32),
    to_unsigned(764025010,32),
    to_unsigned(764217423,32),
    to_unsigned(764409829,32),
    to_unsigned(764602228,32),
    to_unsigned(764794620,32),
    to_unsigned(764987004,32),
    to_unsigned(765179382,32),
    to_unsigned(765371753,32),
    to_unsigned(765564117,32),
    to_unsigned(765756473,32),
    to_unsigned(765948823,32),
    to_unsigned(766141165,32),
    to_unsigned(766333501,32),
    to_unsigned(766525829,32),
    to_unsigned(766718151,32),
    to_unsigned(766910465,32),
    to_unsigned(767102772,32),
    to_unsigned(767295073,32),
    to_unsigned(767487366,32),
    to_unsigned(767679652,32),
    to_unsigned(767871931,32),
    to_unsigned(768064203,32),
    to_unsigned(768256468,32),
    to_unsigned(768448726,32),
    to_unsigned(768640977,32),
    to_unsigned(768833221,32),
    to_unsigned(769025458,32),
    to_unsigned(769217687,32),
    to_unsigned(769409910,32),
    to_unsigned(769602125,32),
    to_unsigned(769794334,32),
    to_unsigned(769986535,32),
    to_unsigned(770178730,32),
    to_unsigned(770370917,32),
    to_unsigned(770563097,32),
    to_unsigned(770755270,32),
    to_unsigned(770947436,32),
    to_unsigned(771139595,32),
    to_unsigned(771331747,32),
    to_unsigned(771523891,32),
    to_unsigned(771716029,32),
    to_unsigned(771908159,32),
    to_unsigned(772100283,32),
    to_unsigned(772292399,32),
    to_unsigned(772484508,32),
    to_unsigned(772676611,32),
    to_unsigned(772868706,32),
    to_unsigned(773060794,32),
    to_unsigned(773252874,32),
    to_unsigned(773444948,32),
    to_unsigned(773637015,32),
    to_unsigned(773829074,32),
    to_unsigned(774021127,32),
    to_unsigned(774213172,32),
    to_unsigned(774405210,32),
    to_unsigned(774597241,32),
    to_unsigned(774789265,32),
    to_unsigned(774981282,32),
    to_unsigned(775173291,32),
    to_unsigned(775365294,32),
    to_unsigned(775557289,32),
    to_unsigned(775749278,32),
    to_unsigned(775941259,32),
    to_unsigned(776133233,32),
    to_unsigned(776325200,32),
    to_unsigned(776517159,32),
    to_unsigned(776709112,32),
    to_unsigned(776901057,32),
    to_unsigned(777092996,32),
    to_unsigned(777284927,32),
    to_unsigned(777476851,32),
    to_unsigned(777668768,32),
    to_unsigned(777860678,32),
    to_unsigned(778052580,32),
    to_unsigned(778244476,32),
    to_unsigned(778436364,32),
    to_unsigned(778628245,32),
    to_unsigned(778820119,32),
    to_unsigned(779011986,32),
    to_unsigned(779203846,32),
    to_unsigned(779395698,32),
    to_unsigned(779587543,32),
    to_unsigned(779779382,32),
    to_unsigned(779971213,32),
    to_unsigned(780163036,32),
    to_unsigned(780354853,32),
    to_unsigned(780546663,32),
    to_unsigned(780738465,32),
    to_unsigned(780930260,32),
    to_unsigned(781122048,32),
    to_unsigned(781313829,32),
    to_unsigned(781505602,32),
    to_unsigned(781697369,32),
    to_unsigned(781889128,32),
    to_unsigned(782080880,32),
    to_unsigned(782272625,32),
    to_unsigned(782464363,32),
    to_unsigned(782656093,32),
    to_unsigned(782847816,32),
    to_unsigned(783039532,32),
    to_unsigned(783231241,32),
    to_unsigned(783422943,32),
    to_unsigned(783614637,32),
    to_unsigned(783806325,32),
    to_unsigned(783998005,32),
    to_unsigned(784189678,32),
    to_unsigned(784381343,32),
    to_unsigned(784573002,32),
    to_unsigned(784764653,32),
    to_unsigned(784956297,32),
    to_unsigned(785147934,32),
    to_unsigned(785339564,32),
    to_unsigned(785531186,32),
    to_unsigned(785722801,32),
    to_unsigned(785914409,32),
    to_unsigned(786106010,32),
    to_unsigned(786297603,32),
    to_unsigned(786489189,32),
    to_unsigned(786680768,32),
    to_unsigned(786872340,32),
    to_unsigned(787063905,32),
    to_unsigned(787255462,32),
    to_unsigned(787447012,32),
    to_unsigned(787638555,32),
    to_unsigned(787830091,32),
    to_unsigned(788021619,32),
    to_unsigned(788213140,32),
    to_unsigned(788404654,32),
    to_unsigned(788596161,32),
    to_unsigned(788787660,32),
    to_unsigned(788979152,32),
    to_unsigned(789170637,32),
    to_unsigned(789362115,32),
    to_unsigned(789553585,32),
    to_unsigned(789745048,32),
    to_unsigned(789936504,32),
    to_unsigned(790127953,32),
    to_unsigned(790319394,32),
    to_unsigned(790510828,32),
    to_unsigned(790702255,32),
    to_unsigned(790893675,32),
    to_unsigned(791085087,32),
    to_unsigned(791276492,32),
    to_unsigned(791467890,32),
    to_unsigned(791659280,32),
    to_unsigned(791850663,32),
    to_unsigned(792042039,32),
    to_unsigned(792233408,32),
    to_unsigned(792424769,32),
    to_unsigned(792616123,32),
    to_unsigned(792807470,32),
    to_unsigned(792998809,32),
    to_unsigned(793190141,32),
    to_unsigned(793381466,32),
    to_unsigned(793572784,32),
    to_unsigned(793764094,32),
    to_unsigned(793955397,32),
    to_unsigned(794146693,32),
    to_unsigned(794337981,32),
    to_unsigned(794529263,32),
    to_unsigned(794720536,32),
    to_unsigned(794911803,32),
    to_unsigned(795103062,32),
    to_unsigned(795294314,32),
    to_unsigned(795485559,32),
    to_unsigned(795676796,32),
    to_unsigned(795868026,32),
    to_unsigned(796059248,32),
    to_unsigned(796250464,32),
    to_unsigned(796441672,32),
    to_unsigned(796632872,32),
    to_unsigned(796824066,32),
    to_unsigned(797015252,32),
    to_unsigned(797206430,32),
    to_unsigned(797397602,32),
    to_unsigned(797588766,32),
    to_unsigned(797779923,32),
    to_unsigned(797971072,32),
    to_unsigned(798162214,32),
    to_unsigned(798353349,32),
    to_unsigned(798544476,32),
    to_unsigned(798735596,32),
    to_unsigned(798926709,32),
    to_unsigned(799117814,32),
    to_unsigned(799308912,32),
    to_unsigned(799500003,32),
    to_unsigned(799691086,32),
    to_unsigned(799882162,32),
    to_unsigned(800073231,32),
    to_unsigned(800264292,32),
    to_unsigned(800455346,32),
    to_unsigned(800646393,32),
    to_unsigned(800837432,32),
    to_unsigned(801028464,32),
    to_unsigned(801219488,32),
    to_unsigned(801410505,32),
    to_unsigned(801601515,32),
    to_unsigned(801792517,32),
    to_unsigned(801983512,32),
    to_unsigned(802174500,32),
    to_unsigned(802365480,32),
    to_unsigned(802556453,32),
    to_unsigned(802747418,32),
    to_unsigned(802938376,32),
    to_unsigned(803129327,32),
    to_unsigned(803320271,32),
    to_unsigned(803511207,32),
    to_unsigned(803702135,32),
    to_unsigned(803893056,32),
    to_unsigned(804083970,32),
    to_unsigned(804274877,32),
    to_unsigned(804465776,32),
    to_unsigned(804656667,32),
    to_unsigned(804847551,32),
    to_unsigned(805038428,32),
    to_unsigned(805229298,32),
    to_unsigned(805420160,32),
    to_unsigned(805611014,32),
    to_unsigned(805801862,32),
    to_unsigned(805992701,32),
    to_unsigned(806183534,32),
    to_unsigned(806374359,32),
    to_unsigned(806565176,32),
    to_unsigned(806755987,32),
    to_unsigned(806946789,32),
    to_unsigned(807137585,32),
    to_unsigned(807328373,32),
    to_unsigned(807519153,32),
    to_unsigned(807709926,32),
    to_unsigned(807900692,32),
    to_unsigned(808091450,32),
    to_unsigned(808282201,32),
    to_unsigned(808472944,32),
    to_unsigned(808663680,32),
    to_unsigned(808854409,32),
    to_unsigned(809045130,32),
    to_unsigned(809235843,32),
    to_unsigned(809426549,32),
    to_unsigned(809617248,32),
    to_unsigned(809807940,32),
    to_unsigned(809998623,32),
    to_unsigned(810189300,32),
    to_unsigned(810379969,32),
    to_unsigned(810570630,32),
    to_unsigned(810761284,32),
    to_unsigned(810951931,32),
    to_unsigned(811142570,32),
    to_unsigned(811333202,32),
    to_unsigned(811523826,32),
    to_unsigned(811714443,32),
    to_unsigned(811905052,32),
    to_unsigned(812095654,32),
    to_unsigned(812286249,32),
    to_unsigned(812476836,32),
    to_unsigned(812667415,32),
    to_unsigned(812857987,32),
    to_unsigned(813048552,32),
    to_unsigned(813239109,32),
    to_unsigned(813429658,32),
    to_unsigned(813620200,32),
    to_unsigned(813810735,32),
    to_unsigned(814001262,32),
    to_unsigned(814191782,32),
    to_unsigned(814382294,32),
    to_unsigned(814572799,32),
    to_unsigned(814763296,32),
    to_unsigned(814953786,32),
    to_unsigned(815144268,32),
    to_unsigned(815334743,32),
    to_unsigned(815525210,32),
    to_unsigned(815715670,32),
    to_unsigned(815906122,32),
    to_unsigned(816096567,32),
    to_unsigned(816287004,32),
    to_unsigned(816477434,32),
    to_unsigned(816667856,32),
    to_unsigned(816858270,32),
    to_unsigned(817048678,32),
    to_unsigned(817239077,32),
    to_unsigned(817429470,32),
    to_unsigned(817619854,32),
    to_unsigned(817810231,32),
    to_unsigned(818000601,32),
    to_unsigned(818190963,32),
    to_unsigned(818381318,32),
    to_unsigned(818571665,32),
    to_unsigned(818762005,32),
    to_unsigned(818952337,32),
    to_unsigned(819142661,32),
    to_unsigned(819332978,32),
    to_unsigned(819523288,32),
    to_unsigned(819713589,32),
    to_unsigned(819903884,32),
    to_unsigned(820094171,32),
    to_unsigned(820284450,32),
    to_unsigned(820474722,32),
    to_unsigned(820664986,32),
    to_unsigned(820855243,32),
    to_unsigned(821045492,32),
    to_unsigned(821235733,32),
    to_unsigned(821425968,32),
    to_unsigned(821616194,32),
    to_unsigned(821806413,32),
    to_unsigned(821996624,32),
    to_unsigned(822186828,32),
    to_unsigned(822377024,32),
    to_unsigned(822567213,32),
    to_unsigned(822757394,32),
    to_unsigned(822947568,32),
    to_unsigned(823137734,32),
    to_unsigned(823327892,32),
    to_unsigned(823518043,32),
    to_unsigned(823708187,32),
    to_unsigned(823898322,32),
    to_unsigned(824088451,32),
    to_unsigned(824278571,32),
    to_unsigned(824468684,32),
    to_unsigned(824658790,32),
    to_unsigned(824848888,32),
    to_unsigned(825038978,32),
    to_unsigned(825229061,32),
    to_unsigned(825419136,32),
    to_unsigned(825609203,32),
    to_unsigned(825799263,32),
    to_unsigned(825989316,32),
    to_unsigned(826179360,32),
    to_unsigned(826369398,32),
    to_unsigned(826559427,32),
    to_unsigned(826749449,32),
    to_unsigned(826939463,32),
    to_unsigned(827129470,32),
    to_unsigned(827319469,32),
    to_unsigned(827509461,32),
    to_unsigned(827699445,32),
    to_unsigned(827889421,32),
    to_unsigned(828079390,32),
    to_unsigned(828269351,32),
    to_unsigned(828459305,32),
    to_unsigned(828649251,32),
    to_unsigned(828839189,32),
    to_unsigned(829029120,32),
    to_unsigned(829219043,32),
    to_unsigned(829408958,32),
    to_unsigned(829598866,32),
    to_unsigned(829788766,32),
    to_unsigned(829978659,32),
    to_unsigned(830168543,32),
    to_unsigned(830358421,32),
    to_unsigned(830548290,32),
    to_unsigned(830738152,32),
    to_unsigned(830928007,32),
    to_unsigned(831117854,32),
    to_unsigned(831307693,32),
    to_unsigned(831497524,32),
    to_unsigned(831687348,32),
    to_unsigned(831877164,32),
    to_unsigned(832066973,32),
    to_unsigned(832256774,32),
    to_unsigned(832446567,32),
    to_unsigned(832636352,32),
    to_unsigned(832826130,32),
    to_unsigned(833015901,32),
    to_unsigned(833205663,32),
    to_unsigned(833395418,32),
    to_unsigned(833585166,32),
    to_unsigned(833774905,32),
    to_unsigned(833964637,32),
    to_unsigned(834154361,32),
    to_unsigned(834344078,32),
    to_unsigned(834533787,32),
    to_unsigned(834723488,32),
    to_unsigned(834913182,32),
    to_unsigned(835102868,32),
    to_unsigned(835292546,32),
    to_unsigned(835482217,32),
    to_unsigned(835671880,32),
    to_unsigned(835861535,32),
    to_unsigned(836051183,32),
    to_unsigned(836240822,32),
    to_unsigned(836430455,32),
    to_unsigned(836620079,32),
    to_unsigned(836809696,32),
    to_unsigned(836999305,32),
    to_unsigned(837188907,32),
    to_unsigned(837378500,32),
    to_unsigned(837568086,32),
    to_unsigned(837757665,32),
    to_unsigned(837947235,32),
    to_unsigned(838136798,32),
    to_unsigned(838326353,32),
    to_unsigned(838515901,32),
    to_unsigned(838705441,32),
    to_unsigned(838894973,32),
    to_unsigned(839084497,32),
    to_unsigned(839274014,32),
    to_unsigned(839463523,32),
    to_unsigned(839653024,32),
    to_unsigned(839842518,32),
    to_unsigned(840032003,32),
    to_unsigned(840221482,32),
    to_unsigned(840410952,32),
    to_unsigned(840600415,32),
    to_unsigned(840789869,32),
    to_unsigned(840979317,32),
    to_unsigned(841168756,32),
    to_unsigned(841358188,32),
    to_unsigned(841547612,32),
    to_unsigned(841737028,32),
    to_unsigned(841926437,32),
    to_unsigned(842115837,32),
    to_unsigned(842305230,32),
    to_unsigned(842494616,32),
    to_unsigned(842683993,32),
    to_unsigned(842873363,32),
    to_unsigned(843062725,32),
    to_unsigned(843252079,32),
    to_unsigned(843441426,32),
    to_unsigned(843630765,32),
    to_unsigned(843820096,32),
    to_unsigned(844009419,32),
    to_unsigned(844198735,32),
    to_unsigned(844388043,32),
    to_unsigned(844577343,32),
    to_unsigned(844766635,32),
    to_unsigned(844955919,32),
    to_unsigned(845145196,32),
    to_unsigned(845334465,32),
    to_unsigned(845523726,32),
    to_unsigned(845712980,32),
    to_unsigned(845902225,32),
    to_unsigned(846091463,32),
    to_unsigned(846280693,32),
    to_unsigned(846469915,32),
    to_unsigned(846659130,32),
    to_unsigned(846848337,32),
    to_unsigned(847037536,32),
    to_unsigned(847226727,32),
    to_unsigned(847415910,32),
    to_unsigned(847605086,32),
    to_unsigned(847794254,32),
    to_unsigned(847983414,32),
    to_unsigned(848172566,32),
    to_unsigned(848361710,32),
    to_unsigned(848550847,32),
    to_unsigned(848739976,32),
    to_unsigned(848929097,32),
    to_unsigned(849118210,32),
    to_unsigned(849307315,32),
    to_unsigned(849496413,32),
    to_unsigned(849685503,32),
    to_unsigned(849874585,32),
    to_unsigned(850063659,32),
    to_unsigned(850252725,32),
    to_unsigned(850441784,32),
    to_unsigned(850630835,32),
    to_unsigned(850819878,32),
    to_unsigned(851008913,32),
    to_unsigned(851197940,32),
    to_unsigned(851386959,32),
    to_unsigned(851575971,32),
    to_unsigned(851764975,32),
    to_unsigned(851953971,32),
    to_unsigned(852142959,32),
    to_unsigned(852331939,32),
    to_unsigned(852520912,32),
    to_unsigned(852709876,32),
    to_unsigned(852898833,32),
    to_unsigned(853087782,32),
    to_unsigned(853276723,32),
    to_unsigned(853465656,32),
    to_unsigned(853654582,32),
    to_unsigned(853843499,32),
    to_unsigned(854032409,32),
    to_unsigned(854221311,32),
    to_unsigned(854410205,32),
    to_unsigned(854599091,32),
    to_unsigned(854787970,32),
    to_unsigned(854976840,32),
    to_unsigned(855165703,32),
    to_unsigned(855354557,32),
    to_unsigned(855543404,32),
    to_unsigned(855732243,32),
    to_unsigned(855921074,32),
    to_unsigned(856109898,32),
    to_unsigned(856298713,32),
    to_unsigned(856487521,32),
    to_unsigned(856676320,32),
    to_unsigned(856865112,32),
    to_unsigned(857053896,32),
    to_unsigned(857242672,32),
    to_unsigned(857431440,32),
    to_unsigned(857620201,32),
    to_unsigned(857808953,32),
    to_unsigned(857997697,32),
    to_unsigned(858186434,32),
    to_unsigned(858375163,32),
    to_unsigned(858563884,32),
    to_unsigned(858752597,32),
    to_unsigned(858941302,32),
    to_unsigned(859129999,32),
    to_unsigned(859318688,32),
    to_unsigned(859507370,32),
    to_unsigned(859696043,32),
    to_unsigned(859884709,32),
    to_unsigned(860073366,32),
    to_unsigned(860262016,32),
    to_unsigned(860450658,32),
    to_unsigned(860639292,32),
    to_unsigned(860827918,32),
    to_unsigned(861016536,32),
    to_unsigned(861205146,32),
    to_unsigned(861393748,32),
    to_unsigned(861582343,32),
    to_unsigned(861770929,32),
    to_unsigned(861959508,32),
    to_unsigned(862148078,32),
    to_unsigned(862336641,32),
    to_unsigned(862525196,32),
    to_unsigned(862713743,32),
    to_unsigned(862902282,32),
    to_unsigned(863090813,32),
    to_unsigned(863279336,32),
    to_unsigned(863467851,32),
    to_unsigned(863656358,32),
    to_unsigned(863844857,32),
    to_unsigned(864033348,32),
    to_unsigned(864221832,32),
    to_unsigned(864410307,32),
    to_unsigned(864598775,32),
    to_unsigned(864787234,32),
    to_unsigned(864975686,32),
    to_unsigned(865164129,32),
    to_unsigned(865352565,32),
    to_unsigned(865540993,32),
    to_unsigned(865729412,32),
    to_unsigned(865917824,32),
    to_unsigned(866106228,32),
    to_unsigned(866294624,32),
    to_unsigned(866483012,32),
    to_unsigned(866671392,32),
    to_unsigned(866859764,32),
    to_unsigned(867048128,32),
    to_unsigned(867236484,32),
    to_unsigned(867424832,32),
    to_unsigned(867613172,32),
    to_unsigned(867801504,32),
    to_unsigned(867989828,32),
    to_unsigned(868178144,32),
    to_unsigned(868366452,32),
    to_unsigned(868554753,32),
    to_unsigned(868743045,32),
    to_unsigned(868931329,32),
    to_unsigned(869119605,32),
    to_unsigned(869307874,32),
    to_unsigned(869496134,32),
    to_unsigned(869684386,32),
    to_unsigned(869872630,32),
    to_unsigned(870060867,32),
    to_unsigned(870249095,32),
    to_unsigned(870437315,32),
    to_unsigned(870625527,32),
    to_unsigned(870813732,32),
    to_unsigned(871001928,32),
    to_unsigned(871190116,32),
    to_unsigned(871378297,32),
    to_unsigned(871566469,32),
    to_unsigned(871754633,32),
    to_unsigned(871942789,32),
    to_unsigned(872130938,32),
    to_unsigned(872319078,32),
    to_unsigned(872507210,32),
    to_unsigned(872695334,32),
    to_unsigned(872883450,32),
    to_unsigned(873071558,32),
    to_unsigned(873259658,32),
    to_unsigned(873447750,32),
    to_unsigned(873635834,32),
    to_unsigned(873823910,32),
    to_unsigned(874011978,32),
    to_unsigned(874200038,32),
    to_unsigned(874388090,32),
    to_unsigned(874576134,32),
    to_unsigned(874764170,32),
    to_unsigned(874952198,32),
    to_unsigned(875140218,32),
    to_unsigned(875328229,32),
    to_unsigned(875516233,32),
    to_unsigned(875704228,32),
    to_unsigned(875892216,32),
    to_unsigned(876080196,32),
    to_unsigned(876268167,32),
    to_unsigned(876456130,32),
    to_unsigned(876644086,32),
    to_unsigned(876832033,32),
    to_unsigned(877019972,32),
    to_unsigned(877207903,32),
    to_unsigned(877395827,32),
    to_unsigned(877583742,32),
    to_unsigned(877771649,32),
    to_unsigned(877959547,32),
    to_unsigned(878147438,32),
    to_unsigned(878335321,32),
    to_unsigned(878523196,32),
    to_unsigned(878711062,32),
    to_unsigned(878898921,32),
    to_unsigned(879086771,32),
    to_unsigned(879274614,32),
    to_unsigned(879462448,32),
    to_unsigned(879650274,32),
    to_unsigned(879838092,32),
    to_unsigned(880025902,32),
    to_unsigned(880213704,32),
    to_unsigned(880401498,32),
    to_unsigned(880589284,32),
    to_unsigned(880777062,32),
    to_unsigned(880964831,32),
    to_unsigned(881152593,32),
    to_unsigned(881340346,32),
    to_unsigned(881528091,32),
    to_unsigned(881715828,32),
    to_unsigned(881903558,32),
    to_unsigned(882091278,32),
    to_unsigned(882278991,32),
    to_unsigned(882466696,32),
    to_unsigned(882654393,32),
    to_unsigned(882842081,32),
    to_unsigned(883029762,32),
    to_unsigned(883217434,32),
    to_unsigned(883405098,32),
    to_unsigned(883592754,32),
    to_unsigned(883780402,32),
    to_unsigned(883968042,32),
    to_unsigned(884155674,32),
    to_unsigned(884343297,32),
    to_unsigned(884530913,32),
    to_unsigned(884718520,32),
    to_unsigned(884906119,32),
    to_unsigned(885093710,32),
    to_unsigned(885281293,32),
    to_unsigned(885468868,32),
    to_unsigned(885656434,32),
    to_unsigned(885843993,32),
    to_unsigned(886031543,32),
    to_unsigned(886219085,32),
    to_unsigned(886406619,32),
    to_unsigned(886594145,32),
    to_unsigned(886781663,32),
    to_unsigned(886969173,32),
    to_unsigned(887156674,32),
    to_unsigned(887344167,32),
    to_unsigned(887531652,32),
    to_unsigned(887719129,32),
    to_unsigned(887906598,32),
    to_unsigned(888094059,32),
    to_unsigned(888281511,32),
    to_unsigned(888468956,32),
    to_unsigned(888656392,32),
    to_unsigned(888843820,32),
    to_unsigned(889031240,32),
    to_unsigned(889218651,32),
    to_unsigned(889406055,32),
    to_unsigned(889593450,32),
    to_unsigned(889780837,32),
    to_unsigned(889968216,32),
    to_unsigned(890155587,32),
    to_unsigned(890342949,32),
    to_unsigned(890530304,32),
    to_unsigned(890717650,32),
    to_unsigned(890904988,32),
    to_unsigned(891092318,32),
    to_unsigned(891279640,32),
    to_unsigned(891466953,32),
    to_unsigned(891654258,32),
    to_unsigned(891841555,32),
    to_unsigned(892028844,32),
    to_unsigned(892216125,32),
    to_unsigned(892403397,32),
    to_unsigned(892590662,32),
    to_unsigned(892777918,32),
    to_unsigned(892965165,32),
    to_unsigned(893152405,32),
    to_unsigned(893339636,32),
    to_unsigned(893526860,32),
    to_unsigned(893714075,32),
    to_unsigned(893901282,32),
    to_unsigned(894088480,32),
    to_unsigned(894275670,32),
    to_unsigned(894462853,32),
    to_unsigned(894650026,32),
    to_unsigned(894837192,32),
    to_unsigned(895024350,32),
    to_unsigned(895211499,32),
    to_unsigned(895398640,32),
    to_unsigned(895585773,32),
    to_unsigned(895772897,32),
    to_unsigned(895960014,32),
    to_unsigned(896147122,32),
    to_unsigned(896334221,32),
    to_unsigned(896521313,32),
    to_unsigned(896708396,32),
    to_unsigned(896895472,32),
    to_unsigned(897082538,32),
    to_unsigned(897269597,32),
    to_unsigned(897456647,32),
    to_unsigned(897643690,32),
    to_unsigned(897830723,32),
    to_unsigned(898017749,32),
    to_unsigned(898204766,32),
    to_unsigned(898391776,32),
    to_unsigned(898578776,32),
    to_unsigned(898765769,32),
    to_unsigned(898952753,32),
    to_unsigned(899139729,32),
    to_unsigned(899326697,32),
    to_unsigned(899513657,32),
    to_unsigned(899700608,32),
    to_unsigned(899887551,32),
    to_unsigned(900074486,32),
    to_unsigned(900261412,32),
    to_unsigned(900448330,32),
    to_unsigned(900635240,32),
    to_unsigned(900822142,32),
    to_unsigned(901009035,32),
    to_unsigned(901195920,32),
    to_unsigned(901382797,32),
    to_unsigned(901569666,32),
    to_unsigned(901756526,32),
    to_unsigned(901943378,32),
    to_unsigned(902130222,32),
    to_unsigned(902317057,32),
    to_unsigned(902503884,32),
    to_unsigned(902690703,32),
    to_unsigned(902877513,32),
    to_unsigned(903064315,32),
    to_unsigned(903251109,32),
    to_unsigned(903437895,32),
    to_unsigned(903624672,32),
    to_unsigned(903811441,32),
    to_unsigned(903998202,32),
    to_unsigned(904184954,32),
    to_unsigned(904371698,32),
    to_unsigned(904558434,32),
    to_unsigned(904745161,32),
    to_unsigned(904931880,32),
    to_unsigned(905118591,32),
    to_unsigned(905305293,32),
    to_unsigned(905491987,32),
    to_unsigned(905678673,32),
    to_unsigned(905865351,32),
    to_unsigned(906052020,32),
    to_unsigned(906238681,32),
    to_unsigned(906425333,32),
    to_unsigned(906611977,32),
    to_unsigned(906798613,32),
    to_unsigned(906985241,32),
    to_unsigned(907171860,32),
    to_unsigned(907358470,32),
    to_unsigned(907545073,32),
    to_unsigned(907731667,32),
    to_unsigned(907918253,32),
    to_unsigned(908104830,32),
    to_unsigned(908291399,32),
    to_unsigned(908477960,32),
    to_unsigned(908664512,32),
    to_unsigned(908851057,32),
    to_unsigned(909037592,32),
    to_unsigned(909224120,32),
    to_unsigned(909410638,32),
    to_unsigned(909597149,32),
    to_unsigned(909783651,32),
    to_unsigned(909970145,32),
    to_unsigned(910156631,32),
    to_unsigned(910343108,32),
    to_unsigned(910529577,32),
    to_unsigned(910716037,32),
    to_unsigned(910902489,32),
    to_unsigned(911088933,32),
    to_unsigned(911275368,32),
    to_unsigned(911461795,32),
    to_unsigned(911648214,32),
    to_unsigned(911834624,32),
    to_unsigned(912021026,32),
    to_unsigned(912207419,32),
    to_unsigned(912393804,32),
    to_unsigned(912580181,32),
    to_unsigned(912766549,32),
    to_unsigned(912952909,32),
    to_unsigned(913139260,32),
    to_unsigned(913325603,32),
    to_unsigned(913511938,32),
    to_unsigned(913698264,32),
    to_unsigned(913884582,32),
    to_unsigned(914070892,32),
    to_unsigned(914257193,32),
    to_unsigned(914443485,32),
    to_unsigned(914629770,32),
    to_unsigned(914816045,32),
    to_unsigned(915002313,32),
    to_unsigned(915188572,32),
    to_unsigned(915374823,32),
    to_unsigned(915561065,32),
    to_unsigned(915747299,32),
    to_unsigned(915933524,32),
    to_unsigned(916119741,32),
    to_unsigned(916305949,32),
    to_unsigned(916492150,32),
    to_unsigned(916678341,32),
    to_unsigned(916864525,32),
    to_unsigned(917050699,32),
    to_unsigned(917236866,32),
    to_unsigned(917423024,32),
    to_unsigned(917609173,32),
    to_unsigned(917795314,32),
    to_unsigned(917981447,32),
    to_unsigned(918167571,32),
    to_unsigned(918353687,32),
    to_unsigned(918539794,32),
    to_unsigned(918725893,32),
    to_unsigned(918911984,32),
    to_unsigned(919098066,32),
    to_unsigned(919284139,32),
    to_unsigned(919470205,32),
    to_unsigned(919656261,32),
    to_unsigned(919842309,32),
    to_unsigned(920028349,32),
    to_unsigned(920214381,32),
    to_unsigned(920400403,32),
    to_unsigned(920586418,32),
    to_unsigned(920772424,32),
    to_unsigned(920958421,32),
    to_unsigned(921144410,32),
    to_unsigned(921330391,32),
    to_unsigned(921516363,32),
    to_unsigned(921702326,32),
    to_unsigned(921888282,32),
    to_unsigned(922074228,32),
    to_unsigned(922260166,32),
    to_unsigned(922446096,32),
    to_unsigned(922632017,32),
    to_unsigned(922817930,32),
    to_unsigned(923003834,32),
    to_unsigned(923189730,32),
    to_unsigned(923375617,32),
    to_unsigned(923561496,32),
    to_unsigned(923747366,32),
    to_unsigned(923933228,32),
    to_unsigned(924119082,32),
    to_unsigned(924304926,32),
    to_unsigned(924490763,32),
    to_unsigned(924676591,32),
    to_unsigned(924862410,32),
    to_unsigned(925048221,32),
    to_unsigned(925234023,32),
    to_unsigned(925419817,32),
    to_unsigned(925605602,32),
    to_unsigned(925791379,32),
    to_unsigned(925977147,32),
    to_unsigned(926162907,32),
    to_unsigned(926348658,32),
    to_unsigned(926534401,32),
    to_unsigned(926720135,32),
    to_unsigned(926905861,32),
    to_unsigned(927091578,32),
    to_unsigned(927277287,32),
    to_unsigned(927462987,32),
    to_unsigned(927648679,32),
    to_unsigned(927834362,32),
    to_unsigned(928020037,32),
    to_unsigned(928205703,32),
    to_unsigned(928391360,32),
    to_unsigned(928577009,32),
    to_unsigned(928762650,32),
    to_unsigned(928948281,32),
    to_unsigned(929133905,32),
    to_unsigned(929319520,32),
    to_unsigned(929505126,32),
    to_unsigned(929690724,32),
    to_unsigned(929876313,32),
    to_unsigned(930061894,32),
    to_unsigned(930247466,32),
    to_unsigned(930433029,32),
    to_unsigned(930618584,32),
    to_unsigned(930804131,32),
    to_unsigned(930989669,32),
    to_unsigned(931175198,32),
    to_unsigned(931360719,32),
    to_unsigned(931546231,32),
    to_unsigned(931731735,32),
    to_unsigned(931917230,32),
    to_unsigned(932102716,32),
    to_unsigned(932288194,32),
    to_unsigned(932473664,32),
    to_unsigned(932659124,32),
    to_unsigned(932844577,32),
    to_unsigned(933030020,32),
    to_unsigned(933215455,32),
    to_unsigned(933400882,32),
    to_unsigned(933586300,32),
    to_unsigned(933771709,32),
    to_unsigned(933957110,32),
    to_unsigned(934142502,32),
    to_unsigned(934327886,32),
    to_unsigned(934513261,32),
    to_unsigned(934698627,32),
    to_unsigned(934883985,32),
    to_unsigned(935069334,32),
    to_unsigned(935254675,32),
    to_unsigned(935440007,32),
    to_unsigned(935625330,32),
    to_unsigned(935810645,32),
    to_unsigned(935995952,32),
    to_unsigned(936181249,32),
    to_unsigned(936366538,32),
    to_unsigned(936551819,32),
    to_unsigned(936737091,32),
    to_unsigned(936922354,32),
    to_unsigned(937107608,32),
    to_unsigned(937292854,32),
    to_unsigned(937478092,32),
    to_unsigned(937663320,32),
    to_unsigned(937848541,32),
    to_unsigned(938033752,32),
    to_unsigned(938218955,32),
    to_unsigned(938404149,32),
    to_unsigned(938589335,32),
    to_unsigned(938774512,32),
    to_unsigned(938959680,32),
    to_unsigned(939144840,32),
    to_unsigned(939329991,32),
    to_unsigned(939515134,32),
    to_unsigned(939700268,32),
    to_unsigned(939885393,32),
    to_unsigned(940070509,32),
    to_unsigned(940255617,32),
    to_unsigned(940440717,32),
    to_unsigned(940625807,32),
    to_unsigned(940810889,32),
    to_unsigned(940995963,32),
    to_unsigned(941181027,32),
    to_unsigned(941366083,32),
    to_unsigned(941551131,32),
    to_unsigned(941736169,32),
    to_unsigned(941921200,32),
    to_unsigned(942106221,32),
    to_unsigned(942291234,32),
    to_unsigned(942476238,32),
    to_unsigned(942661233,32),
    to_unsigned(942846220,32),
    to_unsigned(943031198,32),
    to_unsigned(943216168,32),
    to_unsigned(943401128,32),
    to_unsigned(943586081,32),
    to_unsigned(943771024,32),
    to_unsigned(943955959,32),
    to_unsigned(944140885,32),
    to_unsigned(944325802,32),
    to_unsigned(944510711,32),
    to_unsigned(944695611,32),
    to_unsigned(944880502,32),
    to_unsigned(945065385,32),
    to_unsigned(945250259,32),
    to_unsigned(945435124,32),
    to_unsigned(945619981,32),
    to_unsigned(945804829,32),
    to_unsigned(945989668,32),
    to_unsigned(946174499,32),
    to_unsigned(946359320,32),
    to_unsigned(946544134,32),
    to_unsigned(946728938,32),
    to_unsigned(946913734,32),
    to_unsigned(947098521,32),
    to_unsigned(947283299,32),
    to_unsigned(947468069,32),
    to_unsigned(947652830,32),
    to_unsigned(947837582,32),
    to_unsigned(948022325,32),
    to_unsigned(948207060,32),
    to_unsigned(948391786,32),
    to_unsigned(948576503,32),
    to_unsigned(948761212,32),
    to_unsigned(948945912,32),
    to_unsigned(949130603,32),
    to_unsigned(949315286,32),
    to_unsigned(949499959,32),
    to_unsigned(949684624,32),
    to_unsigned(949869281,32),
    to_unsigned(950053928,32),
    to_unsigned(950238567,32),
    to_unsigned(950423197,32),
    to_unsigned(950607818,32),
    to_unsigned(950792431,32),
    to_unsigned(950977035,32),
    to_unsigned(951161630,32),
    to_unsigned(951346216,32),
    to_unsigned(951530794,32),
    to_unsigned(951715363,32),
    to_unsigned(951899923,32),
    to_unsigned(952084474,32),
    to_unsigned(952269017,32),
    to_unsigned(952453551,32),
    to_unsigned(952638076,32),
    to_unsigned(952822592,32),
    to_unsigned(953007100,32),
    to_unsigned(953191599,32),
    to_unsigned(953376089,32),
    to_unsigned(953560570,32),
    to_unsigned(953745043,32),
    to_unsigned(953929507,32),
    to_unsigned(954113962,32),
    to_unsigned(954298408,32),
    to_unsigned(954482845,32),
    to_unsigned(954667274,32),
    to_unsigned(954851694,32),
    to_unsigned(955036105,32),
    to_unsigned(955220507,32),
    to_unsigned(955404901,32),
    to_unsigned(955589286,32),
    to_unsigned(955773662,32),
    to_unsigned(955958029,32),
    to_unsigned(956142388,32),
    to_unsigned(956326737,32),
    to_unsigned(956511078,32),
    to_unsigned(956695410,32),
    to_unsigned(956879734,32),
    to_unsigned(957064048,32),
    to_unsigned(957248354,32),
    to_unsigned(957432651,32),
    to_unsigned(957616939,32),
    to_unsigned(957801218,32),
    to_unsigned(957985489,32),
    to_unsigned(958169750,32),
    to_unsigned(958354003,32),
    to_unsigned(958538247,32),
    to_unsigned(958722482,32),
    to_unsigned(958906709,32),
    to_unsigned(959090927,32),
    to_unsigned(959275135,32),
    to_unsigned(959459335,32),
    to_unsigned(959643527,32),
    to_unsigned(959827709,32),
    to_unsigned(960011883,32),
    to_unsigned(960196047,32),
    to_unsigned(960380203,32),
    to_unsigned(960564350,32),
    to_unsigned(960748488,32),
    to_unsigned(960932618,32),
    to_unsigned(961116738,32),
    to_unsigned(961300850,32),
    to_unsigned(961484953,32),
    to_unsigned(961669047,32),
    to_unsigned(961853132,32),
    to_unsigned(962037209,32),
    to_unsigned(962221276,32),
    to_unsigned(962405335,32),
    to_unsigned(962589385,32),
    to_unsigned(962773426,32),
    to_unsigned(962957458,32),
    to_unsigned(963141481,32),
    to_unsigned(963325496,32),
    to_unsigned(963509501,32),
    to_unsigned(963693498,32),
    to_unsigned(963877486,32),
    to_unsigned(964061465,32),
    to_unsigned(964245435,32),
    to_unsigned(964429396,32),
    to_unsigned(964613349,32),
    to_unsigned(964797292,32),
    to_unsigned(964981227,32),
    to_unsigned(965165153,32),
    to_unsigned(965349070,32),
    to_unsigned(965532978,32),
    to_unsigned(965716877,32),
    to_unsigned(965900767,32),
    to_unsigned(966084649,32),
    to_unsigned(966268521,32),
    to_unsigned(966452385,32),
    to_unsigned(966636240,32),
    to_unsigned(966820086,32),
    to_unsigned(967003923,32),
    to_unsigned(967187751,32),
    to_unsigned(967371570,32),
    to_unsigned(967555381,32),
    to_unsigned(967739182,32),
    to_unsigned(967922975,32),
    to_unsigned(968106758,32),
    to_unsigned(968290533,32),
    to_unsigned(968474299,32),
    to_unsigned(968658056,32),
    to_unsigned(968841804,32),
    to_unsigned(969025543,32),
    to_unsigned(969209274,32),
    to_unsigned(969392995,32),
    to_unsigned(969576707,32),
    to_unsigned(969760411,32),
    to_unsigned(969944105,32),
    to_unsigned(970127791,32),
    to_unsigned(970311468,32),
    to_unsigned(970495136,32),
    to_unsigned(970678795,32),
    to_unsigned(970862445,32),
    to_unsigned(971046086,32),
    to_unsigned(971229718,32),
    to_unsigned(971413341,32),
    to_unsigned(971596956,32),
    to_unsigned(971780561,32),
    to_unsigned(971964157,32),
    to_unsigned(972147745,32),
    to_unsigned(972331324,32),
    to_unsigned(972514893,32),
    to_unsigned(972698454,32),
    to_unsigned(972882006,32),
    to_unsigned(973065548,32),
    to_unsigned(973249082,32),
    to_unsigned(973432607,32),
    to_unsigned(973616123,32),
    to_unsigned(973799630,32),
    to_unsigned(973983128,32),
    to_unsigned(974166618,32),
    to_unsigned(974350098,32),
    to_unsigned(974533569,32),
    to_unsigned(974717031,32),
    to_unsigned(974900484,32),
    to_unsigned(975083929,32),
    to_unsigned(975267364,32),
    to_unsigned(975450791,32),
    to_unsigned(975634208,32),
    to_unsigned(975817617,32),
    to_unsigned(976001016,32),
    to_unsigned(976184407,32),
    to_unsigned(976367788,32),
    to_unsigned(976551161,32),
    to_unsigned(976734524,32),
    to_unsigned(976917879,32),
    to_unsigned(977101225,32),
    to_unsigned(977284561,32),
    to_unsigned(977467889,32),
    to_unsigned(977651208,32),
    to_unsigned(977834518,32),
    to_unsigned(978017818,32),
    to_unsigned(978201110,32),
    to_unsigned(978384393,32),
    to_unsigned(978567666,32),
    to_unsigned(978750931,32),
    to_unsigned(978934187,32),
    to_unsigned(979117434,32),
    to_unsigned(979300672,32),
    to_unsigned(979483900,32),
    to_unsigned(979667120,32),
    to_unsigned(979850331,32),
    to_unsigned(980033533,32),
    to_unsigned(980216725,32),
    to_unsigned(980399909,32),
    to_unsigned(980583084,32),
    to_unsigned(980766250,32),
    to_unsigned(980949406,32),
    to_unsigned(981132554,32),
    to_unsigned(981315693,32),
    to_unsigned(981498822,32),
    to_unsigned(981681943,32),
    to_unsigned(981865054,32),
    to_unsigned(982048157,32),
    to_unsigned(982231251,32),
    to_unsigned(982414335,32),
    to_unsigned(982597411,32),
    to_unsigned(982780477,32),
    to_unsigned(982963534,32),
    to_unsigned(983146583,32),
    to_unsigned(983329622,32),
    to_unsigned(983512653,32),
    to_unsigned(983695674,32),
    to_unsigned(983878686,32),
    to_unsigned(984061689,32),
    to_unsigned(984244683,32),
    to_unsigned(984427668,32),
    to_unsigned(984610644,32),
    to_unsigned(984793611,32),
    to_unsigned(984976569,32),
    to_unsigned(985159518,32),
    to_unsigned(985342458,32),
    to_unsigned(985525389,32),
    to_unsigned(985708311,32),
    to_unsigned(985891223,32),
    to_unsigned(986074127,32),
    to_unsigned(986257021,32),
    to_unsigned(986439907,32),
    to_unsigned(986622783,32),
    to_unsigned(986805651,32),
    to_unsigned(986988509,32),
    to_unsigned(987171358,32),
    to_unsigned(987354198,32),
    to_unsigned(987537029,32),
    to_unsigned(987719851,32),
    to_unsigned(987902664,32),
    to_unsigned(988085468,32),
    to_unsigned(988268263,32),
    to_unsigned(988451048,32),
    to_unsigned(988633825,32),
    to_unsigned(988816592,32),
    to_unsigned(988999351,32),
    to_unsigned(989182100,32),
    to_unsigned(989364840,32),
    to_unsigned(989547571,32),
    to_unsigned(989730293,32),
    to_unsigned(989913006,32),
    to_unsigned(990095710,32),
    to_unsigned(990278405,32),
    to_unsigned(990461090,32),
    to_unsigned(990643767,32),
    to_unsigned(990826434,32),
    to_unsigned(991009092,32),
    to_unsigned(991191742,32),
    to_unsigned(991374382,32),
    to_unsigned(991557013,32),
    to_unsigned(991739634,32),
    to_unsigned(991922247,32),
    to_unsigned(992104851,32),
    to_unsigned(992287445,32),
    to_unsigned(992470031,32),
    to_unsigned(992652607,32),
    to_unsigned(992835174,32),
    to_unsigned(993017732,32),
    to_unsigned(993200281,32),
    to_unsigned(993382820,32),
    to_unsigned(993565351,32),
    to_unsigned(993747873,32),
    to_unsigned(993930385,32),
    to_unsigned(994112888,32),
    to_unsigned(994295382,32),
    to_unsigned(994477867,32),
    to_unsigned(994660343,32),
    to_unsigned(994842809,32),
    to_unsigned(995025267,32),
    to_unsigned(995207715,32),
    to_unsigned(995390155,32),
    to_unsigned(995572585,32),
    to_unsigned(995755005,32),
    to_unsigned(995937417,32),
    to_unsigned(996119820,32),
    to_unsigned(996302213,32),
    to_unsigned(996484598,32),
    to_unsigned(996666973,32),
    to_unsigned(996849339,32),
    to_unsigned(997031695,32),
    to_unsigned(997214043,32),
    to_unsigned(997396382,32),
    to_unsigned(997578711,32),
    to_unsigned(997761031,32),
    to_unsigned(997943342,32),
    to_unsigned(998125644,32),
    to_unsigned(998307936,32),
    to_unsigned(998490220,32),
    to_unsigned(998672494,32),
    to_unsigned(998854759,32),
    to_unsigned(999037015,32),
    to_unsigned(999219262,32),
    to_unsigned(999401499,32),
    to_unsigned(999583728,32),
    to_unsigned(999765947,32),
    to_unsigned(999948157,32),
    to_unsigned(1000130357,32),
    to_unsigned(1000312549,32),
    to_unsigned(1000494731,32),
    to_unsigned(1000676905,32),
    to_unsigned(1000859069,32),
    to_unsigned(1001041223,32),
    to_unsigned(1001223369,32),
    to_unsigned(1001405505,32),
    to_unsigned(1001587632,32),
    to_unsigned(1001769750,32),
    to_unsigned(1001951859,32),
    to_unsigned(1002133959,32),
    to_unsigned(1002316049,32),
    to_unsigned(1002498130,32),
    to_unsigned(1002680202,32),
    to_unsigned(1002862265,32),
    to_unsigned(1003044318,32),
    to_unsigned(1003226363,32),
    to_unsigned(1003408398,32),
    to_unsigned(1003590423,32),
    to_unsigned(1003772440,32),
    to_unsigned(1003954447,32),
    to_unsigned(1004136446,32),
    to_unsigned(1004318434,32),
    to_unsigned(1004500414,32),
    to_unsigned(1004682385,32),
    to_unsigned(1004864346,32),
    to_unsigned(1005046298,32),
    to_unsigned(1005228241,32),
    to_unsigned(1005410174,32),
    to_unsigned(1005592098,32),
    to_unsigned(1005774013,32),
    to_unsigned(1005955919,32),
    to_unsigned(1006137816,32),
    to_unsigned(1006319703,32),
    to_unsigned(1006501581,32),
    to_unsigned(1006683450,32),
    to_unsigned(1006865309,32),
    to_unsigned(1007047159,32),
    to_unsigned(1007229000,32),
    to_unsigned(1007410832,32),
    to_unsigned(1007592655,32),
    to_unsigned(1007774468,32),
    to_unsigned(1007956272,32),
    to_unsigned(1008138067,32),
    to_unsigned(1008319852,32),
    to_unsigned(1008501628,32),
    to_unsigned(1008683395,32),
    to_unsigned(1008865153,32),
    to_unsigned(1009046901,32),
    to_unsigned(1009228640,32),
    to_unsigned(1009410370,32),
    to_unsigned(1009592090,32),
    to_unsigned(1009773802,32),
    to_unsigned(1009955504,32),
    to_unsigned(1010137196,32),
    to_unsigned(1010318880,32),
    to_unsigned(1010500554,32),
    to_unsigned(1010682219,32),
    to_unsigned(1010863874,32),
    to_unsigned(1011045520,32),
    to_unsigned(1011227157,32),
    to_unsigned(1011408785,32),
    to_unsigned(1011590403,32),
    to_unsigned(1011772012,32),
    to_unsigned(1011953612,32),
    to_unsigned(1012135202,32),
    to_unsigned(1012316784,32),
    to_unsigned(1012498355,32),
    to_unsigned(1012679918,32),
    to_unsigned(1012861471,32),
    to_unsigned(1013043015,32),
    to_unsigned(1013224550,32),
    to_unsigned(1013406075,32),
    to_unsigned(1013587591,32),
    to_unsigned(1013769098,32),
    to_unsigned(1013950595,32),
    to_unsigned(1014132083,32),
    to_unsigned(1014313562,32),
    to_unsigned(1014495031,32),
    to_unsigned(1014676491,32),
    to_unsigned(1014857942,32),
    to_unsigned(1015039383,32),
    to_unsigned(1015220815,32),
    to_unsigned(1015402238,32),
    to_unsigned(1015583651,32),
    to_unsigned(1015765055,32),
    to_unsigned(1015946450,32),
    to_unsigned(1016127836,32),
    to_unsigned(1016309212,32),
    to_unsigned(1016490578,32),
    to_unsigned(1016671936,32),
    to_unsigned(1016853284,32),
    to_unsigned(1017034622,32),
    to_unsigned(1017215952,32),
    to_unsigned(1017397272,32),
    to_unsigned(1017578582,32),
    to_unsigned(1017759884,32),
    to_unsigned(1017941175,32),
    to_unsigned(1018122458,32),
    to_unsigned(1018303731,32),
    to_unsigned(1018484995,32),
    to_unsigned(1018666250,32),
    to_unsigned(1018847495,32),
    to_unsigned(1019028730,32),
    to_unsigned(1019209957,32),
    to_unsigned(1019391174,32),
    to_unsigned(1019572381,32),
    to_unsigned(1019753580,32),
    to_unsigned(1019934769,32),
    to_unsigned(1020115948,32),
    to_unsigned(1020297118,32),
    to_unsigned(1020478279,32),
    to_unsigned(1020659430,32),
    to_unsigned(1020840572,32),
    to_unsigned(1021021705,32),
    to_unsigned(1021202828,32),
    to_unsigned(1021383942,32),
    to_unsigned(1021565047,32),
    to_unsigned(1021746142,32),
    to_unsigned(1021927227,32),
    to_unsigned(1022108304,32),
    to_unsigned(1022289370,32),
    to_unsigned(1022470428,32),
    to_unsigned(1022651476,32),
    to_unsigned(1022832515,32),
    to_unsigned(1023013544,32),
    to_unsigned(1023194564,32),
    to_unsigned(1023375574,32),
    to_unsigned(1023556576,32),
    to_unsigned(1023737567,32),
    to_unsigned(1023918549,32),
    to_unsigned(1024099522,32),
    to_unsigned(1024280486,32),
    to_unsigned(1024461440,32),
    to_unsigned(1024642384,32),
    to_unsigned(1024823320,32),
    to_unsigned(1025004245,32),
    to_unsigned(1025185162,32),
    to_unsigned(1025366069,32),
    to_unsigned(1025546966,32),
    to_unsigned(1025727854,32),
    to_unsigned(1025908733,32),
    to_unsigned(1026089602,32),
    to_unsigned(1026270462,32),
    to_unsigned(1026451312,32),
    to_unsigned(1026632153,32),
    to_unsigned(1026812985,32),
    to_unsigned(1026993807,32),
    to_unsigned(1027174619,32),
    to_unsigned(1027355422,32),
    to_unsigned(1027536216,32),
    to_unsigned(1027717000,32),
    to_unsigned(1027897775,32),
    to_unsigned(1028078540,32),
    to_unsigned(1028259296,32),
    to_unsigned(1028440043,32),
    to_unsigned(1028620780,32),
    to_unsigned(1028801507,32),
    to_unsigned(1028982226,32),
    to_unsigned(1029162934,32),
    to_unsigned(1029343633,32),
    to_unsigned(1029524323,32),
    to_unsigned(1029705003,32),
    to_unsigned(1029885674,32),
    to_unsigned(1030066336,32),
    to_unsigned(1030246987,32),
    to_unsigned(1030427630,32),
    to_unsigned(1030608263,32),
    to_unsigned(1030788886,32),
    to_unsigned(1030969500,32),
    to_unsigned(1031150105,32),
    to_unsigned(1031330700,32),
    to_unsigned(1031511285,32),
    to_unsigned(1031691861,32),
    to_unsigned(1031872428,32),
    to_unsigned(1032052985,32),
    to_unsigned(1032233533,32),
    to_unsigned(1032414071,32),
    to_unsigned(1032594599,32),
    to_unsigned(1032775118,32),
    to_unsigned(1032955628,32),
    to_unsigned(1033136128,32),
    to_unsigned(1033316619,32),
    to_unsigned(1033497100,32),
    to_unsigned(1033677572,32),
    to_unsigned(1033858034,32),
    to_unsigned(1034038486,32),
    to_unsigned(1034218930,32),
    to_unsigned(1034399363,32),
    to_unsigned(1034579787,32),
    to_unsigned(1034760202,32),
    to_unsigned(1034940607,32),
    to_unsigned(1035121003,32),
    to_unsigned(1035301389,32),
    to_unsigned(1035481765,32),
    to_unsigned(1035662132,32),
    to_unsigned(1035842490,32),
    to_unsigned(1036022838,32),
    to_unsigned(1036203176,32),
    to_unsigned(1036383505,32),
    to_unsigned(1036563825,32),
    to_unsigned(1036744135,32),
    to_unsigned(1036924435,32),
    to_unsigned(1037104726,32),
    to_unsigned(1037285007,32),
    to_unsigned(1037465279,32),
    to_unsigned(1037645541,32),
    to_unsigned(1037825794,32),
    to_unsigned(1038006037,32),
    to_unsigned(1038186271,32),
    to_unsigned(1038366495,32),
    to_unsigned(1038546709,32),
    to_unsigned(1038726914,32),
    to_unsigned(1038907110,32),
    to_unsigned(1039087296,32),
    to_unsigned(1039267472,32),
    to_unsigned(1039447639,32),
    to_unsigned(1039627796,32),
    to_unsigned(1039807944,32),
    to_unsigned(1039988082,32),
    to_unsigned(1040168210,32),
    to_unsigned(1040348329,32),
    to_unsigned(1040528439,32),
    to_unsigned(1040708539,32),
    to_unsigned(1040888629,32),
    to_unsigned(1041068710,32),
    to_unsigned(1041248781,32),
    to_unsigned(1041428843,32),
    to_unsigned(1041608895,32),
    to_unsigned(1041788937,32),
    to_unsigned(1041968970,32),
    to_unsigned(1042148993,32),
    to_unsigned(1042329007,32),
    to_unsigned(1042509011,32),
    to_unsigned(1042689006,32),
    to_unsigned(1042868991,32),
    to_unsigned(1043048966,32),
    to_unsigned(1043228932,32),
    to_unsigned(1043408888,32),
    to_unsigned(1043588835,32),
    to_unsigned(1043768772,32),
    to_unsigned(1043948699,32),
    to_unsigned(1044128617,32),
    to_unsigned(1044308525,32),
    to_unsigned(1044488424,32),
    to_unsigned(1044668313,32),
    to_unsigned(1044848192,32),
    to_unsigned(1045028062,32),
    to_unsigned(1045207922,32),
    to_unsigned(1045387773,32),
    to_unsigned(1045567614,32),
    to_unsigned(1045747445,32),
    to_unsigned(1045927267,32),
    to_unsigned(1046107079,32),
    to_unsigned(1046286882,32),
    to_unsigned(1046466675,32),
    to_unsigned(1046646458,32),
    to_unsigned(1046826232,32),
    to_unsigned(1047005996,32),
    to_unsigned(1047185750,32),
    to_unsigned(1047365495,32),
    to_unsigned(1047545231,32),
    to_unsigned(1047724956,32),
    to_unsigned(1047904672,32),
    to_unsigned(1048084378,32),
    to_unsigned(1048264075,32),
    to_unsigned(1048443762,32),
    to_unsigned(1048623439,32),
    to_unsigned(1048803107,32),
    to_unsigned(1048982765,32),
    to_unsigned(1049162414,32),
    to_unsigned(1049342053,32),
    to_unsigned(1049521682,32),
    to_unsigned(1049701301,32),
    to_unsigned(1049880911,32),
    to_unsigned(1050060512,32),
    to_unsigned(1050240102,32),
    to_unsigned(1050419683,32),
    to_unsigned(1050599254,32),
    to_unsigned(1050778816,32),
    to_unsigned(1050958368,32),
    to_unsigned(1051137910,32),
    to_unsigned(1051317443,32),
    to_unsigned(1051496966,32),
    to_unsigned(1051676479,32),
    to_unsigned(1051855983,32),
    to_unsigned(1052035477,32),
    to_unsigned(1052214961,32),
    to_unsigned(1052394436,32),
    to_unsigned(1052573901,32),
    to_unsigned(1052753356,32),
    to_unsigned(1052932802,32),
    to_unsigned(1053112238,32),
    to_unsigned(1053291664,32),
    to_unsigned(1053471081,32),
    to_unsigned(1053650487,32),
    to_unsigned(1053829885,32),
    to_unsigned(1054009272,32),
    to_unsigned(1054188650,32),
    to_unsigned(1054368018,32),
    to_unsigned(1054547377,32),
    to_unsigned(1054726725,32),
    to_unsigned(1054906065,32),
    to_unsigned(1055085394,32),
    to_unsigned(1055264714,32),
    to_unsigned(1055444024,32),
    to_unsigned(1055623324,32),
    to_unsigned(1055802614,32),
    to_unsigned(1055981895,32),
    to_unsigned(1056161166,32),
    to_unsigned(1056340428,32),
    to_unsigned(1056519680,32),
    to_unsigned(1056698922,32),
    to_unsigned(1056878154,32),
    to_unsigned(1057057377,32),
    to_unsigned(1057236589,32),
    to_unsigned(1057415793,32),
    to_unsigned(1057594986,32),
    to_unsigned(1057774170,32),
    to_unsigned(1057953344,32),
    to_unsigned(1058132508,32),
    to_unsigned(1058311663,32),
    to_unsigned(1058490807,32),
    to_unsigned(1058669943,32),
    to_unsigned(1058849068,32),
    to_unsigned(1059028184,32),
    to_unsigned(1059207289,32),
    to_unsigned(1059386386,32),
    to_unsigned(1059565472,32),
    to_unsigned(1059744549,32),
    to_unsigned(1059923616,32),
    to_unsigned(1060102673,32),
    to_unsigned(1060281720,32),
    to_unsigned(1060460758,32),
    to_unsigned(1060639786,32),
    to_unsigned(1060818804,32),
    to_unsigned(1060997813,32),
    to_unsigned(1061176811,32),
    to_unsigned(1061355800,32),
    to_unsigned(1061534780,32),
    to_unsigned(1061713749,32),
    to_unsigned(1061892709,32),
    to_unsigned(1062071659,32),
    to_unsigned(1062250599,32),
    to_unsigned(1062429529,32),
    to_unsigned(1062608450,32),
    to_unsigned(1062787361,32),
    to_unsigned(1062966262,32),
    to_unsigned(1063145153,32),
    to_unsigned(1063324035,32),
    to_unsigned(1063502906,32),
    to_unsigned(1063681768,32),
    to_unsigned(1063860621,32),
    to_unsigned(1064039463,32),
    to_unsigned(1064218296,32),
    to_unsigned(1064397119,32),
    to_unsigned(1064575932,32),
    to_unsigned(1064754735,32),
    to_unsigned(1064933529,32),
    to_unsigned(1065112312,32),
    to_unsigned(1065291086,32),
    to_unsigned(1065469850,32),
    to_unsigned(1065648605,32),
    to_unsigned(1065827349,32),
    to_unsigned(1066006084,32),
    to_unsigned(1066184809,32),
    to_unsigned(1066363524,32),
    to_unsigned(1066542230,32),
    to_unsigned(1066720925,32),
    to_unsigned(1066899611,32),
    to_unsigned(1067078287,32),
    to_unsigned(1067256953,32),
    to_unsigned(1067435610,32),
    to_unsigned(1067614256,32),
    to_unsigned(1067792893,32),
    to_unsigned(1067971520,32),
    to_unsigned(1068150137,32),
    to_unsigned(1068328744,32),
    to_unsigned(1068507341,32),
    to_unsigned(1068685929,32),
    to_unsigned(1068864507,32),
    to_unsigned(1069043075,32),
    to_unsigned(1069221633,32),
    to_unsigned(1069400181,32),
    to_unsigned(1069578720,32),
    to_unsigned(1069757248,32),
    to_unsigned(1069935767,32),
    to_unsigned(1070114276,32),
    to_unsigned(1070292775,32),
    to_unsigned(1070471265,32),
    to_unsigned(1070649744,32),
    to_unsigned(1070828214,32),
    to_unsigned(1071006674,32),
    to_unsigned(1071185124,32),
    to_unsigned(1071363564,32),
    to_unsigned(1071541994,32),
    to_unsigned(1071720414,32),
    to_unsigned(1071898825,32),
    to_unsigned(1072077226,32),
    to_unsigned(1072255617,32),
    to_unsigned(1072433998,32),
    to_unsigned(1072612369,32),
    to_unsigned(1072790730,32),
    to_unsigned(1072969081,32),
    to_unsigned(1073147423,32),
    to_unsigned(1073325755,32),
    to_unsigned(1073504076,32),
    to_unsigned(1073682388,32),
    to_unsigned(1073860690,32),
    to_unsigned(1074038983,32),
    to_unsigned(1074217265,32),
    to_unsigned(1074395537,32),
    to_unsigned(1074573800,32),
    to_unsigned(1074752053,32),
    to_unsigned(1074930296,32),
    to_unsigned(1075108529,32),
    to_unsigned(1075286752,32),
    to_unsigned(1075464965,32),
    to_unsigned(1075643168,32),
    to_unsigned(1075821362,32),
    to_unsigned(1075999545,32),
    to_unsigned(1076177719,32),
    to_unsigned(1076355883,32),
    to_unsigned(1076534036,32),
    to_unsigned(1076712180,32),
    to_unsigned(1076890314,32),
    to_unsigned(1077068439,32),
    to_unsigned(1077246553,32),
    to_unsigned(1077424657,32),
    to_unsigned(1077602752,32),
    to_unsigned(1077780836,32),
    to_unsigned(1077958911,32),
    to_unsigned(1078136976,32),
    to_unsigned(1078315030,32),
    to_unsigned(1078493075,32),
    to_unsigned(1078671110,32),
    to_unsigned(1078849135,32),
    to_unsigned(1079027151,32),
    to_unsigned(1079205156,32),
    to_unsigned(1079383151,32),
    to_unsigned(1079561137,32),
    to_unsigned(1079739112,32),
    to_unsigned(1079917078,32),
    to_unsigned(1080095033,32),
    to_unsigned(1080272979,32),
    to_unsigned(1080450915,32),
    to_unsigned(1080628841,32),
    to_unsigned(1080806757,32),
    to_unsigned(1080984663,32),
    to_unsigned(1081162559,32),
    to_unsigned(1081340445,32),
    to_unsigned(1081518321,32),
    to_unsigned(1081696187,32),
    to_unsigned(1081874043,32),
    to_unsigned(1082051890,32),
    to_unsigned(1082229726,32),
    to_unsigned(1082407553,32),
    to_unsigned(1082585369,32),
    to_unsigned(1082763176,32),
    to_unsigned(1082940972,32),
    to_unsigned(1083118759,32),
    to_unsigned(1083296536,32),
    to_unsigned(1083474302,32),
    to_unsigned(1083652059,32),
    to_unsigned(1083829806,32),
    to_unsigned(1084007543,32),
    to_unsigned(1084185270,32),
    to_unsigned(1084362986,32),
    to_unsigned(1084540693,32),
    to_unsigned(1084718390,32),
    to_unsigned(1084896077,32),
    to_unsigned(1085073754,32),
    to_unsigned(1085251421,32),
    to_unsigned(1085429079,32),
    to_unsigned(1085606726,32),
    to_unsigned(1085784363,32),
    to_unsigned(1085961990,32),
    to_unsigned(1086139607,32),
    to_unsigned(1086317214,32),
    to_unsigned(1086494812,32),
    to_unsigned(1086672399,32),
    to_unsigned(1086849976,32),
    to_unsigned(1087027543,32),
    to_unsigned(1087205100,32),
    to_unsigned(1087382648,32),
    to_unsigned(1087560185,32),
    to_unsigned(1087737712,32),
    to_unsigned(1087915229,32),
    to_unsigned(1088092737,32),
    to_unsigned(1088270234,32),
    to_unsigned(1088447721,32),
    to_unsigned(1088625199,32),
    to_unsigned(1088802666,32),
    to_unsigned(1088980123,32),
    to_unsigned(1089157570,32),
    to_unsigned(1089335007,32),
    to_unsigned(1089512435,32),
    to_unsigned(1089689852,32),
    to_unsigned(1089867259,32),
    to_unsigned(1090044656,32),
    to_unsigned(1090222043,32),
    to_unsigned(1090399420,32),
    to_unsigned(1090576787,32),
    to_unsigned(1090754145,32),
    to_unsigned(1090931492,32),
    to_unsigned(1091108829,32),
    to_unsigned(1091286156,32),
    to_unsigned(1091463473,32),
    to_unsigned(1091640779,32),
    to_unsigned(1091818076,32),
    to_unsigned(1091995363,32),
    to_unsigned(1092172640,32),
    to_unsigned(1092349907,32),
    to_unsigned(1092527164,32),
    to_unsigned(1092704410,32),
    to_unsigned(1092881647,32),
    to_unsigned(1093058873,32),
    to_unsigned(1093236090,32),
    to_unsigned(1093413297,32),
    to_unsigned(1093590493,32),
    to_unsigned(1093767679,32),
    to_unsigned(1093944856,32),
    to_unsigned(1094122022,32),
    to_unsigned(1094299178,32),
    to_unsigned(1094476324,32),
    to_unsigned(1094653461,32),
    to_unsigned(1094830587,32),
    to_unsigned(1095007703,32),
    to_unsigned(1095184809,32),
    to_unsigned(1095361904,32),
    to_unsigned(1095538990,32),
    to_unsigned(1095716066,32),
    to_unsigned(1095893132,32),
    to_unsigned(1096070187,32),
    to_unsigned(1096247233,32),
    to_unsigned(1096424268,32),
    to_unsigned(1096601293,32),
    to_unsigned(1096778309,32),
    to_unsigned(1096955314,32),
    to_unsigned(1097132309,32),
    to_unsigned(1097309294,32),
    to_unsigned(1097486269,32),
    to_unsigned(1097663234,32),
    to_unsigned(1097840189,32),
    to_unsigned(1098017133,32),
    to_unsigned(1098194068,32),
    to_unsigned(1098370992,32),
    to_unsigned(1098547907,32),
    to_unsigned(1098724811,32),
    to_unsigned(1098901705,32),
    to_unsigned(1099078589,32),
    to_unsigned(1099255463,32),
    to_unsigned(1099432327,32),
    to_unsigned(1099609181,32),
    to_unsigned(1099786025,32),
    to_unsigned(1099962858,32),
    to_unsigned(1100139682,32),
    to_unsigned(1100316495,32),
    to_unsigned(1100493298,32),
    to_unsigned(1100670091,32),
    to_unsigned(1100846874,32),
    to_unsigned(1101023647,32),
    to_unsigned(1101200410,32),
    to_unsigned(1101377162,32),
    to_unsigned(1101553905,32),
    to_unsigned(1101730637,32),
    to_unsigned(1101907360,32),
    to_unsigned(1102084072,32),
    to_unsigned(1102260774,32),
    to_unsigned(1102437465,32),
    to_unsigned(1102614147,32),
    to_unsigned(1102790819,32),
    to_unsigned(1102967480,32),
    to_unsigned(1103144132,32),
    to_unsigned(1103320773,32),
    to_unsigned(1103497404,32),
    to_unsigned(1103674025,32),
    to_unsigned(1103850635,32),
    to_unsigned(1104027236,32),
    to_unsigned(1104203826,32),
    to_unsigned(1104380407,32),
    to_unsigned(1104556977,32),
    to_unsigned(1104733537,32),
    to_unsigned(1104910087,32),
    to_unsigned(1105086626,32),
    to_unsigned(1105263156,32),
    to_unsigned(1105439675,32),
    to_unsigned(1105616185,32),
    to_unsigned(1105792684,32),
    to_unsigned(1105969173,32),
    to_unsigned(1106145651,32),
    to_unsigned(1106322120,32),
    to_unsigned(1106498578,32),
    to_unsigned(1106675026,32),
    to_unsigned(1106851464,32),
    to_unsigned(1107027892,32),
    to_unsigned(1107204310,32),
    to_unsigned(1107380717,32),
    to_unsigned(1107557115,32),
    to_unsigned(1107733502,32),
    to_unsigned(1107909879,32),
    to_unsigned(1108086246,32),
    to_unsigned(1108262602,32),
    to_unsigned(1108438949,32),
    to_unsigned(1108615285,32),
    to_unsigned(1108791611,32),
    to_unsigned(1108967927,32),
    to_unsigned(1109144232,32),
    to_unsigned(1109320528,32),
    to_unsigned(1109496813,32),
    to_unsigned(1109673088,32),
    to_unsigned(1109849353,32),
    to_unsigned(1110025608,32),
    to_unsigned(1110201852,32),
    to_unsigned(1110378087,32),
    to_unsigned(1110554311,32),
    to_unsigned(1110730524,32),
    to_unsigned(1110906728,32),
    to_unsigned(1111082921,32),
    to_unsigned(1111259105,32),
    to_unsigned(1111435278,32),
    to_unsigned(1111611440,32),
    to_unsigned(1111787593,32),
    to_unsigned(1111963735,32),
    to_unsigned(1112139867,32),
    to_unsigned(1112315989,32),
    to_unsigned(1112492101,32),
    to_unsigned(1112668202,32),
    to_unsigned(1112844294,32),
    to_unsigned(1113020375,32),
    to_unsigned(1113196445,32),
    to_unsigned(1113372506,32),
    to_unsigned(1113548556,32),
    to_unsigned(1113724596,32),
    to_unsigned(1113900626,32),
    to_unsigned(1114076646,32),
    to_unsigned(1114252655,32),
    to_unsigned(1114428654,32),
    to_unsigned(1114604643,32),
    to_unsigned(1114780622,32),
    to_unsigned(1114956590,32),
    to_unsigned(1115132548,32),
    to_unsigned(1115308496,32),
    to_unsigned(1115484433,32),
    to_unsigned(1115660361,32),
    to_unsigned(1115836278,32),
    to_unsigned(1116012185,32),
    to_unsigned(1116188081,32),
    to_unsigned(1116363968,32),
    to_unsigned(1116539844,32),
    to_unsigned(1116715710,32),
    to_unsigned(1116891565,32),
    to_unsigned(1117067410,32),
    to_unsigned(1117243245,32),
    to_unsigned(1117419070,32),
    to_unsigned(1117594885,32),
    to_unsigned(1117770689,32),
    to_unsigned(1117946483,32),
    to_unsigned(1118122266,32),
    to_unsigned(1118298040,32),
    to_unsigned(1118473803,32),
    to_unsigned(1118649556,32),
    to_unsigned(1118825298,32),
    to_unsigned(1119001030,32),
    to_unsigned(1119176752,32),
    to_unsigned(1119352464,32),
    to_unsigned(1119528165,32),
    to_unsigned(1119703856,32),
    to_unsigned(1119879537,32),
    to_unsigned(1120055208,32),
    to_unsigned(1120230868,32),
    to_unsigned(1120406518,32),
    to_unsigned(1120582157,32),
    to_unsigned(1120757787,32),
    to_unsigned(1120933406,32),
    to_unsigned(1121109014,32),
    to_unsigned(1121284613,32),
    to_unsigned(1121460201,32),
    to_unsigned(1121635779,32),
    to_unsigned(1121811346,32),
    to_unsigned(1121986903,32),
    to_unsigned(1122162450,32),
    to_unsigned(1122337987,32),
    to_unsigned(1122513513,32),
    to_unsigned(1122689029,32),
    to_unsigned(1122864534,32),
    to_unsigned(1123040030,32),
    to_unsigned(1123215515,32),
    to_unsigned(1123390989,32),
    to_unsigned(1123566454,32),
    to_unsigned(1123741907,32),
    to_unsigned(1123917351,32),
    to_unsigned(1124092784,32),
    to_unsigned(1124268207,32),
    to_unsigned(1124443620,32),
    to_unsigned(1124619022,32),
    to_unsigned(1124794414,32),
    to_unsigned(1124969796,32),
    to_unsigned(1125145167,32),
    to_unsigned(1125320528,32),
    to_unsigned(1125495879,32),
    to_unsigned(1125671219,32),
    to_unsigned(1125846549,32),
    to_unsigned(1126021868,32),
    to_unsigned(1126197178,32),
    to_unsigned(1126372476,32),
    to_unsigned(1126547765,32),
    to_unsigned(1126723043,32),
    to_unsigned(1126898311,32),
    to_unsigned(1127073568,32),
    to_unsigned(1127248815,32),
    to_unsigned(1127424052,32),
    to_unsigned(1127599278,32),
    to_unsigned(1127774494,32),
    to_unsigned(1127949700,32),
    to_unsigned(1128124895,32),
    to_unsigned(1128300080,32),
    to_unsigned(1128475255,32),
    to_unsigned(1128650419,32),
    to_unsigned(1128825573,32),
    to_unsigned(1129000716,32),
    to_unsigned(1129175849,32),
    to_unsigned(1129350972,32),
    to_unsigned(1129526084,32),
    to_unsigned(1129701186,32),
    to_unsigned(1129876277,32),
    to_unsigned(1130051358,32),
    to_unsigned(1130226429,32),
    to_unsigned(1130401489,32),
    to_unsigned(1130576539,32),
    to_unsigned(1130751579,32),
    to_unsigned(1130926608,32),
    to_unsigned(1131101627,32),
    to_unsigned(1131276635,32),
    to_unsigned(1131451633,32),
    to_unsigned(1131626620,32),
    to_unsigned(1131801598,32),
    to_unsigned(1131976564,32),
    to_unsigned(1132151521,32),
    to_unsigned(1132326467,32),
    to_unsigned(1132501402,32),
    to_unsigned(1132676327,32),
    to_unsigned(1132851242,32),
    to_unsigned(1133026146,32),
    to_unsigned(1133201040,32),
    to_unsigned(1133375924,32),
    to_unsigned(1133550797,32),
    to_unsigned(1133725659,32),
    to_unsigned(1133900511,32),
    to_unsigned(1134075353,32),
    to_unsigned(1134250185,32),
    to_unsigned(1134425005,32),
    to_unsigned(1134599816,32),
    to_unsigned(1134774616,32),
    to_unsigned(1134949406,32),
    to_unsigned(1135124185,32),
    to_unsigned(1135298954,32),
    to_unsigned(1135473712,32),
    to_unsigned(1135648460,32),
    to_unsigned(1135823197,32),
    to_unsigned(1135997924,32),
    to_unsigned(1136172641,32),
    to_unsigned(1136347347,32),
    to_unsigned(1136522043,32),
    to_unsigned(1136696728,32),
    to_unsigned(1136871403,32),
    to_unsigned(1137046067,32),
    to_unsigned(1137220721,32),
    to_unsigned(1137395365,32),
    to_unsigned(1137569998,32),
    to_unsigned(1137744620,32),
    to_unsigned(1137919232,32),
    to_unsigned(1138093834,32),
    to_unsigned(1138268425,32),
    to_unsigned(1138443006,32),
    to_unsigned(1138617576,32),
    to_unsigned(1138792136,32),
    to_unsigned(1138966685,32),
    to_unsigned(1139141224,32),
    to_unsigned(1139315752,32),
    to_unsigned(1139490270,32),
    to_unsigned(1139664777,32),
    to_unsigned(1139839274,32),
    to_unsigned(1140013761,32),
    to_unsigned(1140188237,32),
    to_unsigned(1140362702,32),
    to_unsigned(1140537157,32),
    to_unsigned(1140711602,32),
    to_unsigned(1140886036,32),
    to_unsigned(1141060459,32),
    to_unsigned(1141234873,32),
    to_unsigned(1141409275,32),
    to_unsigned(1141583667,32),
    to_unsigned(1141758049,32),
    to_unsigned(1141932420,32),
    to_unsigned(1142106781,32),
    to_unsigned(1142281131,32),
    to_unsigned(1142455470,32),
    to_unsigned(1142629799,32),
    to_unsigned(1142804118,32),
    to_unsigned(1142978426,32),
    to_unsigned(1143152724,32),
    to_unsigned(1143327011,32),
    to_unsigned(1143501287,32),
    to_unsigned(1143675553,32),
    to_unsigned(1143849809,32),
    to_unsigned(1144024054,32),
    to_unsigned(1144198288,32),
    to_unsigned(1144372512,32),
    to_unsigned(1144546726,32),
    to_unsigned(1144720929,32),
    to_unsigned(1144895121,32),
    to_unsigned(1145069303,32),
    to_unsigned(1145243475,32),
    to_unsigned(1145417636,32),
    to_unsigned(1145591786,32),
    to_unsigned(1145765926,32),
    to_unsigned(1145940055,32),
    to_unsigned(1146114174,32),
    to_unsigned(1146288282,32),
    to_unsigned(1146462380,32),
    to_unsigned(1146636467,32),
    to_unsigned(1146810543,32),
    to_unsigned(1146984609,32),
    to_unsigned(1147158665,32),
    to_unsigned(1147332710,32),
    to_unsigned(1147506744,32),
    to_unsigned(1147680768,32),
    to_unsigned(1147854782,32),
    to_unsigned(1148028784,32),
    to_unsigned(1148202777,32),
    to_unsigned(1148376758,32),
    to_unsigned(1148550729,32),
    to_unsigned(1148724690,32),
    to_unsigned(1148898640,32),
    to_unsigned(1149072579,32),
    to_unsigned(1149246508,32),
    to_unsigned(1149420427,32),
    to_unsigned(1149594334,32),
    to_unsigned(1149768231,32),
    to_unsigned(1149942118,32),
    to_unsigned(1150115994,32),
    to_unsigned(1150289860,32),
    to_unsigned(1150463714,32),
    to_unsigned(1150637559,32),
    to_unsigned(1150811393,32),
    to_unsigned(1150985216,32),
    to_unsigned(1151159028,32),
    to_unsigned(1151332830,32),
    to_unsigned(1151506622,32),
    to_unsigned(1151680403,32),
    to_unsigned(1151854173,32),
    to_unsigned(1152027932,32),
    to_unsigned(1152201682,32),
    to_unsigned(1152375420,32),
    to_unsigned(1152549148,32),
    to_unsigned(1152722865,32),
    to_unsigned(1152896572,32),
    to_unsigned(1153070268,32),
    to_unsigned(1153243954,32),
    to_unsigned(1153417628,32),
    to_unsigned(1153591293,32),
    to_unsigned(1153764946,32),
    to_unsigned(1153938590,32),
    to_unsigned(1154112222,32),
    to_unsigned(1154285844,32),
    to_unsigned(1154459455,32),
    to_unsigned(1154633056,32),
    to_unsigned(1154806646,32),
    to_unsigned(1154980225,32),
    to_unsigned(1155153794,32),
    to_unsigned(1155327352,32),
    to_unsigned(1155500900,32),
    to_unsigned(1155674437,32),
    to_unsigned(1155847963,32),
    to_unsigned(1156021479,32),
    to_unsigned(1156194984,32),
    to_unsigned(1156368478,32),
    to_unsigned(1156541962,32),
    to_unsigned(1156715435,32),
    to_unsigned(1156888898,32),
    to_unsigned(1157062350,32),
    to_unsigned(1157235791,32),
    to_unsigned(1157409222,32),
    to_unsigned(1157582642,32),
    to_unsigned(1157756051,32),
    to_unsigned(1157929450,32),
    to_unsigned(1158102838,32),
    to_unsigned(1158276216,32),
    to_unsigned(1158449582,32),
    to_unsigned(1158622939,32),
    to_unsigned(1158796284,32),
    to_unsigned(1158969619,32),
    to_unsigned(1159142943,32),
    to_unsigned(1159316257,32),
    to_unsigned(1159489560,32),
    to_unsigned(1159662852,32),
    to_unsigned(1159836133,32),
    to_unsigned(1160009404,32),
    to_unsigned(1160182665,32),
    to_unsigned(1160355914,32),
    to_unsigned(1160529153,32),
    to_unsigned(1160702381,32),
    to_unsigned(1160875599,32),
    to_unsigned(1161048806,32),
    to_unsigned(1161222002,32),
    to_unsigned(1161395188,32),
    to_unsigned(1161568362,32),
    to_unsigned(1161741527,32),
    to_unsigned(1161914680,32),
    to_unsigned(1162087823,32),
    to_unsigned(1162260955,32),
    to_unsigned(1162434077,32),
    to_unsigned(1162607188,32),
    to_unsigned(1162780288,32),
    to_unsigned(1162953377,32),
    to_unsigned(1163126456,32),
    to_unsigned(1163299524,32),
    to_unsigned(1163472581,32),
    to_unsigned(1163645628,32),
    to_unsigned(1163818664,32),
    to_unsigned(1163991689,32),
    to_unsigned(1164164704,32),
    to_unsigned(1164337708,32),
    to_unsigned(1164510701,32),
    to_unsigned(1164683683,32),
    to_unsigned(1164856655,32),
    to_unsigned(1165029616,32),
    to_unsigned(1165202566,32),
    to_unsigned(1165375506,32),
    to_unsigned(1165548435,32),
    to_unsigned(1165721353,32),
    to_unsigned(1165894261,32),
    to_unsigned(1166067157,32),
    to_unsigned(1166240043,32),
    to_unsigned(1166412919,32),
    to_unsigned(1166585783,32),
    to_unsigned(1166758637,32),
    to_unsigned(1166931480,32),
    to_unsigned(1167104313,32),
    to_unsigned(1167277135,32),
    to_unsigned(1167449946,32),
    to_unsigned(1167622746,32),
    to_unsigned(1167795535,32),
    to_unsigned(1167968314,32),
    to_unsigned(1168141082,32),
    to_unsigned(1168313839,32),
    to_unsigned(1168486586,32),
    to_unsigned(1168659322,32),
    to_unsigned(1168832047,32),
    to_unsigned(1169004761,32),
    to_unsigned(1169177465,32),
    to_unsigned(1169350158,32),
    to_unsigned(1169522840,32),
    to_unsigned(1169695511,32),
    to_unsigned(1169868172,32),
    to_unsigned(1170040822,32),
    to_unsigned(1170213461,32),
    to_unsigned(1170386089,32),
    to_unsigned(1170558707,32),
    to_unsigned(1170731314,32),
    to_unsigned(1170903910,32),
    to_unsigned(1171076495,32),
    to_unsigned(1171249069,32),
    to_unsigned(1171421633,32),
    to_unsigned(1171594186,32),
    to_unsigned(1171766728,32),
    to_unsigned(1171939260,32),
    to_unsigned(1172111781,32),
    to_unsigned(1172284291,32),
    to_unsigned(1172456790,32),
    to_unsigned(1172629278,32),
    to_unsigned(1172801756,32),
    to_unsigned(1172974222,32),
    to_unsigned(1173146678,32),
    to_unsigned(1173319124,32),
    to_unsigned(1173491558,32),
    to_unsigned(1173663982,32),
    to_unsigned(1173836395,32),
    to_unsigned(1174008797,32),
    to_unsigned(1174181188,32),
    to_unsigned(1174353569,32),
    to_unsigned(1174525938,32),
    to_unsigned(1174698297,32),
    to_unsigned(1174870645,32),
    to_unsigned(1175042983,32),
    to_unsigned(1175215309,32),
    to_unsigned(1175387625,32),
    to_unsigned(1175559930,32),
    to_unsigned(1175732224,32),
    to_unsigned(1175904507,32),
    to_unsigned(1176076780,32),
    to_unsigned(1176249041,32),
    to_unsigned(1176421292,32),
    to_unsigned(1176593532,32),
    to_unsigned(1176765762,32),
    to_unsigned(1176937980,32),
    to_unsigned(1177110188,32),
    to_unsigned(1177282384,32),
    to_unsigned(1177454570,32),
    to_unsigned(1177626746,32),
    to_unsigned(1177798910,32),
    to_unsigned(1177971063,32),
    to_unsigned(1178143206,32),
    to_unsigned(1178315338,32),
    to_unsigned(1178487459,32),
    to_unsigned(1178659569,32),
    to_unsigned(1178831668,32),
    to_unsigned(1179003757,32),
    to_unsigned(1179175835,32),
    to_unsigned(1179347901,32),
    to_unsigned(1179519957,32),
    to_unsigned(1179692002,32),
    to_unsigned(1179864037,32),
    to_unsigned(1180036060,32),
    to_unsigned(1180208073,32),
    to_unsigned(1180380075,32),
    to_unsigned(1180552066,32),
    to_unsigned(1180724046,32),
    to_unsigned(1180896015,32),
    to_unsigned(1181067973,32),
    to_unsigned(1181239921,32),
    to_unsigned(1181411857,32),
    to_unsigned(1181583783,32),
    to_unsigned(1181755698,32),
    to_unsigned(1181927602,32),
    to_unsigned(1182099495,32),
    to_unsigned(1182271378,32),
    to_unsigned(1182443249,32),
    to_unsigned(1182615110,32),
    to_unsigned(1182786959,32),
    to_unsigned(1182958798,32),
    to_unsigned(1183130626,32),
    to_unsigned(1183302443,32),
    to_unsigned(1183474249,32),
    to_unsigned(1183646045,32),
    to_unsigned(1183817829,32),
    to_unsigned(1183989603,32),
    to_unsigned(1184161366,32),
    to_unsigned(1184333117,32),
    to_unsigned(1184504858,32),
    to_unsigned(1184676588,32),
    to_unsigned(1184848308,32),
    to_unsigned(1185020016,32),
    to_unsigned(1185191713,32),
    to_unsigned(1185363400,32),
    to_unsigned(1185535075,32),
    to_unsigned(1185706740,32),
    to_unsigned(1185878394,32),
    to_unsigned(1186050037,32),
    to_unsigned(1186221669,32),
    to_unsigned(1186393290,32),
    to_unsigned(1186564900,32),
    to_unsigned(1186736499,32),
    to_unsigned(1186908087,32),
    to_unsigned(1187079665,32),
    to_unsigned(1187251231,32),
    to_unsigned(1187422787,32),
    to_unsigned(1187594332,32),
    to_unsigned(1187765866,32),
    to_unsigned(1187937388,32),
    to_unsigned(1188108900,32),
    to_unsigned(1188280401,32),
    to_unsigned(1188451892,32),
    to_unsigned(1188623371,32),
    to_unsigned(1188794839,32),
    to_unsigned(1188966296,32),
    to_unsigned(1189137743,32),
    to_unsigned(1189309178,32),
    to_unsigned(1189480603,32),
    to_unsigned(1189652016,32),
    to_unsigned(1189823419,32),
    to_unsigned(1189994811,32),
    to_unsigned(1190166192,32),
    to_unsigned(1190337561,32),
    to_unsigned(1190508920,32),
    to_unsigned(1190680268,32),
    to_unsigned(1190851605,32),
    to_unsigned(1191022931,32),
    to_unsigned(1191194247,32),
    to_unsigned(1191365551,32),
    to_unsigned(1191536844,32),
    to_unsigned(1191708126,32),
    to_unsigned(1191879398,32),
    to_unsigned(1192050658,32),
    to_unsigned(1192221907,32),
    to_unsigned(1192393146,32),
    to_unsigned(1192564373,32),
    to_unsigned(1192735590,32),
    to_unsigned(1192906796,32),
    to_unsigned(1193077990,32),
    to_unsigned(1193249174,32),
    to_unsigned(1193420346,32),
    to_unsigned(1193591508,32),
    to_unsigned(1193762659,32),
    to_unsigned(1193933799,32),
    to_unsigned(1194104927,32),
    to_unsigned(1194276045,32),
    to_unsigned(1194447152,32),
    to_unsigned(1194618248,32),
    to_unsigned(1194789333,32),
    to_unsigned(1194960407,32),
    to_unsigned(1195131470,32),
    to_unsigned(1195302522,32),
    to_unsigned(1195473563,32),
    to_unsigned(1195644593,32),
    to_unsigned(1195815611,32),
    to_unsigned(1195986619,32),
    to_unsigned(1196157616,32),
    to_unsigned(1196328602,32),
    to_unsigned(1196499577,32),
    to_unsigned(1196670541,32),
    to_unsigned(1196841494,32),
    to_unsigned(1197012436,32),
    to_unsigned(1197183367,32),
    to_unsigned(1197354287,32),
    to_unsigned(1197525196,32),
    to_unsigned(1197696094,32),
    to_unsigned(1197866981,32),
    to_unsigned(1198037857,32),
    to_unsigned(1198208722,32),
    to_unsigned(1198379576,32),
    to_unsigned(1198550419,32),
    to_unsigned(1198721251,32),
    to_unsigned(1198892072,32),
    to_unsigned(1199062881,32),
    to_unsigned(1199233680,32),
    to_unsigned(1199404468,32),
    to_unsigned(1199575245,32),
    to_unsigned(1199746011,32),
    to_unsigned(1199916765,32),
    to_unsigned(1200087509,32),
    to_unsigned(1200258242,32),
    to_unsigned(1200428963,32),
    to_unsigned(1200599674,32),
    to_unsigned(1200770374,32),
    to_unsigned(1200941062,32),
    to_unsigned(1201111740,32),
    to_unsigned(1201282406,32),
    to_unsigned(1201453061,32),
    to_unsigned(1201623706,32),
    to_unsigned(1201794339,32),
    to_unsigned(1201964961,32),
    to_unsigned(1202135573,32),
    to_unsigned(1202306173,32),
    to_unsigned(1202476762,32),
    to_unsigned(1202647340,32),
    to_unsigned(1202817907,32),
    to_unsigned(1202988463,32),
    to_unsigned(1203159008,32),
    to_unsigned(1203329542,32),
    to_unsigned(1203500064,32),
    to_unsigned(1203670576,32),
    to_unsigned(1203841077,32),
    to_unsigned(1204011566,32),
    to_unsigned(1204182045,32),
    to_unsigned(1204352512,32),
    to_unsigned(1204522969,32),
    to_unsigned(1204693414,32),
    to_unsigned(1204863848,32),
    to_unsigned(1205034271,32),
    to_unsigned(1205204684,32),
    to_unsigned(1205375085,32),
    to_unsigned(1205545474,32),
    to_unsigned(1205715853,32),
    to_unsigned(1205886221,32),
    to_unsigned(1206056578,32),
    to_unsigned(1206226923,32),
    to_unsigned(1206397258,32),
    to_unsigned(1206567581,32),
    to_unsigned(1206737894,32),
    to_unsigned(1206908195,32),
    to_unsigned(1207078485,32),
    to_unsigned(1207248764,32),
    to_unsigned(1207419032,32),
    to_unsigned(1207589289,32),
    to_unsigned(1207759535,32),
    to_unsigned(1207929769,32),
    to_unsigned(1208099993,32),
    to_unsigned(1208270205,32),
    to_unsigned(1208440407,32),
    to_unsigned(1208610597,32),
    to_unsigned(1208780776,32),
    to_unsigned(1208950944,32),
    to_unsigned(1209121101,32),
    to_unsigned(1209291247,32),
    to_unsigned(1209461381,32),
    to_unsigned(1209631505,32),
    to_unsigned(1209801617,32),
    to_unsigned(1209971719,32),
    to_unsigned(1210141809,32),
    to_unsigned(1210311888,32),
    to_unsigned(1210481956,32),
    to_unsigned(1210652013,32),
    to_unsigned(1210822058,32),
    to_unsigned(1210992093,32),
    to_unsigned(1211162116,32),
    to_unsigned(1211332129,32),
    to_unsigned(1211502130,32),
    to_unsigned(1211672120,32),
    to_unsigned(1211842099,32),
    to_unsigned(1212012066,32),
    to_unsigned(1212182023,32),
    to_unsigned(1212351968,32),
    to_unsigned(1212521903,32),
    to_unsigned(1212691826,32),
    to_unsigned(1212861738,32),
    to_unsigned(1213031639,32),
    to_unsigned(1213201529,32),
    to_unsigned(1213371407,32),
    to_unsigned(1213541275,32),
    to_unsigned(1213711131,32),
    to_unsigned(1213880976,32),
    to_unsigned(1214050810,32),
    to_unsigned(1214220633,32),
    to_unsigned(1214390444,32),
    to_unsigned(1214560245,32),
    to_unsigned(1214730034,32),
    to_unsigned(1214899812,32),
    to_unsigned(1215069579,32),
    to_unsigned(1215239335,32),
    to_unsigned(1215409080,32),
    to_unsigned(1215578813,32),
    to_unsigned(1215748535,32),
    to_unsigned(1215918247,32),
    to_unsigned(1216087946,32),
    to_unsigned(1216257635,32),
    to_unsigned(1216427313,32),
    to_unsigned(1216596979,32),
    to_unsigned(1216766634,32),
    to_unsigned(1216936278,32),
    to_unsigned(1217105911,32),
    to_unsigned(1217275533,32),
    to_unsigned(1217445143,32),
    to_unsigned(1217614743,32),
    to_unsigned(1217784331,32),
    to_unsigned(1217953908,32),
    to_unsigned(1218123473,32),
    to_unsigned(1218293028,32),
    to_unsigned(1218462571,32),
    to_unsigned(1218632103,32),
    to_unsigned(1218801624,32),
    to_unsigned(1218971134,32),
    to_unsigned(1219140632,32),
    to_unsigned(1219310120,32),
    to_unsigned(1219479596,32),
    to_unsigned(1219649061,32),
    to_unsigned(1219818514,32),
    to_unsigned(1219987957,32),
    to_unsigned(1220157388,32),
    to_unsigned(1220326808,32),
    to_unsigned(1220496217,32),
    to_unsigned(1220665615,32),
    to_unsigned(1220835001,32),
    to_unsigned(1221004376,32),
    to_unsigned(1221173740,32),
    to_unsigned(1221343093,32),
    to_unsigned(1221512434,32),
    to_unsigned(1221681764,32),
    to_unsigned(1221851083,32),
    to_unsigned(1222020391,32),
    to_unsigned(1222189688,32),
    to_unsigned(1222358973,32),
    to_unsigned(1222528247,32),
    to_unsigned(1222697510,32),
    to_unsigned(1222866762,32),
    to_unsigned(1223036002,32),
    to_unsigned(1223205231,32),
    to_unsigned(1223374449,32),
    to_unsigned(1223543656,32),
    to_unsigned(1223712851,32),
    to_unsigned(1223882035,32),
    to_unsigned(1224051208,32),
    to_unsigned(1224220370,32),
    to_unsigned(1224389520,32),
    to_unsigned(1224558659,32),
    to_unsigned(1224727787,32),
    to_unsigned(1224896904,32),
    to_unsigned(1225066009,32),
    to_unsigned(1225235103,32),
    to_unsigned(1225404186,32),
    to_unsigned(1225573258,32),
    to_unsigned(1225742318,32),
    to_unsigned(1225911367,32),
    to_unsigned(1226080405,32),
    to_unsigned(1226249431,32),
    to_unsigned(1226418446,32),
    to_unsigned(1226587450,32),
    to_unsigned(1226756443,32),
    to_unsigned(1226925424,32),
    to_unsigned(1227094395,32),
    to_unsigned(1227263353,32),
    to_unsigned(1227432301,32),
    to_unsigned(1227601237,32),
    to_unsigned(1227770162,32),
    to_unsigned(1227939076,32),
    to_unsigned(1228107978,32),
    to_unsigned(1228276870,32),
    to_unsigned(1228445749,32),
    to_unsigned(1228614618,32),
    to_unsigned(1228783475,32),
    to_unsigned(1228952321,32),
    to_unsigned(1229121156,32),
    to_unsigned(1229289979,32),
    to_unsigned(1229458791,32),
    to_unsigned(1229627592,32),
    to_unsigned(1229796382,32),
    to_unsigned(1229965160,32),
    to_unsigned(1230133927,32),
    to_unsigned(1230302682,32),
    to_unsigned(1230471426,32),
    to_unsigned(1230640159,32),
    to_unsigned(1230808881,32),
    to_unsigned(1230977591,32),
    to_unsigned(1231146290,32),
    to_unsigned(1231314978,32),
    to_unsigned(1231483654,32),
    to_unsigned(1231652319,32),
    to_unsigned(1231820973,32),
    to_unsigned(1231989616,32),
    to_unsigned(1232158247,32),
    to_unsigned(1232326866,32),
    to_unsigned(1232495475,32),
    to_unsigned(1232664072,32),
    to_unsigned(1232832658,32),
    to_unsigned(1233001232,32),
    to_unsigned(1233169795,32),
    to_unsigned(1233338347,32),
    to_unsigned(1233506887,32),
    to_unsigned(1233675417,32),
    to_unsigned(1233843934,32),
    to_unsigned(1234012441,32),
    to_unsigned(1234180936,32),
    to_unsigned(1234349419,32),
    to_unsigned(1234517892,32),
    to_unsigned(1234686353,32),
    to_unsigned(1234854803,32),
    to_unsigned(1235023241,32),
    to_unsigned(1235191668,32),
    to_unsigned(1235360084,32),
    to_unsigned(1235528488,32),
    to_unsigned(1235696881,32),
    to_unsigned(1235865262,32),
    to_unsigned(1236033632,32),
    to_unsigned(1236201991,32),
    to_unsigned(1236370339,32),
    to_unsigned(1236538675,32),
    to_unsigned(1236707000,32),
    to_unsigned(1236875313,32),
    to_unsigned(1237043615,32),
    to_unsigned(1237211906,32),
    to_unsigned(1237380185,32),
    to_unsigned(1237548453,32),
    to_unsigned(1237716709,32),
    to_unsigned(1237884954,32),
    to_unsigned(1238053188,32),
    to_unsigned(1238221411,32),
    to_unsigned(1238389622,32),
    to_unsigned(1238557821,32),
    to_unsigned(1238726009,32),
    to_unsigned(1238894186,32),
    to_unsigned(1239062352,32),
    to_unsigned(1239230506,32),
    to_unsigned(1239398648,32),
    to_unsigned(1239566780,32),
    to_unsigned(1239734900,32),
    to_unsigned(1239903008,32),
    to_unsigned(1240071105,32),
    to_unsigned(1240239191,32),
    to_unsigned(1240407265,32),
    to_unsigned(1240575328,32),
    to_unsigned(1240743380,32),
    to_unsigned(1240911420,32),
    to_unsigned(1241079448,32),
    to_unsigned(1241247466,32),
    to_unsigned(1241415472,32),
    to_unsigned(1241583466,32),
    to_unsigned(1241751449,32),
    to_unsigned(1241919421,32),
    to_unsigned(1242087381,32),
    to_unsigned(1242255330,32),
    to_unsigned(1242423267,32),
    to_unsigned(1242591193,32),
    to_unsigned(1242759108,32),
    to_unsigned(1242927011,32),
    to_unsigned(1243094902,32),
    to_unsigned(1243262783,32),
    to_unsigned(1243430651,32),
    to_unsigned(1243598509,32),
    to_unsigned(1243766355,32),
    to_unsigned(1243934189,32),
    to_unsigned(1244102012,32),
    to_unsigned(1244269824,32),
    to_unsigned(1244437624,32),
    to_unsigned(1244605413,32),
    to_unsigned(1244773190,32),
    to_unsigned(1244940956,32),
    to_unsigned(1245108711,32),
    to_unsigned(1245276454,32),
    to_unsigned(1245444185,32),
    to_unsigned(1245611906,32),
    to_unsigned(1245779614,32),
    to_unsigned(1245947312,32),
    to_unsigned(1246114997,32),
    to_unsigned(1246282672,32),
    to_unsigned(1246450334,32),
    to_unsigned(1246617986,32),
    to_unsigned(1246785626,32),
    to_unsigned(1246953254,32),
    to_unsigned(1247120871,32),
    to_unsigned(1247288477,32),
    to_unsigned(1247456071,32),
    to_unsigned(1247623654,32),
    to_unsigned(1247791225,32),
    to_unsigned(1247958785,32),
    to_unsigned(1248126333,32),
    to_unsigned(1248293870,32),
    to_unsigned(1248461395,32),
    to_unsigned(1248628909,32),
    to_unsigned(1248796411,32),
    to_unsigned(1248963902,32),
    to_unsigned(1249131381,32),
    to_unsigned(1249298849,32),
    to_unsigned(1249466305,32),
    to_unsigned(1249633750,32),
    to_unsigned(1249801184,32),
    to_unsigned(1249968606,32),
    to_unsigned(1250136016,32),
    to_unsigned(1250303415,32),
    to_unsigned(1250470803,32),
    to_unsigned(1250638179,32),
    to_unsigned(1250805543,32),
    to_unsigned(1250972896,32),
    to_unsigned(1251140238,32),
    to_unsigned(1251307568,32),
    to_unsigned(1251474886,32),
    to_unsigned(1251642193,32),
    to_unsigned(1251809489,32),
    to_unsigned(1251976773,32),
    to_unsigned(1252144045,32),
    to_unsigned(1252311306,32),
    to_unsigned(1252478555,32),
    to_unsigned(1252645793,32),
    to_unsigned(1252813020,32),
    to_unsigned(1252980235,32),
    to_unsigned(1253147438,32),
    to_unsigned(1253314630,32),
    to_unsigned(1253481810,32),
    to_unsigned(1253648979,32),
    to_unsigned(1253816136,32),
    to_unsigned(1253983282,32),
    to_unsigned(1254150416,32),
    to_unsigned(1254317539,32),
    to_unsigned(1254484650,32),
    to_unsigned(1254651750,32),
    to_unsigned(1254818838,32),
    to_unsigned(1254985915,32),
    to_unsigned(1255152980,32),
    to_unsigned(1255320033,32),
    to_unsigned(1255487075,32),
    to_unsigned(1255654106,32),
    to_unsigned(1255821125,32),
    to_unsigned(1255988132,32),
    to_unsigned(1256155128,32),
    to_unsigned(1256322112,32),
    to_unsigned(1256489085,32),
    to_unsigned(1256656046,32),
    to_unsigned(1256822996,32),
    to_unsigned(1256989934,32),
    to_unsigned(1257156860,32),
    to_unsigned(1257323775,32),
    to_unsigned(1257490678,32),
    to_unsigned(1257657570,32),
    to_unsigned(1257824451,32),
    to_unsigned(1257991319,32),
    to_unsigned(1258158176,32),
    to_unsigned(1258325022,32),
    to_unsigned(1258491856,32),
    to_unsigned(1258658679,32),
    to_unsigned(1258825489,32),
    to_unsigned(1258992289,32),
    to_unsigned(1259159077,32),
    to_unsigned(1259325853,32),
    to_unsigned(1259492617,32),
    to_unsigned(1259659370,32),
    to_unsigned(1259826112,32),
    to_unsigned(1259992842,32),
    to_unsigned(1260159560,32),
    to_unsigned(1260326267,32),
    to_unsigned(1260492962,32),
    to_unsigned(1260659645,32),
    to_unsigned(1260826317,32),
    to_unsigned(1260992977,32),
    to_unsigned(1261159626,32),
    to_unsigned(1261326263,32),
    to_unsigned(1261492889,32),
    to_unsigned(1261659503,32),
    to_unsigned(1261826105,32),
    to_unsigned(1261992696,32),
    to_unsigned(1262159275,32),
    to_unsigned(1262325843,32),
    to_unsigned(1262492399,32),
    to_unsigned(1262658943,32),
    to_unsigned(1262825476,32),
    to_unsigned(1262991997,32),
    to_unsigned(1263158507,32),
    to_unsigned(1263325005,32),
    to_unsigned(1263491491,32),
    to_unsigned(1263657966,32),
    to_unsigned(1263824429,32),
    to_unsigned(1263990880,32),
    to_unsigned(1264157320,32),
    to_unsigned(1264323748,32),
    to_unsigned(1264490165,32),
    to_unsigned(1264656570,32),
    to_unsigned(1264822963,32),
    to_unsigned(1264989345,32),
    to_unsigned(1265155715,32),
    to_unsigned(1265322074,32),
    to_unsigned(1265488421,32),
    to_unsigned(1265654756,32),
    to_unsigned(1265821079,32),
    to_unsigned(1265987391,32),
    to_unsigned(1266153692,32),
    to_unsigned(1266319980,32),
    to_unsigned(1266486257,32),
    to_unsigned(1266652523,32),
    to_unsigned(1266818777,32),
    to_unsigned(1266985019,32),
    to_unsigned(1267151249,32),
    to_unsigned(1267317468,32),
    to_unsigned(1267483675,32),
    to_unsigned(1267649871,32),
    to_unsigned(1267816055,32),
    to_unsigned(1267982227,32),
    to_unsigned(1268148387,32),
    to_unsigned(1268314536,32),
    to_unsigned(1268480673,32),
    to_unsigned(1268646799,32),
    to_unsigned(1268812913,32),
    to_unsigned(1268979015,32),
    to_unsigned(1269145106,32),
    to_unsigned(1269311185,32),
    to_unsigned(1269477252,32),
    to_unsigned(1269643308,32),
    to_unsigned(1269809352,32),
    to_unsigned(1269975384,32),
    to_unsigned(1270141404,32),
    to_unsigned(1270307413,32),
    to_unsigned(1270473411,32),
    to_unsigned(1270639396,32),
    to_unsigned(1270805370,32),
    to_unsigned(1270971332,32),
    to_unsigned(1271137283,32),
    to_unsigned(1271303222,32),
    to_unsigned(1271469149,32),
    to_unsigned(1271635064,32),
    to_unsigned(1271800968,32),
    to_unsigned(1271966860,32),
    to_unsigned(1272132740,32),
    to_unsigned(1272298609,32),
    to_unsigned(1272464466,32),
    to_unsigned(1272630311,32),
    to_unsigned(1272796145,32),
    to_unsigned(1272961967,32),
    to_unsigned(1273127777,32),
    to_unsigned(1273293576,32),
    to_unsigned(1273459362,32),
    to_unsigned(1273625137,32),
    to_unsigned(1273790901,32),
    to_unsigned(1273956652,32),
    to_unsigned(1274122392,32),
    to_unsigned(1274288121,32),
    to_unsigned(1274453837,32),
    to_unsigned(1274619542,32),
    to_unsigned(1274785235,32),
    to_unsigned(1274950917,32),
    to_unsigned(1275116586,32),
    to_unsigned(1275282244,32),
    to_unsigned(1275447890,32),
    to_unsigned(1275613525,32),
    to_unsigned(1275779148,32),
    to_unsigned(1275944759,32),
    to_unsigned(1276110358,32),
    to_unsigned(1276275946,32),
    to_unsigned(1276441522,32),
    to_unsigned(1276607086,32),
    to_unsigned(1276772638,32),
    to_unsigned(1276938179,32),
    to_unsigned(1277103708,32),
    to_unsigned(1277269225,32),
    to_unsigned(1277434730,32),
    to_unsigned(1277600224,32),
    to_unsigned(1277765706,32),
    to_unsigned(1277931176,32),
    to_unsigned(1278096635,32),
    to_unsigned(1278262081,32),
    to_unsigned(1278427516,32),
    to_unsigned(1278592940,32),
    to_unsigned(1278758351,32),
    to_unsigned(1278923751,32),
    to_unsigned(1279089139,32),
    to_unsigned(1279254515,32),
    to_unsigned(1279419879,32),
    to_unsigned(1279585232,32),
    to_unsigned(1279750573,32),
    to_unsigned(1279915902,32),
    to_unsigned(1280081220,32),
    to_unsigned(1280246525,32),
    to_unsigned(1280411819,32),
    to_unsigned(1280577101,32),
    to_unsigned(1280742371,32),
    to_unsigned(1280907630,32),
    to_unsigned(1281072877,32),
    to_unsigned(1281238112,32),
    to_unsigned(1281403335,32),
    to_unsigned(1281568546,32),
    to_unsigned(1281733746,32),
    to_unsigned(1281898934,32),
    to_unsigned(1282064110,32),
    to_unsigned(1282229274,32),
    to_unsigned(1282394427,32),
    to_unsigned(1282559568,32),
    to_unsigned(1282724697,32),
    to_unsigned(1282889814,32),
    to_unsigned(1283054919,32),
    to_unsigned(1283220013,32),
    to_unsigned(1283385094,32),
    to_unsigned(1283550164,32),
    to_unsigned(1283715223,32),
    to_unsigned(1283880269,32),
    to_unsigned(1284045304,32),
    to_unsigned(1284210326,32),
    to_unsigned(1284375337,32),
    to_unsigned(1284540337,32),
    to_unsigned(1284705324,32),
    to_unsigned(1284870299,32),
    to_unsigned(1285035263,32),
    to_unsigned(1285200215,32),
    to_unsigned(1285365155,32),
    to_unsigned(1285530084,32),
    to_unsigned(1285695000,32),
    to_unsigned(1285859905,32),
    to_unsigned(1286024798,32),
    to_unsigned(1286189679,32),
    to_unsigned(1286354548,32),
    to_unsigned(1286519405,32),
    to_unsigned(1286684251,32),
    to_unsigned(1286849085,32),
    to_unsigned(1287013906,32),
    to_unsigned(1287178717,32),
    to_unsigned(1287343515,32),
    to_unsigned(1287508301,32),
    to_unsigned(1287673076,32),
    to_unsigned(1287837838,32),
    to_unsigned(1288002589,32),
    to_unsigned(1288167328,32),
    to_unsigned(1288332056,32),
    to_unsigned(1288496771,32),
    to_unsigned(1288661475,32),
    to_unsigned(1288826166,32),
    to_unsigned(1288990846,32),
    to_unsigned(1289155514,32),
    to_unsigned(1289320170,32),
    to_unsigned(1289484815,32),
    to_unsigned(1289649447,32),
    to_unsigned(1289814068,32),
    to_unsigned(1289978676,32),
    to_unsigned(1290143273,32),
    to_unsigned(1290307858,32),
    to_unsigned(1290472431,32),
    to_unsigned(1290636993,32),
    to_unsigned(1290801542,32),
    to_unsigned(1290966080,32),
    to_unsigned(1291130605,32),
    to_unsigned(1291295119,32),
    to_unsigned(1291459621,32),
    to_unsigned(1291624111,32),
    to_unsigned(1291788589,32),
    to_unsigned(1291953056,32),
    to_unsigned(1292117510,32),
    to_unsigned(1292281953,32),
    to_unsigned(1292446384,32),
    to_unsigned(1292610802,32),
    to_unsigned(1292775209,32),
    to_unsigned(1292939604,32),
    to_unsigned(1293103988,32),
    to_unsigned(1293268359,32),
    to_unsigned(1293432718,32),
    to_unsigned(1293597066,32),
    to_unsigned(1293761402,32),
    to_unsigned(1293925725,32),
    to_unsigned(1294090037,32),
    to_unsigned(1294254337,32),
    to_unsigned(1294418625,32),
    to_unsigned(1294582901,32),
    to_unsigned(1294747166,32),
    to_unsigned(1294911418,32),
    to_unsigned(1295075658,32),
    to_unsigned(1295239887,32),
    to_unsigned(1295404104,32),
    to_unsigned(1295568308,32),
    to_unsigned(1295732501,32),
    to_unsigned(1295896682,32),
    to_unsigned(1296060851,32),
    to_unsigned(1296225008,32),
    to_unsigned(1296389153,32),
    to_unsigned(1296553287,32),
    to_unsigned(1296717408,32),
    to_unsigned(1296881517,32),
    to_unsigned(1297045615,32),
    to_unsigned(1297209701,32),
    to_unsigned(1297373774,32),
    to_unsigned(1297537836,32),
    to_unsigned(1297701886,32),
    to_unsigned(1297865924,32),
    to_unsigned(1298029950,32),
    to_unsigned(1298193964,32),
    to_unsigned(1298357966,32),
    to_unsigned(1298521956,32),
    to_unsigned(1298685934,32),
    to_unsigned(1298849900,32),
    to_unsigned(1299013855,32),
    to_unsigned(1299177797,32),
    to_unsigned(1299341728,32),
    to_unsigned(1299505646,32),
    to_unsigned(1299669553,32),
    to_unsigned(1299833447,32),
    to_unsigned(1299997330,32),
    to_unsigned(1300161201,32),
    to_unsigned(1300325059,32),
    to_unsigned(1300488906,32),
    to_unsigned(1300652741,32),
    to_unsigned(1300816564,32),
    to_unsigned(1300980375,32),
    to_unsigned(1301144174,32),
    to_unsigned(1301307961,32),
    to_unsigned(1301471736,32),
    to_unsigned(1301635499,32),
    to_unsigned(1301799250,32),
    to_unsigned(1301962990,32),
    to_unsigned(1302126717,32),
    to_unsigned(1302290432,32),
    to_unsigned(1302454135,32),
    to_unsigned(1302617827,32),
    to_unsigned(1302781506,32),
    to_unsigned(1302945173,32),
    to_unsigned(1303108829,32),
    to_unsigned(1303272472,32),
    to_unsigned(1303436104,32),
    to_unsigned(1303599723,32),
    to_unsigned(1303763331,32),
    to_unsigned(1303926926,32),
    to_unsigned(1304090510,32),
    to_unsigned(1304254081,32),
    to_unsigned(1304417641,32),
    to_unsigned(1304581188,32),
    to_unsigned(1304744724,32),
    to_unsigned(1304908247,32),
    to_unsigned(1305071759,32),
    to_unsigned(1305235258,32),
    to_unsigned(1305398746,32),
    to_unsigned(1305562221,32),
    to_unsigned(1305725685,32),
    to_unsigned(1305889137,32),
    to_unsigned(1306052576,32),
    to_unsigned(1306216004,32),
    to_unsigned(1306379419,32),
    to_unsigned(1306542823,32),
    to_unsigned(1306706214,32),
    to_unsigned(1306869594,32),
    to_unsigned(1307032961,32),
    to_unsigned(1307196317,32),
    to_unsigned(1307359660,32),
    to_unsigned(1307522992,32),
    to_unsigned(1307686311,32),
    to_unsigned(1307849619,32),
    to_unsigned(1308012914,32),
    to_unsigned(1308176197,32),
    to_unsigned(1308339469,32),
    to_unsigned(1308502728,32),
    to_unsigned(1308665975,32),
    to_unsigned(1308829211,32),
    to_unsigned(1308992434,32),
    to_unsigned(1309155645,32),
    to_unsigned(1309318844,32),
    to_unsigned(1309482031,32),
    to_unsigned(1309645206,32),
    to_unsigned(1309808369,32),
    to_unsigned(1309971520,32),
    to_unsigned(1310134659,32),
    to_unsigned(1310297786,32),
    to_unsigned(1310460901,32),
    to_unsigned(1310624004,32),
    to_unsigned(1310787095,32),
    to_unsigned(1310950174,32),
    to_unsigned(1311113240,32),
    to_unsigned(1311276295,32),
    to_unsigned(1311439338,32),
    to_unsigned(1311602368,32),
    to_unsigned(1311765387,32),
    to_unsigned(1311928393,32),
    to_unsigned(1312091387,32),
    to_unsigned(1312254370,32),
    to_unsigned(1312417340,32),
    to_unsigned(1312580298,32),
    to_unsigned(1312743244,32),
    to_unsigned(1312906178,32),
    to_unsigned(1313069100,32),
    to_unsigned(1313232010,32),
    to_unsigned(1313394908,32),
    to_unsigned(1313557794,32),
    to_unsigned(1313720668,32),
    to_unsigned(1313883529,32),
    to_unsigned(1314046379,32),
    to_unsigned(1314209216,32),
    to_unsigned(1314372042,32),
    to_unsigned(1314534855,32),
    to_unsigned(1314697656,32),
    to_unsigned(1314860445,32),
    to_unsigned(1315023222,32),
    to_unsigned(1315185987,32),
    to_unsigned(1315348740,32),
    to_unsigned(1315511481,32),
    to_unsigned(1315674210,32),
    to_unsigned(1315836926,32),
    to_unsigned(1315999631,32),
    to_unsigned(1316162323,32),
    to_unsigned(1316325003,32),
    to_unsigned(1316487672,32),
    to_unsigned(1316650328,32),
    to_unsigned(1316812972,32),
    to_unsigned(1316975604,32),
    to_unsigned(1317138223,32),
    to_unsigned(1317300831,32),
    to_unsigned(1317463427,32),
    to_unsigned(1317626010,32),
    to_unsigned(1317788582,32),
    to_unsigned(1317951141,32),
    to_unsigned(1318113688,32),
    to_unsigned(1318276223,32),
    to_unsigned(1318438746,32),
    to_unsigned(1318601257,32),
    to_unsigned(1318763755,32),
    to_unsigned(1318926242,32),
    to_unsigned(1319088716,32),
    to_unsigned(1319251179,32),
    to_unsigned(1319413629,32),
    to_unsigned(1319576067,32),
    to_unsigned(1319738493,32),
    to_unsigned(1319900907,32),
    to_unsigned(1320063308,32),
    to_unsigned(1320225698,32),
    to_unsigned(1320388075,32),
    to_unsigned(1320550440,32),
    to_unsigned(1320712793,32),
    to_unsigned(1320875134,32),
    to_unsigned(1321037463,32),
    to_unsigned(1321199780,32),
    to_unsigned(1321362084,32),
    to_unsigned(1321524377,32),
    to_unsigned(1321686657,32),
    to_unsigned(1321848925,32),
    to_unsigned(1322011181,32),
    to_unsigned(1322173425,32),
    to_unsigned(1322335657,32),
    to_unsigned(1322497876,32),
    to_unsigned(1322660083,32),
    to_unsigned(1322822279,32),
    to_unsigned(1322984462,32),
    to_unsigned(1323146632,32),
    to_unsigned(1323308791,32),
    to_unsigned(1323470938,32),
    to_unsigned(1323633072,32),
    to_unsigned(1323795194,32),
    to_unsigned(1323957304,32),
    to_unsigned(1324119402,32),
    to_unsigned(1324281488,32),
    to_unsigned(1324443561,32),
    to_unsigned(1324605623,32),
    to_unsigned(1324767672,32),
    to_unsigned(1324929709,32),
    to_unsigned(1325091734,32),
    to_unsigned(1325253746,32),
    to_unsigned(1325415747,32),
    to_unsigned(1325577735,32),
    to_unsigned(1325739711,32),
    to_unsigned(1325901675,32),
    to_unsigned(1326063627,32),
    to_unsigned(1326225566,32),
    to_unsigned(1326387493,32),
    to_unsigned(1326549409,32),
    to_unsigned(1326711311,32),
    to_unsigned(1326873202,32),
    to_unsigned(1327035081,32),
    to_unsigned(1327196947,32),
    to_unsigned(1327358801,32),
    to_unsigned(1327520643,32),
    to_unsigned(1327682473,32),
    to_unsigned(1327844291,32),
    to_unsigned(1328006096,32),
    to_unsigned(1328167889,32),
    to_unsigned(1328329670,32),
    to_unsigned(1328491439,32),
    to_unsigned(1328653195,32),
    to_unsigned(1328814939,32),
    to_unsigned(1328976672,32),
    to_unsigned(1329138391,32),
    to_unsigned(1329300099,32),
    to_unsigned(1329461794,32),
    to_unsigned(1329623478,32),
    to_unsigned(1329785149,32),
    to_unsigned(1329946807,32),
    to_unsigned(1330108454,32),
    to_unsigned(1330270088,32),
    to_unsigned(1330431710,32),
    to_unsigned(1330593320,32),
    to_unsigned(1330754918,32),
    to_unsigned(1330916503,32),
    to_unsigned(1331078076,32),
    to_unsigned(1331239637,32),
    to_unsigned(1331401186,32),
    to_unsigned(1331562722,32),
    to_unsigned(1331724247,32),
    to_unsigned(1331885759,32),
    to_unsigned(1332047258,32),
    to_unsigned(1332208746,32),
    to_unsigned(1332370221,32),
    to_unsigned(1332531684,32),
    to_unsigned(1332693135,32),
    to_unsigned(1332854573,32),
    to_unsigned(1333016000,32),
    to_unsigned(1333177414,32),
    to_unsigned(1333338815,32),
    to_unsigned(1333500205,32),
    to_unsigned(1333661582,32),
    to_unsigned(1333822947,32),
    to_unsigned(1333984300,32),
    to_unsigned(1334145640,32),
    to_unsigned(1334306968,32),
    to_unsigned(1334468284,32),
    to_unsigned(1334629588,32),
    to_unsigned(1334790879,32),
    to_unsigned(1334952158,32),
    to_unsigned(1335113425,32),
    to_unsigned(1335274680,32),
    to_unsigned(1335435922,32),
    to_unsigned(1335597152,32),
    to_unsigned(1335758370,32),
    to_unsigned(1335919575,32),
    to_unsigned(1336080768,32),
    to_unsigned(1336241949,32),
    to_unsigned(1336403118,32),
    to_unsigned(1336564274,32),
    to_unsigned(1336725418,32),
    to_unsigned(1336886550,32),
    to_unsigned(1337047670,32),
    to_unsigned(1337208777,32),
    to_unsigned(1337369872,32),
    to_unsigned(1337530954,32),
    to_unsigned(1337692025,32),
    to_unsigned(1337853083,32),
    to_unsigned(1338014128,32),
    to_unsigned(1338175162,32),
    to_unsigned(1338336183,32),
    to_unsigned(1338497192,32),
    to_unsigned(1338658188,32),
    to_unsigned(1338819172,32),
    to_unsigned(1338980144,32),
    to_unsigned(1339141104,32),
    to_unsigned(1339302051,32),
    to_unsigned(1339462986,32),
    to_unsigned(1339623909,32),
    to_unsigned(1339784819,32),
    to_unsigned(1339945717,32),
    to_unsigned(1340106603,32),
    to_unsigned(1340267476,32),
    to_unsigned(1340428337,32),
    to_unsigned(1340589186,32),
    to_unsigned(1340750023,32),
    to_unsigned(1340910847,32),
    to_unsigned(1341071658,32),
    to_unsigned(1341232458,32),
    to_unsigned(1341393245,32),
    to_unsigned(1341554020,32),
    to_unsigned(1341714782,32),
    to_unsigned(1341875532,32),
    to_unsigned(1342036270,32),
    to_unsigned(1342196996,32),
    to_unsigned(1342357709,32),
    to_unsigned(1342518410,32),
    to_unsigned(1342679098,32),
    to_unsigned(1342839774,32),
    to_unsigned(1343000438,32),
    to_unsigned(1343161089,32),
    to_unsigned(1343321728,32),
    to_unsigned(1343482355,32),
    to_unsigned(1343642970,32),
    to_unsigned(1343803572,32),
    to_unsigned(1343964161,32),
    to_unsigned(1344124739,32),
    to_unsigned(1344285304,32),
    to_unsigned(1344445856,32),
    to_unsigned(1344606396,32),
    to_unsigned(1344766924,32),
    to_unsigned(1344927440,32),
    to_unsigned(1345087943,32),
    to_unsigned(1345248434,32),
    to_unsigned(1345408912,32),
    to_unsigned(1345569378,32),
    to_unsigned(1345729832,32),
    to_unsigned(1345890273,32),
    to_unsigned(1346050702,32),
    to_unsigned(1346211119,32),
    to_unsigned(1346371523,32),
    to_unsigned(1346531915,32),
    to_unsigned(1346692295,32),
    to_unsigned(1346852662,32),
    to_unsigned(1347013016,32),
    to_unsigned(1347173359,32),
    to_unsigned(1347333689,32),
    to_unsigned(1347494006,32),
    to_unsigned(1347654311,32),
    to_unsigned(1347814604,32),
    to_unsigned(1347974885,32),
    to_unsigned(1348135153,32),
    to_unsigned(1348295408,32),
    to_unsigned(1348455651,32),
    to_unsigned(1348615882,32),
    to_unsigned(1348776101,32),
    to_unsigned(1348936307,32),
    to_unsigned(1349096500,32),
    to_unsigned(1349256682,32),
    to_unsigned(1349416850,32),
    to_unsigned(1349577007,32),
    to_unsigned(1349737151,32),
    to_unsigned(1349897282,32),
    to_unsigned(1350057402,32),
    to_unsigned(1350217508,32),
    to_unsigned(1350377603,32),
    to_unsigned(1350537685,32),
    to_unsigned(1350697754,32),
    to_unsigned(1350857812,32),
    to_unsigned(1351017856,32),
    to_unsigned(1351177889,32),
    to_unsigned(1351337908,32),
    to_unsigned(1351497916,32),
    to_unsigned(1351657911,32),
    to_unsigned(1351817894,32),
    to_unsigned(1351977864,32),
    to_unsigned(1352137822,32),
    to_unsigned(1352297767,32),
    to_unsigned(1352457700,32),
    to_unsigned(1352617620,32),
    to_unsigned(1352777528,32),
    to_unsigned(1352937424,32),
    to_unsigned(1353097307,32),
    to_unsigned(1353257178,32),
    to_unsigned(1353417036,32),
    to_unsigned(1353576882,32),
    to_unsigned(1353736716,32),
    to_unsigned(1353896536,32),
    to_unsigned(1354056345,32),
    to_unsigned(1354216141,32),
    to_unsigned(1354375925,32),
    to_unsigned(1354535696,32),
    to_unsigned(1354695455,32),
    to_unsigned(1354855201,32),
    to_unsigned(1355014935,32),
    to_unsigned(1355174656,32),
    to_unsigned(1355334365,32),
    to_unsigned(1355494062,32),
    to_unsigned(1355653746,32),
    to_unsigned(1355813417,32),
    to_unsigned(1355973076,32),
    to_unsigned(1356132723,32),
    to_unsigned(1356292357,32),
    to_unsigned(1356451979,32),
    to_unsigned(1356611588,32),
    to_unsigned(1356771185,32),
    to_unsigned(1356930769,32),
    to_unsigned(1357090341,32),
    to_unsigned(1357249900,32),
    to_unsigned(1357409447,32),
    to_unsigned(1357568981,32),
    to_unsigned(1357728503,32),
    to_unsigned(1357888013,32),
    to_unsigned(1358047510,32),
    to_unsigned(1358206994,32),
    to_unsigned(1358366466,32),
    to_unsigned(1358525925,32),
    to_unsigned(1358685372,32),
    to_unsigned(1358844807,32),
    to_unsigned(1359004229,32),
    to_unsigned(1359163638,32),
    to_unsigned(1359323036,32),
    to_unsigned(1359482420,32),
    to_unsigned(1359641792,32),
    to_unsigned(1359801152,32),
    to_unsigned(1359960499,32),
    to_unsigned(1360119833,32),
    to_unsigned(1360279155,32),
    to_unsigned(1360438465,32),
    to_unsigned(1360597762,32),
    to_unsigned(1360757046,32),
    to_unsigned(1360916318,32),
    to_unsigned(1361075578,32),
    to_unsigned(1361234825,32),
    to_unsigned(1361394059,32),
    to_unsigned(1361553281,32),
    to_unsigned(1361712491,32),
    to_unsigned(1361871688,32),
    to_unsigned(1362030872,32),
    to_unsigned(1362190044,32),
    to_unsigned(1362349204,32),
    to_unsigned(1362508350,32),
    to_unsigned(1362667485,32),
    to_unsigned(1362826607,32),
    to_unsigned(1362985716,32),
    to_unsigned(1363144813,32),
    to_unsigned(1363303897,32),
    to_unsigned(1363462968,32),
    to_unsigned(1363622028,32),
    to_unsigned(1363781074,32),
    to_unsigned(1363940108,32),
    to_unsigned(1364099130,32),
    to_unsigned(1364258139,32),
    to_unsigned(1364417135,32),
    to_unsigned(1364576119,32),
    to_unsigned(1364735091,32),
    to_unsigned(1364894050,32),
    to_unsigned(1365052996,32),
    to_unsigned(1365211930,32),
    to_unsigned(1365370851,32),
    to_unsigned(1365529760,32),
    to_unsigned(1365688656,32),
    to_unsigned(1365847539,32),
    to_unsigned(1366006410,32),
    to_unsigned(1366165269,32),
    to_unsigned(1366324115,32),
    to_unsigned(1366482948,32),
    to_unsigned(1366641769,32),
    to_unsigned(1366800577,32),
    to_unsigned(1366959373,32),
    to_unsigned(1367118156,32),
    to_unsigned(1367276926,32),
    to_unsigned(1367435684,32),
    to_unsigned(1367594429,32),
    to_unsigned(1367753162,32),
    to_unsigned(1367911882,32),
    to_unsigned(1368070590,32),
    to_unsigned(1368229285,32),
    to_unsigned(1368387968,32),
    to_unsigned(1368546638,32),
    to_unsigned(1368705295,32),
    to_unsigned(1368863940,32),
    to_unsigned(1369022572,32),
    to_unsigned(1369181192,32),
    to_unsigned(1369339799,32),
    to_unsigned(1369498393,32),
    to_unsigned(1369656975,32),
    to_unsigned(1369815544,32),
    to_unsigned(1369974101,32),
    to_unsigned(1370132645,32),
    to_unsigned(1370291176,32),
    to_unsigned(1370449695,32),
    to_unsigned(1370608201,32),
    to_unsigned(1370766695,32),
    to_unsigned(1370925176,32),
    to_unsigned(1371083645,32),
    to_unsigned(1371242101,32),
    to_unsigned(1371400544,32),
    to_unsigned(1371558975,32),
    to_unsigned(1371717393,32),
    to_unsigned(1371875798,32),
    to_unsigned(1372034191,32),
    to_unsigned(1372192571,32),
    to_unsigned(1372350939,32),
    to_unsigned(1372509294,32),
    to_unsigned(1372667636,32),
    to_unsigned(1372825966,32),
    to_unsigned(1372984283,32),
    to_unsigned(1373142588,32),
    to_unsigned(1373300880,32),
    to_unsigned(1373459159,32),
    to_unsigned(1373617425,32),
    to_unsigned(1373775680,32),
    to_unsigned(1373933921,32),
    to_unsigned(1374092150,32),
    to_unsigned(1374250366,32),
    to_unsigned(1374408569,32),
    to_unsigned(1374566760,32),
    to_unsigned(1374724939,32),
    to_unsigned(1374883104,32),
    to_unsigned(1375041257,32),
    to_unsigned(1375199397,32),
    to_unsigned(1375357525,32),
    to_unsigned(1375515640,32),
    to_unsigned(1375673743,32),
    to_unsigned(1375831832,32),
    to_unsigned(1375989910,32),
    to_unsigned(1376147974,32),
    to_unsigned(1376306026,32),
    to_unsigned(1376464065,32),
    to_unsigned(1376622092,32),
    to_unsigned(1376780105,32),
    to_unsigned(1376938107,32),
    to_unsigned(1377096095,32),
    to_unsigned(1377254071,32),
    to_unsigned(1377412034,32),
    to_unsigned(1377569985,32),
    to_unsigned(1377727923,32),
    to_unsigned(1377885848,32),
    to_unsigned(1378043761,32),
    to_unsigned(1378201661,32),
    to_unsigned(1378359548,32),
    to_unsigned(1378517422,32),
    to_unsigned(1378675284,32),
    to_unsigned(1378833134,32),
    to_unsigned(1378990970,32),
    to_unsigned(1379148794,32),
    to_unsigned(1379306605,32),
    to_unsigned(1379464404,32),
    to_unsigned(1379622190,32),
    to_unsigned(1379779963,32),
    to_unsigned(1379937723,32),
    to_unsigned(1380095471,32),
    to_unsigned(1380253206,32),
    to_unsigned(1380410929,32),
    to_unsigned(1380568638,32),
    to_unsigned(1380726335,32),
    to_unsigned(1380884020,32),
    to_unsigned(1381041691,32),
    to_unsigned(1381199350,32),
    to_unsigned(1381356997,32),
    to_unsigned(1381514630,32),
    to_unsigned(1381672251,32),
    to_unsigned(1381829859,32),
    to_unsigned(1381987455,32),
    to_unsigned(1382145038,32),
    to_unsigned(1382302608,32),
    to_unsigned(1382460165,32),
    to_unsigned(1382617710,32),
    to_unsigned(1382775242,32),
    to_unsigned(1382932761,32),
    to_unsigned(1383090268,32),
    to_unsigned(1383247761,32),
    to_unsigned(1383405242,32),
    to_unsigned(1383562711,32),
    to_unsigned(1383720167,32),
    to_unsigned(1383877609,32),
    to_unsigned(1384035040,32),
    to_unsigned(1384192457,32),
    to_unsigned(1384349862,32),
    to_unsigned(1384507254,32),
    to_unsigned(1384664633,32),
    to_unsigned(1384822000,32),
    to_unsigned(1384979354,32),
    to_unsigned(1385136695,32),
    to_unsigned(1385294023,32),
    to_unsigned(1385451339,32),
    to_unsigned(1385608642,32),
    to_unsigned(1385765932,32),
    to_unsigned(1385923210,32),
    to_unsigned(1386080475,32),
    to_unsigned(1386237727,32),
    to_unsigned(1386394966,32),
    to_unsigned(1386552192,32),
    to_unsigned(1386709406,32),
    to_unsigned(1386866607,32),
    to_unsigned(1387023795,32),
    to_unsigned(1387180971,32),
    to_unsigned(1387338134,32),
    to_unsigned(1387495284,32),
    to_unsigned(1387652421,32),
    to_unsigned(1387809545,32),
    to_unsigned(1387966657,32),
    to_unsigned(1388123756,32),
    to_unsigned(1388280842,32),
    to_unsigned(1388437916,32),
    to_unsigned(1388594977,32),
    to_unsigned(1388752025,32),
    to_unsigned(1388909060,32),
    to_unsigned(1389066082,32),
    to_unsigned(1389223092,32),
    to_unsigned(1389380089,32),
    to_unsigned(1389537073,32),
    to_unsigned(1389694044,32),
    to_unsigned(1389851003,32),
    to_unsigned(1390007949,32),
    to_unsigned(1390164882,32),
    to_unsigned(1390321802,32),
    to_unsigned(1390478709,32),
    to_unsigned(1390635604,32),
    to_unsigned(1390792486,32),
    to_unsigned(1390949355,32),
    to_unsigned(1391106211,32),
    to_unsigned(1391263055,32),
    to_unsigned(1391419886,32),
    to_unsigned(1391576704,32),
    to_unsigned(1391733509,32),
    to_unsigned(1391890301,32),
    to_unsigned(1392047081,32),
    to_unsigned(1392203847,32),
    to_unsigned(1392360601,32),
    to_unsigned(1392517343,32),
    to_unsigned(1392674071,32),
    to_unsigned(1392830787,32),
    to_unsigned(1392987489,32),
    to_unsigned(1393144179,32),
    to_unsigned(1393300857,32),
    to_unsigned(1393457521,32),
    to_unsigned(1393614173,32),
    to_unsigned(1393770811,32),
    to_unsigned(1393927437,32),
    to_unsigned(1394084050,32),
    to_unsigned(1394240651,32),
    to_unsigned(1394397238,32),
    to_unsigned(1394553813,32),
    to_unsigned(1394710375,32),
    to_unsigned(1394866924,32),
    to_unsigned(1395023460,32),
    to_unsigned(1395179983,32),
    to_unsigned(1395336494,32),
    to_unsigned(1395492992,32),
    to_unsigned(1395649477,32),
    to_unsigned(1395805949,32),
    to_unsigned(1395962408,32),
    to_unsigned(1396118854,32),
    to_unsigned(1396275288,32),
    to_unsigned(1396431709,32),
    to_unsigned(1396588117,32),
    to_unsigned(1396744512,32),
    to_unsigned(1396900894,32),
    to_unsigned(1397057263,32),
    to_unsigned(1397213620,32),
    to_unsigned(1397369964,32),
    to_unsigned(1397526295,32),
    to_unsigned(1397682613,32),
    to_unsigned(1397838918,32),
    to_unsigned(1397995210,32),
    to_unsigned(1398151490,32),
    to_unsigned(1398307756,32),
    to_unsigned(1398464010,32),
    to_unsigned(1398620251,32),
    to_unsigned(1398776479,32),
    to_unsigned(1398932694,32),
    to_unsigned(1399088897,32),
    to_unsigned(1399245086,32),
    to_unsigned(1399401263,32),
    to_unsigned(1399557427,32),
    to_unsigned(1399713578,32),
    to_unsigned(1399869716,32),
    to_unsigned(1400025841,32),
    to_unsigned(1400181953,32),
    to_unsigned(1400338053,32),
    to_unsigned(1400494139,32),
    to_unsigned(1400650213,32),
    to_unsigned(1400806274,32),
    to_unsigned(1400962322,32),
    to_unsigned(1401118357,32),
    to_unsigned(1401274379,32),
    to_unsigned(1401430388,32),
    to_unsigned(1401586385,32),
    to_unsigned(1401742368,32),
    to_unsigned(1401898339,32),
    to_unsigned(1402054297,32),
    to_unsigned(1402210242,32),
    to_unsigned(1402366174,32),
    to_unsigned(1402522093,32),
    to_unsigned(1402677999,32),
    to_unsigned(1402833892,32),
    to_unsigned(1402989773,32),
    to_unsigned(1403145640,32),
    to_unsigned(1403301495,32),
    to_unsigned(1403457337,32),
    to_unsigned(1403613165,32),
    to_unsigned(1403768981,32),
    to_unsigned(1403924784,32),
    to_unsigned(1404080575,32),
    to_unsigned(1404236352,32),
    to_unsigned(1404392116,32),
    to_unsigned(1404547867,32),
    to_unsigned(1404703606,32),
    to_unsigned(1404859332,32),
    to_unsigned(1405015044,32),
    to_unsigned(1405170744,32),
    to_unsigned(1405326431,32),
    to_unsigned(1405482105,32),
    to_unsigned(1405637766,32),
    to_unsigned(1405793414,32),
    to_unsigned(1405949049,32),
    to_unsigned(1406104671,32),
    to_unsigned(1406260281,32),
    to_unsigned(1406415877,32),
    to_unsigned(1406571460,32),
    to_unsigned(1406727031,32),
    to_unsigned(1406882589,32),
    to_unsigned(1407038133,32),
    to_unsigned(1407193665,32),
    to_unsigned(1407349184,32),
    to_unsigned(1407504690,32),
    to_unsigned(1407660183,32),
    to_unsigned(1407815663,32),
    to_unsigned(1407971130,32),
    to_unsigned(1408126584,32),
    to_unsigned(1408282025,32),
    to_unsigned(1408437453,32),
    to_unsigned(1408592868,32),
    to_unsigned(1408748271,32),
    to_unsigned(1408903660,32),
    to_unsigned(1409059036,32),
    to_unsigned(1409214400,32),
    to_unsigned(1409369750,32),
    to_unsigned(1409525088,32),
    to_unsigned(1409680413,32),
    to_unsigned(1409835724,32),
    to_unsigned(1409991023,32),
    to_unsigned(1410146309,32),
    to_unsigned(1410301582,32),
    to_unsigned(1410456841,32),
    to_unsigned(1410612088,32),
    to_unsigned(1410767322,32),
    to_unsigned(1410922543,32),
    to_unsigned(1411077751,32),
    to_unsigned(1411232946,32),
    to_unsigned(1411388128,32),
    to_unsigned(1411543297,32),
    to_unsigned(1411698453,32),
    to_unsigned(1411853596,32),
    to_unsigned(1412008726,32),
    to_unsigned(1412163843,32),
    to_unsigned(1412318947,32),
    to_unsigned(1412474039,32),
    to_unsigned(1412629117,32),
    to_unsigned(1412784182,32),
    to_unsigned(1412939234,32),
    to_unsigned(1413094273,32),
    to_unsigned(1413249300,32),
    to_unsigned(1413404313,32),
    to_unsigned(1413559313,32),
    to_unsigned(1413714300,32),
    to_unsigned(1413869275,32),
    to_unsigned(1414024236,32),
    to_unsigned(1414179184,32),
    to_unsigned(1414334119,32),
    to_unsigned(1414489042,32),
    to_unsigned(1414643951,32),
    to_unsigned(1414798847,32),
    to_unsigned(1414953730,32),
    to_unsigned(1415108601,32),
    to_unsigned(1415263458,32),
    to_unsigned(1415418302,32),
    to_unsigned(1415573133,32),
    to_unsigned(1415727952,32),
    to_unsigned(1415882757,32),
    to_unsigned(1416037549,32),
    to_unsigned(1416192328,32),
    to_unsigned(1416347094,32),
    to_unsigned(1416501847,32),
    to_unsigned(1416656588,32),
    to_unsigned(1416811315,32),
    to_unsigned(1416966029,32),
    to_unsigned(1417120730,32),
    to_unsigned(1417275418,32),
    to_unsigned(1417430093,32),
    to_unsigned(1417584755,32),
    to_unsigned(1417739404,32),
    to_unsigned(1417894040,32),
    to_unsigned(1418048662,32),
    to_unsigned(1418203272,32),
    to_unsigned(1418357869,32),
    to_unsigned(1418512453,32),
    to_unsigned(1418667024,32),
    to_unsigned(1418821581,32),
    to_unsigned(1418976126,32),
    to_unsigned(1419130657,32),
    to_unsigned(1419285176,32),
    to_unsigned(1419439682,32),
    to_unsigned(1419594174,32),
    to_unsigned(1419748653,32),
    to_unsigned(1419903120,32),
    to_unsigned(1420057573,32),
    to_unsigned(1420212013,32),
    to_unsigned(1420366441,32),
    to_unsigned(1420520855,32),
    to_unsigned(1420675256,32),
    to_unsigned(1420829644,32),
    to_unsigned(1420984019,32),
    to_unsigned(1421138381,32),
    to_unsigned(1421292730,32),
    to_unsigned(1421447065,32),
    to_unsigned(1421601388,32),
    to_unsigned(1421755698,32),
    to_unsigned(1421909994,32),
    to_unsigned(1422064278,32),
    to_unsigned(1422218548,32),
    to_unsigned(1422372806,32),
    to_unsigned(1422527050,32),
    to_unsigned(1422681281,32),
    to_unsigned(1422835499,32),
    to_unsigned(1422989704,32),
    to_unsigned(1423143896,32),
    to_unsigned(1423298075,32),
    to_unsigned(1423452241,32),
    to_unsigned(1423606394,32),
    to_unsigned(1423760533,32),
    to_unsigned(1423914660,32),
    to_unsigned(1424068773,32),
    to_unsigned(1424222874,32),
    to_unsigned(1424376961,32),
    to_unsigned(1424531035,32),
    to_unsigned(1424685096,32),
    to_unsigned(1424839144,32),
    to_unsigned(1424993179,32),
    to_unsigned(1425147201,32),
    to_unsigned(1425301210,32),
    to_unsigned(1425455206,32),
    to_unsigned(1425609188,32),
    to_unsigned(1425763157,32),
    to_unsigned(1425917114,32),
    to_unsigned(1426071057,32),
    to_unsigned(1426224987,32),
    to_unsigned(1426378904,32),
    to_unsigned(1426532808,32),
    to_unsigned(1426686699,32),
    to_unsigned(1426840576,32),
    to_unsigned(1426994441,32),
    to_unsigned(1427148292,32),
    to_unsigned(1427302130,32),
    to_unsigned(1427455956,32),
    to_unsigned(1427609768,32),
    to_unsigned(1427763567,32),
    to_unsigned(1427917352,32),
    to_unsigned(1428071125,32),
    to_unsigned(1428224885,32),
    to_unsigned(1428378631,32),
    to_unsigned(1428532364,32),
    to_unsigned(1428686085,32),
    to_unsigned(1428839792,32),
    to_unsigned(1428993486,32),
    to_unsigned(1429147166,32),
    to_unsigned(1429300834,32),
    to_unsigned(1429454488,32),
    to_unsigned(1429608130,32),
    to_unsigned(1429761758,32),
    to_unsigned(1429915373,32),
    to_unsigned(1430068975,32),
    to_unsigned(1430222564,32),
    to_unsigned(1430376139,32),
    to_unsigned(1430529702,32),
    to_unsigned(1430683251,32),
    to_unsigned(1430836787,32),
    to_unsigned(1430990310,32),
    to_unsigned(1431143820,32),
    to_unsigned(1431297317,32),
    to_unsigned(1431450801,32),
    to_unsigned(1431604271,32),
    to_unsigned(1431757728,32),
    to_unsigned(1431911172,32),
    to_unsigned(1432064603,32),
    to_unsigned(1432218021,32),
    to_unsigned(1432371426,32),
    to_unsigned(1432524817,32),
    to_unsigned(1432678195,32),
    to_unsigned(1432831561,32),
    to_unsigned(1432984912,32),
    to_unsigned(1433138251,32),
    to_unsigned(1433291577,32),
    to_unsigned(1433444889,32),
    to_unsigned(1433598188,32),
    to_unsigned(1433751475,32),
    to_unsigned(1433904747,32),
    to_unsigned(1434058007,32),
    to_unsigned(1434211254,32),
    to_unsigned(1434364487,32),
    to_unsigned(1434517707,32),
    to_unsigned(1434670914,32),
    to_unsigned(1434824108,32),
    to_unsigned(1434977288,32),
    to_unsigned(1435130456,32),
    to_unsigned(1435283610,32),
    to_unsigned(1435436751,32),
    to_unsigned(1435589879,32),
    to_unsigned(1435742994,32),
    to_unsigned(1435896095,32),
    to_unsigned(1436049183,32),
    to_unsigned(1436202258,32),
    to_unsigned(1436355320,32),
    to_unsigned(1436508369,32),
    to_unsigned(1436661404,32),
    to_unsigned(1436814426,32),
    to_unsigned(1436967435,32),
    to_unsigned(1437120431,32),
    to_unsigned(1437273414,32),
    to_unsigned(1437426383,32),
    to_unsigned(1437579339,32),
    to_unsigned(1437732282,32),
    to_unsigned(1437885212,32),
    to_unsigned(1438038128,32),
    to_unsigned(1438191032,32),
    to_unsigned(1438343922,32),
    to_unsigned(1438496799,32),
    to_unsigned(1438649662,32),
    to_unsigned(1438802513,32),
    to_unsigned(1438955350,32),
    to_unsigned(1439108174,32),
    to_unsigned(1439260985,32),
    to_unsigned(1439413782,32),
    to_unsigned(1439566566,32),
    to_unsigned(1439719338,32),
    to_unsigned(1439872095,32),
    to_unsigned(1440024840,32),
    to_unsigned(1440177571,32),
    to_unsigned(1440330289,32),
    to_unsigned(1440482994,32),
    to_unsigned(1440635686,32),
    to_unsigned(1440788364,32),
    to_unsigned(1440941029,32),
    to_unsigned(1441093681,32),
    to_unsigned(1441246320,32),
    to_unsigned(1441398945,32),
    to_unsigned(1441551557,32),
    to_unsigned(1441704156,32),
    to_unsigned(1441856742,32),
    to_unsigned(1442009314,32),
    to_unsigned(1442161874,32),
    to_unsigned(1442314419,32),
    to_unsigned(1442466952,32),
    to_unsigned(1442619471,32),
    to_unsigned(1442771978,32),
    to_unsigned(1442924470,32),
    to_unsigned(1443076950,32),
    to_unsigned(1443229416,32),
    to_unsigned(1443381869,32),
    to_unsigned(1443534309,32),
    to_unsigned(1443686736,32),
    to_unsigned(1443839149,32),
    to_unsigned(1443991549,32),
    to_unsigned(1444143936,32),
    to_unsigned(1444296309,32),
    to_unsigned(1444448669,32),
    to_unsigned(1444601016,32),
    to_unsigned(1444753350,32),
    to_unsigned(1444905670,32),
    to_unsigned(1445057977,32),
    to_unsigned(1445210271,32),
    to_unsigned(1445362551,32),
    to_unsigned(1445514818,32),
    to_unsigned(1445667072,32),
    to_unsigned(1445819313,32),
    to_unsigned(1445971540,32),
    to_unsigned(1446123754,32),
    to_unsigned(1446275955,32),
    to_unsigned(1446428142,32),
    to_unsigned(1446580317,32),
    to_unsigned(1446732477,32),
    to_unsigned(1446884625,32),
    to_unsigned(1447036759,32),
    to_unsigned(1447188880,32),
    to_unsigned(1447340988,32),
    to_unsigned(1447493082,32),
    to_unsigned(1447645163,32),
    to_unsigned(1447797231,32),
    to_unsigned(1447949285,32),
    to_unsigned(1448101326,32),
    to_unsigned(1448253354,32),
    to_unsigned(1448405369,32),
    to_unsigned(1448557370,32),
    to_unsigned(1448709358,32),
    to_unsigned(1448861332,32),
    to_unsigned(1449013294,32),
    to_unsigned(1449165241,32),
    to_unsigned(1449317176,32),
    to_unsigned(1449469097,32),
    to_unsigned(1449621005,32),
    to_unsigned(1449772900,32),
    to_unsigned(1449924781,32),
    to_unsigned(1450076649,32),
    to_unsigned(1450228504,32),
    to_unsigned(1450380345,32),
    to_unsigned(1450532173,32),
    to_unsigned(1450683988,32),
    to_unsigned(1450835789,32),
    to_unsigned(1450987577,32),
    to_unsigned(1451139352,32),
    to_unsigned(1451291113,32),
    to_unsigned(1451442861,32),
    to_unsigned(1451594596,32),
    to_unsigned(1451746317,32),
    to_unsigned(1451898025,32),
    to_unsigned(1452049719,32),
    to_unsigned(1452201401,32),
    to_unsigned(1452353069,32),
    to_unsigned(1452504723,32),
    to_unsigned(1452656364,32),
    to_unsigned(1452807992,32),
    to_unsigned(1452959607,32),
    to_unsigned(1453111208,32),
    to_unsigned(1453262795,32),
    to_unsigned(1453414370,32),
    to_unsigned(1453565931,32),
    to_unsigned(1453717479,32),
    to_unsigned(1453869013,32),
    to_unsigned(1454020534,32),
    to_unsigned(1454172042,32),
    to_unsigned(1454323536,32),
    to_unsigned(1454475017,32),
    to_unsigned(1454626484,32),
    to_unsigned(1454777938,32),
    to_unsigned(1454929379,32),
    to_unsigned(1455080806,32),
    to_unsigned(1455232220,32),
    to_unsigned(1455383621,32),
    to_unsigned(1455535008,32),
    to_unsigned(1455686382,32),
    to_unsigned(1455837743,32),
    to_unsigned(1455989090,32),
    to_unsigned(1456140424,32),
    to_unsigned(1456291744,32),
    to_unsigned(1456443051,32),
    to_unsigned(1456594344,32),
    to_unsigned(1456745625,32),
    to_unsigned(1456896891,32),
    to_unsigned(1457048145,32),
    to_unsigned(1457199385,32),
    to_unsigned(1457350611,32),
    to_unsigned(1457501825,32),
    to_unsigned(1457653024,32),
    to_unsigned(1457804211,32),
    to_unsigned(1457955384,32),
    to_unsigned(1458106543,32),
    to_unsigned(1458257690,32),
    to_unsigned(1458408823,32),
    to_unsigned(1458559942,32),
    to_unsigned(1458711048,32),
    to_unsigned(1458862141,32),
    to_unsigned(1459013220,32),
    to_unsigned(1459164286,32),
    to_unsigned(1459315338,32),
    to_unsigned(1459466377,32),
    to_unsigned(1459617402,32),
    to_unsigned(1459768414,32),
    to_unsigned(1459919413,32),
    to_unsigned(1460070398,32),
    to_unsigned(1460221370,32),
    to_unsigned(1460372329,32),
    to_unsigned(1460523274,32),
    to_unsigned(1460674205,32),
    to_unsigned(1460825124,32),
    to_unsigned(1460976028,32),
    to_unsigned(1461126920,32),
    to_unsigned(1461277797,32),
    to_unsigned(1461428662,32),
    to_unsigned(1461579513,32),
    to_unsigned(1461730350,32),
    to_unsigned(1461881175,32),
    to_unsigned(1462031985,32),
    to_unsigned(1462182783,32),
    to_unsigned(1462333566,32),
    to_unsigned(1462484337,32),
    to_unsigned(1462635094,32),
    to_unsigned(1462785837,32),
    to_unsigned(1462936567,32),
    to_unsigned(1463087284,32),
    to_unsigned(1463237987,32),
    to_unsigned(1463388677,32),
    to_unsigned(1463539353,32),
    to_unsigned(1463690016,32),
    to_unsigned(1463840665,32),
    to_unsigned(1463991301,32),
    to_unsigned(1464141923,32),
    to_unsigned(1464292532,32),
    to_unsigned(1464443128,32),
    to_unsigned(1464593710,32),
    to_unsigned(1464744279,32),
    to_unsigned(1464894834,32),
    to_unsigned(1465045375,32),
    to_unsigned(1465195904,32),
    to_unsigned(1465346418,32),
    to_unsigned(1465496920,32),
    to_unsigned(1465647407,32),
    to_unsigned(1465797882,32),
    to_unsigned(1465948343,32),
    to_unsigned(1466098790,32),
    to_unsigned(1466249224,32),
    to_unsigned(1466399644,32),
    to_unsigned(1466550051,32),
    to_unsigned(1466700445,32),
    to_unsigned(1466850825,32),
    to_unsigned(1467001191,32),
    to_unsigned(1467151544,32),
    to_unsigned(1467301884,32),
    to_unsigned(1467452210,32),
    to_unsigned(1467602522,32),
    to_unsigned(1467752821,32),
    to_unsigned(1467903107,32),
    to_unsigned(1468053379,32),
    to_unsigned(1468203638,32),
    to_unsigned(1468353883,32),
    to_unsigned(1468504114,32),
    to_unsigned(1468654332,32),
    to_unsigned(1468804537,32),
    to_unsigned(1468954728,32),
    to_unsigned(1469104906,32),
    to_unsigned(1469255070,32),
    to_unsigned(1469405220,32),
    to_unsigned(1469555357,32),
    to_unsigned(1469705481,32),
    to_unsigned(1469855591,32),
    to_unsigned(1470005688,32),
    to_unsigned(1470155771,32),
    to_unsigned(1470305840,32),
    to_unsigned(1470455896,32),
    to_unsigned(1470605939,32),
    to_unsigned(1470755968,32),
    to_unsigned(1470905983,32),
    to_unsigned(1471055985,32),
    to_unsigned(1471205973,32),
    to_unsigned(1471355948,32),
    to_unsigned(1471505910,32),
    to_unsigned(1471655857,32),
    to_unsigned(1471805792,32),
    to_unsigned(1471955713,32),
    to_unsigned(1472105620,32),
    to_unsigned(1472255514,32),
    to_unsigned(1472405394,32),
    to_unsigned(1472555260,32),
    to_unsigned(1472705113,32),
    to_unsigned(1472854953,32),
    to_unsigned(1473004779,32),
    to_unsigned(1473154592,32),
    to_unsigned(1473304391,32),
    to_unsigned(1473454176,32),
    to_unsigned(1473603948,32),
    to_unsigned(1473753706,32),
    to_unsigned(1473903451,32),
    to_unsigned(1474053182,32),
    to_unsigned(1474202900,32),
    to_unsigned(1474352604,32),
    to_unsigned(1474502295,32),
    to_unsigned(1474651972,32),
    to_unsigned(1474801635,32),
    to_unsigned(1474951285,32),
    to_unsigned(1475100921,32),
    to_unsigned(1475250544,32),
    to_unsigned(1475400154,32),
    to_unsigned(1475549749,32),
    to_unsigned(1475699331,32),
    to_unsigned(1475848900,32),
    to_unsigned(1475998455,32),
    to_unsigned(1476147996,32),
    to_unsigned(1476297524,32),
    to_unsigned(1476447038,32),
    to_unsigned(1476596539,32),
    to_unsigned(1476746026,32),
    to_unsigned(1476895500,32),
    to_unsigned(1477044960,32),
    to_unsigned(1477194406,32),
    to_unsigned(1477343839,32),
    to_unsigned(1477493258,32),
    to_unsigned(1477642664,32),
    to_unsigned(1477792056,32),
    to_unsigned(1477941435,32),
    to_unsigned(1478090800,32),
    to_unsigned(1478240151,32),
    to_unsigned(1478389489,32),
    to_unsigned(1478538813,32),
    to_unsigned(1478688123,32),
    to_unsigned(1478837420,32),
    to_unsigned(1478986704,32),
    to_unsigned(1479135974,32),
    to_unsigned(1479285230,32),
    to_unsigned(1479434472,32),
    to_unsigned(1479583701,32),
    to_unsigned(1479732917,32),
    to_unsigned(1479882119,32),
    to_unsigned(1480031307,32),
    to_unsigned(1480180481,32),
    to_unsigned(1480329642,32),
    to_unsigned(1480478790,32),
    to_unsigned(1480627924,32),
    to_unsigned(1480777044,32),
    to_unsigned(1480926150,32),
    to_unsigned(1481075243,32),
    to_unsigned(1481224323,32),
    to_unsigned(1481373388,32),
    to_unsigned(1481522440,32),
    to_unsigned(1481671479,32),
    to_unsigned(1481820504,32),
    to_unsigned(1481969515,32),
    to_unsigned(1482118513,32),
    to_unsigned(1482267497,32),
    to_unsigned(1482416467,32),
    to_unsigned(1482565424,32),
    to_unsigned(1482714367,32),
    to_unsigned(1482863296,32),
    to_unsigned(1483012212,32),
    to_unsigned(1483161114,32),
    to_unsigned(1483310003,32),
    to_unsigned(1483458878,32),
    to_unsigned(1483607739,32),
    to_unsigned(1483756587,32),
    to_unsigned(1483905421,32),
    to_unsigned(1484054241,32),
    to_unsigned(1484203048,32),
    to_unsigned(1484351841,32),
    to_unsigned(1484500621,32),
    to_unsigned(1484649387,32),
    to_unsigned(1484798139,32),
    to_unsigned(1484946877,32),
    to_unsigned(1485095602,32),
    to_unsigned(1485244313,32),
    to_unsigned(1485393011,32),
    to_unsigned(1485541695,32),
    to_unsigned(1485690365,32),
    to_unsigned(1485839022,32),
    to_unsigned(1485987665,32),
    to_unsigned(1486136294,32),
    to_unsigned(1486284910,32),
    to_unsigned(1486433512,32),
    to_unsigned(1486582100,32),
    to_unsigned(1486730675,32),
    to_unsigned(1486879236,32),
    to_unsigned(1487027783,32),
    to_unsigned(1487176317,32),
    to_unsigned(1487324837,32),
    to_unsigned(1487473343,32),
    to_unsigned(1487621836,32),
    to_unsigned(1487770315,32),
    to_unsigned(1487918780,32),
    to_unsigned(1488067232,32),
    to_unsigned(1488215670,32),
    to_unsigned(1488364094,32),
    to_unsigned(1488512504,32),
    to_unsigned(1488660901,32),
    to_unsigned(1488809284,32),
    to_unsigned(1488957654,32),
    to_unsigned(1489106010,32),
    to_unsigned(1489254352,32),
    to_unsigned(1489402680,32),
    to_unsigned(1489550995,32),
    to_unsigned(1489699296,32),
    to_unsigned(1489847584,32),
    to_unsigned(1489995857,32),
    to_unsigned(1490144117,32),
    to_unsigned(1490292364,32),
    to_unsigned(1490440596,32),
    to_unsigned(1490588815,32),
    to_unsigned(1490737020,32),
    to_unsigned(1490885212,32),
    to_unsigned(1491033390,32),
    to_unsigned(1491181554,32),
    to_unsigned(1491329704,32),
    to_unsigned(1491477841,32),
    to_unsigned(1491625964,32),
    to_unsigned(1491774073,32),
    to_unsigned(1491922169,32),
    to_unsigned(1492070251,32),
    to_unsigned(1492218319,32),
    to_unsigned(1492366373,32),
    to_unsigned(1492514414,32),
    to_unsigned(1492662441,32),
    to_unsigned(1492810454,32),
    to_unsigned(1492958453,32),
    to_unsigned(1493106439,32),
    to_unsigned(1493254411,32),
    to_unsigned(1493402370,32),
    to_unsigned(1493550314,32),
    to_unsigned(1493698245,32),
    to_unsigned(1493846162,32),
    to_unsigned(1493994066,32),
    to_unsigned(1494141956,32),
    to_unsigned(1494289832,32),
    to_unsigned(1494437694,32),
    to_unsigned(1494585542,32),
    to_unsigned(1494733377,32),
    to_unsigned(1494881198,32),
    to_unsigned(1495029005,32),
    to_unsigned(1495176799,32),
    to_unsigned(1495324579,32),
    to_unsigned(1495472345,32),
    to_unsigned(1495620097,32),
    to_unsigned(1495767836,32),
    to_unsigned(1495915560,32),
    to_unsigned(1496063271,32),
    to_unsigned(1496210969,32),
    to_unsigned(1496358652,32),
    to_unsigned(1496506322,32),
    to_unsigned(1496653978,32),
    to_unsigned(1496801620,32),
    to_unsigned(1496949249,32),
    to_unsigned(1497096864,32),
    to_unsigned(1497244465,32),
    to_unsigned(1497392052,32),
    to_unsigned(1497539625,32),
    to_unsigned(1497687185,32),
    to_unsigned(1497834731,32),
    to_unsigned(1497982263,32),
    to_unsigned(1498129782,32),
    to_unsigned(1498277286,32),
    to_unsigned(1498424777,32),
    to_unsigned(1498572254,32),
    to_unsigned(1498719718,32),
    to_unsigned(1498867167,32),
    to_unsigned(1499014603,32),
    to_unsigned(1499162025,32),
    to_unsigned(1499309433,32),
    to_unsigned(1499456828,32),
    to_unsigned(1499604208,32),
    to_unsigned(1499751575,32),
    to_unsigned(1499898928,32),
    to_unsigned(1500046267,32),
    to_unsigned(1500193593,32),
    to_unsigned(1500340905,32),
    to_unsigned(1500488203,32),
    to_unsigned(1500635487,32),
    to_unsigned(1500782757,32),
    to_unsigned(1500930014,32),
    to_unsigned(1501077256,32),
    to_unsigned(1501224485,32),
    to_unsigned(1501371700,32),
    to_unsigned(1501518902,32),
    to_unsigned(1501666089,32),
    to_unsigned(1501813263,32),
    to_unsigned(1501960423,32),
    to_unsigned(1502107569,32),
    to_unsigned(1502254701,32),
    to_unsigned(1502401820,32),
    to_unsigned(1502548925,32),
    to_unsigned(1502696016,32),
    to_unsigned(1502843093,32),
    to_unsigned(1502990156,32),
    to_unsigned(1503137205,32),
    to_unsigned(1503284241,32),
    to_unsigned(1503431263,32),
    to_unsigned(1503578271,32),
    to_unsigned(1503725265,32),
    to_unsigned(1503872245,32),
    to_unsigned(1504019212,32),
    to_unsigned(1504166165,32),
    to_unsigned(1504313104,32),
    to_unsigned(1504460029,32),
    to_unsigned(1504606940,32),
    to_unsigned(1504753837,32),
    to_unsigned(1504900721,32),
    to_unsigned(1505047591,32),
    to_unsigned(1505194446,32),
    to_unsigned(1505341288,32),
    to_unsigned(1505488117,32),
    to_unsigned(1505634931,32),
    to_unsigned(1505781732,32),
    to_unsigned(1505928518,32),
    to_unsigned(1506075291,32),
    to_unsigned(1506222050,32),
    to_unsigned(1506368795,32),
    to_unsigned(1506515527,32),
    to_unsigned(1506662244,32),
    to_unsigned(1506808948,32),
    to_unsigned(1506955638,32),
    to_unsigned(1507102314,32),
    to_unsigned(1507248976,32),
    to_unsigned(1507395624,32),
    to_unsigned(1507542258,32),
    to_unsigned(1507688879,32),
    to_unsigned(1507835486,32),
    to_unsigned(1507982078,32),
    to_unsigned(1508128657,32),
    to_unsigned(1508275222,32),
    to_unsigned(1508421774,32),
    to_unsigned(1508568311,32),
    to_unsigned(1508714834,32),
    to_unsigned(1508861344,32),
    to_unsigned(1509007840,32),
    to_unsigned(1509154322,32),
    to_unsigned(1509300790,32),
    to_unsigned(1509447244,32),
    to_unsigned(1509593684,32),
    to_unsigned(1509740110,32),
    to_unsigned(1509886523,32),
    to_unsigned(1510032921,32),
    to_unsigned(1510179306,32),
    to_unsigned(1510325677,32),
    to_unsigned(1510472034,32),
    to_unsigned(1510618377,32),
    to_unsigned(1510764706,32),
    to_unsigned(1510911022,32),
    to_unsigned(1511057323,32),
    to_unsigned(1511203611,32),
    to_unsigned(1511349884,32),
    to_unsigned(1511496144,32),
    to_unsigned(1511642390,32),
    to_unsigned(1511788622,32),
    to_unsigned(1511934840,32),
    to_unsigned(1512081044,32),
    to_unsigned(1512227234,32),
    to_unsigned(1512373411,32),
    to_unsigned(1512519573,32),
    to_unsigned(1512665722,32),
    to_unsigned(1512811857,32),
    to_unsigned(1512957977,32),
    to_unsigned(1513104084,32),
    to_unsigned(1513250177,32),
    to_unsigned(1513396256,32),
    to_unsigned(1513542321,32),
    to_unsigned(1513688373,32),
    to_unsigned(1513834410,32),
    to_unsigned(1513980433,32),
    to_unsigned(1514126443,32),
    to_unsigned(1514272438,32),
    to_unsigned(1514418420,32),
    to_unsigned(1514564388,32),
    to_unsigned(1514710341,32),
    to_unsigned(1514856281,32),
    to_unsigned(1515002207,32),
    to_unsigned(1515148119,32),
    to_unsigned(1515294017,32),
    to_unsigned(1515439902,32),
    to_unsigned(1515585772,32),
    to_unsigned(1515731628,32),
    to_unsigned(1515877470,32),
    to_unsigned(1516023299,32),
    to_unsigned(1516169113,32),
    to_unsigned(1516314914,32),
    to_unsigned(1516460701,32),
    to_unsigned(1516606473,32),
    to_unsigned(1516752232,32),
    to_unsigned(1516897977,32),
    to_unsigned(1517043708,32),
    to_unsigned(1517189425,32),
    to_unsigned(1517335128,32),
    to_unsigned(1517480817,32),
    to_unsigned(1517626492,32),
    to_unsigned(1517772153,32),
    to_unsigned(1517917800,32),
    to_unsigned(1518063433,32),
    to_unsigned(1518209053,32),
    to_unsigned(1518354658,32),
    to_unsigned(1518500249,32),
    to_unsigned(1518645827,32),
    to_unsigned(1518791390,32),
    to_unsigned(1518936940,32),
    to_unsigned(1519082475,32),
    to_unsigned(1519227997,32),
    to_unsigned(1519373504,32),
    to_unsigned(1519518998,32),
    to_unsigned(1519664478,32),
    to_unsigned(1519809943,32),
    to_unsigned(1519955395,32),
    to_unsigned(1520100833,32),
    to_unsigned(1520246257,32),
    to_unsigned(1520391666,32),
    to_unsigned(1520537062,32),
    to_unsigned(1520682444,32),
    to_unsigned(1520827812,32),
    to_unsigned(1520973166,32),
    to_unsigned(1521118506,32),
    to_unsigned(1521263832,32),
    to_unsigned(1521409144,32),
    to_unsigned(1521554442,32),
    to_unsigned(1521699726,32),
    to_unsigned(1521844996,32),
    to_unsigned(1521990252,32),
    to_unsigned(1522135494,32),
    to_unsigned(1522280722,32),
    to_unsigned(1522425936,32),
    to_unsigned(1522571136,32),
    to_unsigned(1522716322,32),
    to_unsigned(1522861494,32),
    to_unsigned(1523006652,32),
    to_unsigned(1523151796,32),
    to_unsigned(1523296926,32),
    to_unsigned(1523442042,32),
    to_unsigned(1523587144,32),
    to_unsigned(1523732232,32),
    to_unsigned(1523877306,32),
    to_unsigned(1524022366,32),
    to_unsigned(1524167412,32),
    to_unsigned(1524312444,32),
    to_unsigned(1524457462,32),
    to_unsigned(1524602466,32),
    to_unsigned(1524747456,32),
    to_unsigned(1524892432,32),
    to_unsigned(1525037394,32),
    to_unsigned(1525182342,32),
    to_unsigned(1525327276,32),
    to_unsigned(1525472196,32),
    to_unsigned(1525617102,32),
    to_unsigned(1525761994,32),
    to_unsigned(1525906871,32),
    to_unsigned(1526051735,32),
    to_unsigned(1526196585,32),
    to_unsigned(1526341421,32),
    to_unsigned(1526486243,32),
    to_unsigned(1526631050,32),
    to_unsigned(1526775844,32),
    to_unsigned(1526920623,32),
    to_unsigned(1527065389,32),
    to_unsigned(1527210141,32),
    to_unsigned(1527354878,32),
    to_unsigned(1527499602,32),
    to_unsigned(1527644311,32),
    to_unsigned(1527789006,32),
    to_unsigned(1527933688,32),
    to_unsigned(1528078355,32),
    to_unsigned(1528223008,32),
    to_unsigned(1528367647,32),
    to_unsigned(1528512273,32),
    to_unsigned(1528656884,32),
    to_unsigned(1528801481,32),
    to_unsigned(1528946064,32),
    to_unsigned(1529090633,32),
    to_unsigned(1529235188,32),
    to_unsigned(1529379728,32),
    to_unsigned(1529524255,32),
    to_unsigned(1529668768,32),
    to_unsigned(1529813266,32),
    to_unsigned(1529957751,32),
    to_unsigned(1530102222,32),
    to_unsigned(1530246678,32),
    to_unsigned(1530391120,32),
    to_unsigned(1530535549,32),
    to_unsigned(1530679963,32),
    to_unsigned(1530824363,32),
    to_unsigned(1530968749,32),
    to_unsigned(1531113121,32),
    to_unsigned(1531257479,32),
    to_unsigned(1531401823,32),
    to_unsigned(1531546153,32),
    to_unsigned(1531690469,32),
    to_unsigned(1531834771,32),
    to_unsigned(1531979058,32),
    to_unsigned(1532123332,32),
    to_unsigned(1532267591,32),
    to_unsigned(1532411836,32),
    to_unsigned(1532556068,32),
    to_unsigned(1532700285,32),
    to_unsigned(1532844488,32),
    to_unsigned(1532988677,32),
    to_unsigned(1533132852,32),
    to_unsigned(1533277013,32),
    to_unsigned(1533421159,32),
    to_unsigned(1533565292,32),
    to_unsigned(1533709411,32),
    to_unsigned(1533853515,32),
    to_unsigned(1533997605,32),
    to_unsigned(1534141681,32),
    to_unsigned(1534285744,32),
    to_unsigned(1534429792,32),
    to_unsigned(1534573826,32),
    to_unsigned(1534717845,32),
    to_unsigned(1534861851,32),
    to_unsigned(1535005843,32),
    to_unsigned(1535149820,32),
    to_unsigned(1535293784,32),
    to_unsigned(1535437733,32),
    to_unsigned(1535581668,32),
    to_unsigned(1535725589,32),
    to_unsigned(1535869496,32),
    to_unsigned(1536013389,32),
    to_unsigned(1536157267,32),
    to_unsigned(1536301132,32),
    to_unsigned(1536444982,32),
    to_unsigned(1536588819,32),
    to_unsigned(1536732641,32),
    to_unsigned(1536876449,32),
    to_unsigned(1537020243,32),
    to_unsigned(1537164023,32),
    to_unsigned(1537307788,32),
    to_unsigned(1537451540,32),
    to_unsigned(1537595277,32),
    to_unsigned(1537739001,32),
    to_unsigned(1537882710,32),
    to_unsigned(1538026405,32),
    to_unsigned(1538170086,32),
    to_unsigned(1538313753,32),
    to_unsigned(1538457405,32),
    to_unsigned(1538601044,32),
    to_unsigned(1538744668,32),
    to_unsigned(1538888278,32),
    to_unsigned(1539031874,32),
    to_unsigned(1539175456,32),
    to_unsigned(1539319024,32),
    to_unsigned(1539462577,32),
    to_unsigned(1539606117,32),
    to_unsigned(1539749642,32),
    to_unsigned(1539893153,32),
    to_unsigned(1540036650,32),
    to_unsigned(1540180133,32),
    to_unsigned(1540323602,32),
    to_unsigned(1540467056,32),
    to_unsigned(1540610497,32),
    to_unsigned(1540753923,32),
    to_unsigned(1540897335,32),
    to_unsigned(1541040733,32),
    to_unsigned(1541184116,32),
    to_unsigned(1541327486,32),
    to_unsigned(1541470841,32),
    to_unsigned(1541614182,32),
    to_unsigned(1541757509,32),
    to_unsigned(1541900822,32),
    to_unsigned(1542044121,32),
    to_unsigned(1542187405,32),
    to_unsigned(1542330676,32),
    to_unsigned(1542473932,32),
    to_unsigned(1542617174,32),
    to_unsigned(1542760402,32),
    to_unsigned(1542903615,32),
    to_unsigned(1543046815,32),
    to_unsigned(1543190000,32),
    to_unsigned(1543333171,32),
    to_unsigned(1543476328,32),
    to_unsigned(1543619471,32),
    to_unsigned(1543762599,32),
    to_unsigned(1543905714,32),
    to_unsigned(1544048814,32),
    to_unsigned(1544191900,32),
    to_unsigned(1544334971,32),
    to_unsigned(1544478029,32),
    to_unsigned(1544621072,32),
    to_unsigned(1544764101,32),
    to_unsigned(1544907116,32),
    to_unsigned(1545050117,32),
    to_unsigned(1545193104,32),
    to_unsigned(1545336076,32),
    to_unsigned(1545479034,32),
    to_unsigned(1545621978,32),
    to_unsigned(1545764908,32),
    to_unsigned(1545907823,32),
    to_unsigned(1546050725,32),
    to_unsigned(1546193612,32),
    to_unsigned(1546336485,32),
    to_unsigned(1546479343,32),
    to_unsigned(1546622188,32),
    to_unsigned(1546765018,32),
    to_unsigned(1546907834,32),
    to_unsigned(1547050636,32),
    to_unsigned(1547193423,32),
    to_unsigned(1547336197,32),
    to_unsigned(1547478956,32),
    to_unsigned(1547621701,32),
    to_unsigned(1547764431,32),
    to_unsigned(1547907148,32),
    to_unsigned(1548049850,32),
    to_unsigned(1548192538,32),
    to_unsigned(1548335212,32),
    to_unsigned(1548477871,32),
    to_unsigned(1548620517,32),
    to_unsigned(1548763148,32),
    to_unsigned(1548905765,32),
    to_unsigned(1549048367,32),
    to_unsigned(1549190956,32),
    to_unsigned(1549333530,32),
    to_unsigned(1549476090,32),
    to_unsigned(1549618635,32),
    to_unsigned(1549761167,32),
    to_unsigned(1549903684,32),
    to_unsigned(1550046187,32),
    to_unsigned(1550188675,32),
    to_unsigned(1550331150,32),
    to_unsigned(1550473610,32),
    to_unsigned(1550616056,32),
    to_unsigned(1550758488,32),
    to_unsigned(1550900905,32),
    to_unsigned(1551043308,32),
    to_unsigned(1551185697,32),
    to_unsigned(1551328072,32),
    to_unsigned(1551470432,32),
    to_unsigned(1551612778,32),
    to_unsigned(1551755110,32),
    to_unsigned(1551897427,32),
    to_unsigned(1552039731,32),
    to_unsigned(1552182020,32),
    to_unsigned(1552324295,32),
    to_unsigned(1552466555,32),
    to_unsigned(1552608801,32),
    to_unsigned(1552751033,32),
    to_unsigned(1552893251,32),
    to_unsigned(1553035454,32),
    to_unsigned(1553177644,32),
    to_unsigned(1553319819,32),
    to_unsigned(1553461979,32),
    to_unsigned(1553604125,32),
    to_unsigned(1553746257,32),
    to_unsigned(1553888375,32),
    to_unsigned(1554030479,32),
    to_unsigned(1554172568,32),
    to_unsigned(1554314643,32),
    to_unsigned(1554456703,32),
    to_unsigned(1554598750,32),
    to_unsigned(1554740782,32),
    to_unsigned(1554882800,32),
    to_unsigned(1555024803,32),
    to_unsigned(1555166792,32),
    to_unsigned(1555308767,32),
    to_unsigned(1555450728,32),
    to_unsigned(1555592674,32),
    to_unsigned(1555734606,32),
    to_unsigned(1555876524,32),
    to_unsigned(1556018427,32),
    to_unsigned(1556160316,32),
    to_unsigned(1556302191,32),
    to_unsigned(1556444051,32),
    to_unsigned(1556585897,32),
    to_unsigned(1556727729,32),
    to_unsigned(1556869547,32),
    to_unsigned(1557011350,32),
    to_unsigned(1557153139,32),
    to_unsigned(1557294914,32),
    to_unsigned(1557436674,32),
    to_unsigned(1557578420,32),
    to_unsigned(1557720151,32),
    to_unsigned(1557861869,32),
    to_unsigned(1558003572,32),
    to_unsigned(1558145260,32),
    to_unsigned(1558286935,32),
    to_unsigned(1558428595,32),
    to_unsigned(1558570241,32),
    to_unsigned(1558711872,32),
    to_unsigned(1558853489,32),
    to_unsigned(1558995092,32),
    to_unsigned(1559136680,32),
    to_unsigned(1559278254,32),
    to_unsigned(1559419814,32),
    to_unsigned(1559561360,32),
    to_unsigned(1559702891,32),
    to_unsigned(1559844407,32),
    to_unsigned(1559985910,32),
    to_unsigned(1560127398,32),
    to_unsigned(1560268872,32),
    to_unsigned(1560410331,32),
    to_unsigned(1560551776,32),
    to_unsigned(1560693207,32),
    to_unsigned(1560834623,32),
    to_unsigned(1560976025,32),
    to_unsigned(1561117413,32),
    to_unsigned(1561258786,32),
    to_unsigned(1561400145,32),
    to_unsigned(1561541490,32),
    to_unsigned(1561682820,32),
    to_unsigned(1561824136,32),
    to_unsigned(1561965437,32),
    to_unsigned(1562106725,32),
    to_unsigned(1562247997,32),
    to_unsigned(1562389256,32),
    to_unsigned(1562530500,32),
    to_unsigned(1562671730,32),
    to_unsigned(1562812945,32),
    to_unsigned(1562954146,32),
    to_unsigned(1563095333,32),
    to_unsigned(1563236505,32),
    to_unsigned(1563377663,32),
    to_unsigned(1563518806,32),
    to_unsigned(1563659936,32),
    to_unsigned(1563801050,32),
    to_unsigned(1563942151,32),
    to_unsigned(1564083237,32),
    to_unsigned(1564224309,32),
    to_unsigned(1564365366,32),
    to_unsigned(1564506409,32),
    to_unsigned(1564647437,32),
    to_unsigned(1564788452,32),
    to_unsigned(1564929451,32),
    to_unsigned(1565070437,32),
    to_unsigned(1565211408,32),
    to_unsigned(1565352364,32),
    to_unsigned(1565493307,32),
    to_unsigned(1565634234,32),
    to_unsigned(1565775148,32),
    to_unsigned(1565916047,32),
    to_unsigned(1566056931,32),
    to_unsigned(1566197802,32),
    to_unsigned(1566338658,32),
    to_unsigned(1566479499,32),
    to_unsigned(1566620326,32),
    to_unsigned(1566761139,32),
    to_unsigned(1566901937,32),
    to_unsigned(1567042721,32),
    to_unsigned(1567183490,32),
    to_unsigned(1567324246,32),
    to_unsigned(1567464986,32),
    to_unsigned(1567605712,32),
    to_unsigned(1567746424,32),
    to_unsigned(1567887122,32),
    to_unsigned(1568027805,32),
    to_unsigned(1568168473,32),
    to_unsigned(1568309127,32),
    to_unsigned(1568449767,32),
    to_unsigned(1568590393,32),
    to_unsigned(1568731004,32),
    to_unsigned(1568871600,32),
    to_unsigned(1569012182,32),
    to_unsigned(1569152750,32),
    to_unsigned(1569293303,32),
    to_unsigned(1569433842,32),
    to_unsigned(1569574366,32),
    to_unsigned(1569714876,32),
    to_unsigned(1569855372,32),
    to_unsigned(1569995853,32),
    to_unsigned(1570136320,32),
    to_unsigned(1570276772,32),
    to_unsigned(1570417210,32),
    to_unsigned(1570557633,32),
    to_unsigned(1570698042,32),
    to_unsigned(1570838436,32),
    to_unsigned(1570978817,32),
    to_unsigned(1571119182,32),
    to_unsigned(1571259533,32),
    to_unsigned(1571399870,32),
    to_unsigned(1571540192,32),
    to_unsigned(1571680500,32),
    to_unsigned(1571820794,32),
    to_unsigned(1571961073,32),
    to_unsigned(1572101337,32),
    to_unsigned(1572241587,32),
    to_unsigned(1572381823,32),
    to_unsigned(1572522044,32),
    to_unsigned(1572662251,32),
    to_unsigned(1572802443,32),
    to_unsigned(1572942621,32),
    to_unsigned(1573082784,32),
    to_unsigned(1573222933,32),
    to_unsigned(1573363067,32),
    to_unsigned(1573503187,32),
    to_unsigned(1573643293,32),
    to_unsigned(1573783384,32),
    to_unsigned(1573923460,32),
    to_unsigned(1574063522,32),
    to_unsigned(1574203570,32),
    to_unsigned(1574343603,32),
    to_unsigned(1574483622,32),
    to_unsigned(1574623626,32),
    to_unsigned(1574763616,32),
    to_unsigned(1574903591,32),
    to_unsigned(1575043552,32),
    to_unsigned(1575183498,32),
    to_unsigned(1575323430,32),
    to_unsigned(1575463347,32),
    to_unsigned(1575603250,32),
    to_unsigned(1575743139,32),
    to_unsigned(1575883012,32),
    to_unsigned(1576022872,32),
    to_unsigned(1576162717,32),
    to_unsigned(1576302547,32),
    to_unsigned(1576442363,32),
    to_unsigned(1576582165,32),
    to_unsigned(1576721952,32),
    to_unsigned(1576861724,32),
    to_unsigned(1577001482,32),
    to_unsigned(1577141226,32),
    to_unsigned(1577280955,32),
    to_unsigned(1577420669,32),
    to_unsigned(1577560369,32),
    to_unsigned(1577700055,32),
    to_unsigned(1577839726,32),
    to_unsigned(1577979382,32),
    to_unsigned(1578119024,32),
    to_unsigned(1578258651,32),
    to_unsigned(1578398264,32),
    to_unsigned(1578537863,32),
    to_unsigned(1578677447,32),
    to_unsigned(1578817016,32),
    to_unsigned(1578956571,32),
    to_unsigned(1579096112,32),
    to_unsigned(1579235638,32),
    to_unsigned(1579375149,32),
    to_unsigned(1579514646,32),
    to_unsigned(1579654128,32),
    to_unsigned(1579793596,32),
    to_unsigned(1579933049,32),
    to_unsigned(1580072488,32),
    to_unsigned(1580211912,32),
    to_unsigned(1580351322,32),
    to_unsigned(1580490717,32),
    to_unsigned(1580630098,32),
    to_unsigned(1580769464,32),
    to_unsigned(1580908816,32),
    to_unsigned(1581048153,32),
    to_unsigned(1581187475,32),
    to_unsigned(1581326783,32),
    to_unsigned(1581466077,32),
    to_unsigned(1581605356,32),
    to_unsigned(1581744620,32),
    to_unsigned(1581883870,32),
    to_unsigned(1582023105,32),
    to_unsigned(1582162326,32),
    to_unsigned(1582301533,32),
    to_unsigned(1582440724,32),
    to_unsigned(1582579901,32),
    to_unsigned(1582719064,32),
    to_unsigned(1582858212,32),
    to_unsigned(1582997346,32),
    to_unsigned(1583136465,32),
    to_unsigned(1583275569,32),
    to_unsigned(1583414659,32),
    to_unsigned(1583553734,32),
    to_unsigned(1583692795,32),
    to_unsigned(1583831841,32),
    to_unsigned(1583970873,32),
    to_unsigned(1584109890,32),
    to_unsigned(1584248892,32),
    to_unsigned(1584387880,32),
    to_unsigned(1584526854,32),
    to_unsigned(1584665812,32),
    to_unsigned(1584804757,32),
    to_unsigned(1584943686,32),
    to_unsigned(1585082602,32),
    to_unsigned(1585221502,32),
    to_unsigned(1585360388,32),
    to_unsigned(1585499260,32),
    to_unsigned(1585638116,32),
    to_unsigned(1585776959,32),
    to_unsigned(1585915786,32),
    to_unsigned(1586054599,32),
    to_unsigned(1586193398,32),
    to_unsigned(1586332182,32),
    to_unsigned(1586470951,32),
    to_unsigned(1586609706,32),
    to_unsigned(1586748446,32),
    to_unsigned(1586887172,32),
    to_unsigned(1587025883,32),
    to_unsigned(1587164579,32),
    to_unsigned(1587303261,32),
    to_unsigned(1587441928,32),
    to_unsigned(1587580581,32),
    to_unsigned(1587719219,32),
    to_unsigned(1587857843,32),
    to_unsigned(1587996452,32),
    to_unsigned(1588135046,32),
    to_unsigned(1588273626,32),
    to_unsigned(1588412191,32),
    to_unsigned(1588550741,32),
    to_unsigned(1588689277,32),
    to_unsigned(1588827798,32),
    to_unsigned(1588966305,32),
    to_unsigned(1589104797,32),
    to_unsigned(1589243275,32),
    to_unsigned(1589381738,32),
    to_unsigned(1589520186,32),
    to_unsigned(1589658619,32),
    to_unsigned(1589797038,32),
    to_unsigned(1589935443,32),
    to_unsigned(1590073833,32),
    to_unsigned(1590212208,32),
    to_unsigned(1590350568,32),
    to_unsigned(1590488914,32),
    to_unsigned(1590627246,32),
    to_unsigned(1590765563,32),
    to_unsigned(1590903865,32),
    to_unsigned(1591042152,32),
    to_unsigned(1591180425,32),
    to_unsigned(1591318683,32),
    to_unsigned(1591456927,32),
    to_unsigned(1591595156,32),
    to_unsigned(1591733370,32),
    to_unsigned(1591871570,32),
    to_unsigned(1592009755,32),
    to_unsigned(1592147925,32),
    to_unsigned(1592286081,32),
    to_unsigned(1592424222,32),
    to_unsigned(1592562349,32),
    to_unsigned(1592700461,32),
    to_unsigned(1592838558,32),
    to_unsigned(1592976641,32),
    to_unsigned(1593114709,32),
    to_unsigned(1593252762,32),
    to_unsigned(1593390801,32),
    to_unsigned(1593528825,32),
    to_unsigned(1593666834,32),
    to_unsigned(1593804829,32),
    to_unsigned(1593942809,32),
    to_unsigned(1594080774,32),
    to_unsigned(1594218725,32),
    to_unsigned(1594356661,32),
    to_unsigned(1594494583,32),
    to_unsigned(1594632490,32),
    to_unsigned(1594770382,32),
    to_unsigned(1594908259,32),
    to_unsigned(1595046122,32),
    to_unsigned(1595183970,32),
    to_unsigned(1595321804,32),
    to_unsigned(1595459623,32),
    to_unsigned(1595597427,32),
    to_unsigned(1595735216,32),
    to_unsigned(1595872991,32),
    to_unsigned(1596010751,32),
    to_unsigned(1596148497,32),
    to_unsigned(1596286228,32),
    to_unsigned(1596423944,32),
    to_unsigned(1596561645,32),
    to_unsigned(1596699332,32),
    to_unsigned(1596837004,32),
    to_unsigned(1596974662,32),
    to_unsigned(1597112305,32),
    to_unsigned(1597249933,32),
    to_unsigned(1597387546,32),
    to_unsigned(1597525145,32),
    to_unsigned(1597662729,32),
    to_unsigned(1597800298,32),
    to_unsigned(1597937853,32),
    to_unsigned(1598075393,32),
    to_unsigned(1598212918,32),
    to_unsigned(1598350429,32),
    to_unsigned(1598487925,32),
    to_unsigned(1598625406,32),
    to_unsigned(1598762873,32),
    to_unsigned(1598900325,32),
    to_unsigned(1599037762,32),
    to_unsigned(1599175184,32),
    to_unsigned(1599312592,32),
    to_unsigned(1599449985,32),
    to_unsigned(1599587363,32),
    to_unsigned(1599724727,32),
    to_unsigned(1599862076,32),
    to_unsigned(1599999410,32),
    to_unsigned(1600136730,32),
    to_unsigned(1600274035,32),
    to_unsigned(1600411325,32),
    to_unsigned(1600548600,32),
    to_unsigned(1600685861,32),
    to_unsigned(1600823107,32),
    to_unsigned(1600960338,32),
    to_unsigned(1601097555,32),
    to_unsigned(1601234757,32),
    to_unsigned(1601371944,32),
    to_unsigned(1601509116,32),
    to_unsigned(1601646274,32),
    to_unsigned(1601783417,32),
    to_unsigned(1601920545,32),
    to_unsigned(1602057658,32),
    to_unsigned(1602194757,32),
    to_unsigned(1602331841,32),
    to_unsigned(1602468911,32),
    to_unsigned(1602605965,32),
    to_unsigned(1602743005,32),
    to_unsigned(1602880030,32),
    to_unsigned(1603017041,32),
    to_unsigned(1603154036,32),
    to_unsigned(1603291017,32),
    to_unsigned(1603427983,32),
    to_unsigned(1603564935,32),
    to_unsigned(1603701872,32),
    to_unsigned(1603838794,32),
    to_unsigned(1603975701,32),
    to_unsigned(1604112593,32),
    to_unsigned(1604249471,32),
    to_unsigned(1604386334,32),
    to_unsigned(1604523182,32),
    to_unsigned(1604660016,32),
    to_unsigned(1604796835,32),
    to_unsigned(1604933639,32),
    to_unsigned(1605070428,32),
    to_unsigned(1605207202,32),
    to_unsigned(1605343962,32),
    to_unsigned(1605480707,32),
    to_unsigned(1605617437,32),
    to_unsigned(1605754153,32),
    to_unsigned(1605890853,32),
    to_unsigned(1606027539,32),
    to_unsigned(1606164211,32),
    to_unsigned(1606300867,32),
    to_unsigned(1606437509,32),
    to_unsigned(1606574136,32),
    to_unsigned(1606710748,32),
    to_unsigned(1606847345,32),
    to_unsigned(1606983928,32),
    to_unsigned(1607120495,32),
    to_unsigned(1607257048,32),
    to_unsigned(1607393587,32),
    to_unsigned(1607530110,32),
    to_unsigned(1607666619,32),
    to_unsigned(1607803113,32),
    to_unsigned(1607939592,32),
    to_unsigned(1608076056,32),
    to_unsigned(1608212506,32),
    to_unsigned(1608348941,32),
    to_unsigned(1608485361,32),
    to_unsigned(1608621766,32),
    to_unsigned(1608758157,32),
    to_unsigned(1608894532,32),
    to_unsigned(1609030893,32),
    to_unsigned(1609167239,32),
    to_unsigned(1609303571,32),
    to_unsigned(1609439887,32),
    to_unsigned(1609576189,32),
    to_unsigned(1609712476,32),
    to_unsigned(1609848748,32),
    to_unsigned(1609985005,32),
    to_unsigned(1610121248,32),
    to_unsigned(1610257475,32),
    to_unsigned(1610393688,32),
    to_unsigned(1610529887,32),
    to_unsigned(1610666070,32),
    to_unsigned(1610802238,32),
    to_unsigned(1610938392,32),
    to_unsigned(1611074531,32),
    to_unsigned(1611210655,32),
    to_unsigned(1611346764,32),
    to_unsigned(1611482859,32),
    to_unsigned(1611618939,32),
    to_unsigned(1611755003,32),
    to_unsigned(1611891053,32),
    to_unsigned(1612027089,32),
    to_unsigned(1612163109,32),
    to_unsigned(1612299115,32),
    to_unsigned(1612435105,32),
    to_unsigned(1612571081,32),
    to_unsigned(1612707043,32),
    to_unsigned(1612842989,32),
    to_unsigned(1612978920,32),
    to_unsigned(1613114837,32),
    to_unsigned(1613250739,32),
    to_unsigned(1613386626,32),
    to_unsigned(1613522498,32),
    to_unsigned(1613658355,32),
    to_unsigned(1613794198,32),
    to_unsigned(1613930025,32),
    to_unsigned(1614065838,32),
    to_unsigned(1614201636,32),
    to_unsigned(1614337419,32),
    to_unsigned(1614473188,32),
    to_unsigned(1614608941,32),
    to_unsigned(1614744680,32),
    to_unsigned(1614880404,32),
    to_unsigned(1615016113,32),
    to_unsigned(1615151807,32),
    to_unsigned(1615287486,32),
    to_unsigned(1615423150,32),
    to_unsigned(1615558800,32),
    to_unsigned(1615694435,32),
    to_unsigned(1615830055,32),
    to_unsigned(1615965660,32),
    to_unsigned(1616101250,32),
    to_unsigned(1616236825,32),
    to_unsigned(1616372385,32),
    to_unsigned(1616507931,32),
    to_unsigned(1616643462,32),
    to_unsigned(1616778978,32),
    to_unsigned(1616914479,32),
    to_unsigned(1617049965,32),
    to_unsigned(1617185436,32),
    to_unsigned(1617320893,32),
    to_unsigned(1617456334,32),
    to_unsigned(1617591761,32),
    to_unsigned(1617727173,32),
    to_unsigned(1617862570,32),
    to_unsigned(1617997952,32),
    to_unsigned(1618133319,32),
    to_unsigned(1618268671,32),
    to_unsigned(1618404009,32),
    to_unsigned(1618539331,32),
    to_unsigned(1618674639,32),
    to_unsigned(1618809932,32),
    to_unsigned(1618945210,32),
    to_unsigned(1619080473,32),
    to_unsigned(1619215721,32),
    to_unsigned(1619350954,32),
    to_unsigned(1619486173,32),
    to_unsigned(1619621376,32),
    to_unsigned(1619756565,32),
    to_unsigned(1619891739,32),
    to_unsigned(1620026897,32),
    to_unsigned(1620162041,32),
    to_unsigned(1620297170,32),
    to_unsigned(1620432285,32),
    to_unsigned(1620567384,32),
    to_unsigned(1620702468,32),
    to_unsigned(1620837538,32),
    to_unsigned(1620972592,32),
    to_unsigned(1621107632,32),
    to_unsigned(1621242657,32),
    to_unsigned(1621377667,32),
    to_unsigned(1621512662,32),
    to_unsigned(1621647642,32),
    to_unsigned(1621782607,32),
    to_unsigned(1621917557,32),
    to_unsigned(1622052493,32),
    to_unsigned(1622187413,32),
    to_unsigned(1622322319,32),
    to_unsigned(1622457209,32),
    to_unsigned(1622592085,32),
    to_unsigned(1622726946,32),
    to_unsigned(1622861792,32),
    to_unsigned(1622996623,32),
    to_unsigned(1623131439,32),
    to_unsigned(1623266240,32),
    to_unsigned(1623401026,32),
    to_unsigned(1623535797,32),
    to_unsigned(1623670554,32),
    to_unsigned(1623805295,32),
    to_unsigned(1623940022,32),
    to_unsigned(1624074733,32),
    to_unsigned(1624209430,32),
    to_unsigned(1624344112,32),
    to_unsigned(1624478779,32),
    to_unsigned(1624613430,32),
    to_unsigned(1624748067,32),
    to_unsigned(1624882689,32),
    to_unsigned(1625017296,32),
    to_unsigned(1625151889,32),
    to_unsigned(1625286466,32),
    to_unsigned(1625421028,32),
    to_unsigned(1625555575,32),
    to_unsigned(1625690108,32),
    to_unsigned(1625824625,32),
    to_unsigned(1625959128,32),
    to_unsigned(1626093615,32),
    to_unsigned(1626228088,32),
    to_unsigned(1626362545,32),
    to_unsigned(1626496988,32),
    to_unsigned(1626631416,32),
    to_unsigned(1626765829,32),
    to_unsigned(1626900227,32),
    to_unsigned(1627034609,32),
    to_unsigned(1627168977,32),
    to_unsigned(1627303330,32),
    to_unsigned(1627437668,32),
    to_unsigned(1627571991,32),
    to_unsigned(1627706300,32),
    to_unsigned(1627840593,32),
    to_unsigned(1627974871,32),
    to_unsigned(1628109134,32),
    to_unsigned(1628243382,32),
    to_unsigned(1628377616,32),
    to_unsigned(1628511834,32),
    to_unsigned(1628646037,32),
    to_unsigned(1628780226,32),
    to_unsigned(1628914399,32),
    to_unsigned(1629048557,32),
    to_unsigned(1629182701,32),
    to_unsigned(1629316829,32),
    to_unsigned(1629450943,32),
    to_unsigned(1629585041,32),
    to_unsigned(1629719125,32),
    to_unsigned(1629853194,32),
    to_unsigned(1629987247,32),
    to_unsigned(1630121286,32),
    to_unsigned(1630255309,32),
    to_unsigned(1630389318,32),
    to_unsigned(1630523312,32),
    to_unsigned(1630657290,32),
    to_unsigned(1630791254,32),
    to_unsigned(1630925203,32),
    to_unsigned(1631059136,32),
    to_unsigned(1631193055,32),
    to_unsigned(1631326959,32),
    to_unsigned(1631460847,32),
    to_unsigned(1631594721,32),
    to_unsigned(1631728580,32),
    to_unsigned(1631862424,32),
    to_unsigned(1631996252,32),
    to_unsigned(1632130066,32),
    to_unsigned(1632263865,32),
    to_unsigned(1632397648,32),
    to_unsigned(1632531417,32),
    to_unsigned(1632665171,32),
    to_unsigned(1632798910,32),
    to_unsigned(1632932633,32),
    to_unsigned(1633066342,32),
    to_unsigned(1633200036,32),
    to_unsigned(1633333714,32),
    to_unsigned(1633467378,32),
    to_unsigned(1633601027,32),
    to_unsigned(1633734660,32),
    to_unsigned(1633868279,32),
    to_unsigned(1634001882,32),
    to_unsigned(1634135471,32),
    to_unsigned(1634269044,32),
    to_unsigned(1634402603,32),
    to_unsigned(1634536146,32),
    to_unsigned(1634669675,32),
    to_unsigned(1634803188,32),
    to_unsigned(1634936687,32),
    to_unsigned(1635070170,32),
    to_unsigned(1635203638,32),
    to_unsigned(1635337092,32),
    to_unsigned(1635470530,32),
    to_unsigned(1635603953,32),
    to_unsigned(1635737362,32),
    to_unsigned(1635870755,32),
    to_unsigned(1636004133,32),
    to_unsigned(1636137496,32),
    to_unsigned(1636270844,32),
    to_unsigned(1636404177,32),
    to_unsigned(1636537495,32),
    to_unsigned(1636670798,32),
    to_unsigned(1636804086,32),
    to_unsigned(1636937359,32),
    to_unsigned(1637070617,32),
    to_unsigned(1637203860,32),
    to_unsigned(1637337087,32),
    to_unsigned(1637470300,32),
    to_unsigned(1637603498,32),
    to_unsigned(1637736680,32),
    to_unsigned(1637869848,32),
    to_unsigned(1638003000,32),
    to_unsigned(1638136137,32),
    to_unsigned(1638269260,32),
    to_unsigned(1638402367,32),
    to_unsigned(1638535459,32),
    to_unsigned(1638668537,32),
    to_unsigned(1638801599,32),
    to_unsigned(1638934646,32),
    to_unsigned(1639067678,32),
    to_unsigned(1639200695,32),
    to_unsigned(1639333696,32),
    to_unsigned(1639466683,32),
    to_unsigned(1639599655,32),
    to_unsigned(1639732612,32),
    to_unsigned(1639865553,32),
    to_unsigned(1639998480,32),
    to_unsigned(1640131391,32),
    to_unsigned(1640264287,32),
    to_unsigned(1640397169,32),
    to_unsigned(1640530035,32),
    to_unsigned(1640662886,32),
    to_unsigned(1640795722,32),
    to_unsigned(1640928543,32),
    to_unsigned(1641061349,32),
    to_unsigned(1641194139,32),
    to_unsigned(1641326915,32),
    to_unsigned(1641459676,32),
    to_unsigned(1641592421,32),
    to_unsigned(1641725152,32),
    to_unsigned(1641857867,32),
    to_unsigned(1641990567,32),
    to_unsigned(1642123252,32),
    to_unsigned(1642255922,32),
    to_unsigned(1642388577,32),
    to_unsigned(1642521217,32),
    to_unsigned(1642653842,32),
    to_unsigned(1642786452,32),
    to_unsigned(1642919046,32),
    to_unsigned(1643051626,32),
    to_unsigned(1643184190,32),
    to_unsigned(1643316739,32),
    to_unsigned(1643449274,32),
    to_unsigned(1643581793,32),
    to_unsigned(1643714297,32),
    to_unsigned(1643846785,32),
    to_unsigned(1643979259,32),
    to_unsigned(1644111718,32),
    to_unsigned(1644244161,32),
    to_unsigned(1644376590,32),
    to_unsigned(1644509003,32),
    to_unsigned(1644641401,32),
    to_unsigned(1644773784,32),
    to_unsigned(1644906152,32),
    to_unsigned(1645038505,32),
    to_unsigned(1645170842,32),
    to_unsigned(1645303165,32),
    to_unsigned(1645435472,32),
    to_unsigned(1645567765,32),
    to_unsigned(1645700042,32),
    to_unsigned(1645832304,32),
    to_unsigned(1645964551,32),
    to_unsigned(1646096783,32),
    to_unsigned(1646228999,32),
    to_unsigned(1646361201,32),
    to_unsigned(1646493387,32),
    to_unsigned(1646625559,32),
    to_unsigned(1646757715,32),
    to_unsigned(1646889856,32),
    to_unsigned(1647021982,32),
    to_unsigned(1647154092,32),
    to_unsigned(1647286188,32),
    to_unsigned(1647418268,32),
    to_unsigned(1647550334,32),
    to_unsigned(1647682384,32),
    to_unsigned(1647814419,32),
    to_unsigned(1647946439,32),
    to_unsigned(1648078443,32),
    to_unsigned(1648210433,32),
    to_unsigned(1648342407,32),
    to_unsigned(1648474367,32),
    to_unsigned(1648606311,32),
    to_unsigned(1648738240,32),
    to_unsigned(1648870154,32),
    to_unsigned(1649002052,32),
    to_unsigned(1649133936,32),
    to_unsigned(1649265804,32),
    to_unsigned(1649397657,32),
    to_unsigned(1649529495,32),
    to_unsigned(1649661318,32),
    to_unsigned(1649793126,32),
    to_unsigned(1649924918,32),
    to_unsigned(1650056696,32),
    to_unsigned(1650188458,32),
    to_unsigned(1650320205,32),
    to_unsigned(1650451937,32),
    to_unsigned(1650583653,32),
    to_unsigned(1650715355,32),
    to_unsigned(1650847041,32),
    to_unsigned(1650978712,32),
    to_unsigned(1651110368,32),
    to_unsigned(1651242009,32),
    to_unsigned(1651373635,32),
    to_unsigned(1651505245,32),
    to_unsigned(1651636840,32),
    to_unsigned(1651768421,32),
    to_unsigned(1651899985,32),
    to_unsigned(1652031535,32),
    to_unsigned(1652163070,32),
    to_unsigned(1652294589,32),
    to_unsigned(1652426093,32),
    to_unsigned(1652557582,32),
    to_unsigned(1652689056,32),
    to_unsigned(1652820515,32),
    to_unsigned(1652951958,32),
    to_unsigned(1653083386,32),
    to_unsigned(1653214799,32),
    to_unsigned(1653346197,32),
    to_unsigned(1653477580,32),
    to_unsigned(1653608947,32),
    to_unsigned(1653740299,32),
    to_unsigned(1653871636,32),
    to_unsigned(1654002958,32),
    to_unsigned(1654134265,32),
    to_unsigned(1654265556,32),
    to_unsigned(1654396832,32),
    to_unsigned(1654528093,32),
    to_unsigned(1654659339,32),
    to_unsigned(1654790570,32),
    to_unsigned(1654921785,32),
    to_unsigned(1655052985,32),
    to_unsigned(1655184170,32),
    to_unsigned(1655315340,32),
    to_unsigned(1655446494,32),
    to_unsigned(1655577634,32),
    to_unsigned(1655708758,32),
    to_unsigned(1655839867,32),
    to_unsigned(1655970960,32),
    to_unsigned(1656102039,32),
    to_unsigned(1656233102,32),
    to_unsigned(1656364150,32),
    to_unsigned(1656495183,32),
    to_unsigned(1656626200,32),
    to_unsigned(1656757203,32),
    to_unsigned(1656888190,32),
    to_unsigned(1657019161,32),
    to_unsigned(1657150118,32),
    to_unsigned(1657281059,32),
    to_unsigned(1657411986,32),
    to_unsigned(1657542896,32),
    to_unsigned(1657673792,32),
    to_unsigned(1657804673,32),
    to_unsigned(1657935538,32),
    to_unsigned(1658066388,32),
    to_unsigned(1658197222,32),
    to_unsigned(1658328042,32),
    to_unsigned(1658458846,32),
    to_unsigned(1658589635,32),
    to_unsigned(1658720409,32),
    to_unsigned(1658851167,32),
    to_unsigned(1658981911,32),
    to_unsigned(1659112639,32),
    to_unsigned(1659243351,32),
    to_unsigned(1659374049,32),
    to_unsigned(1659504731,32),
    to_unsigned(1659635398,32),
    to_unsigned(1659766050,32),
    to_unsigned(1659896686,32),
    to_unsigned(1660027308,32),
    to_unsigned(1660157914,32),
    to_unsigned(1660288504,32),
    to_unsigned(1660419080,32),
    to_unsigned(1660549640,32),
    to_unsigned(1660680185,32),
    to_unsigned(1660810714,32),
    to_unsigned(1660941229,32),
    to_unsigned(1661071728,32),
    to_unsigned(1661202212,32),
    to_unsigned(1661332680,32),
    to_unsigned(1661463134,32),
    to_unsigned(1661593572,32),
    to_unsigned(1661723994,32),
    to_unsigned(1661854402,32),
    to_unsigned(1661984794,32),
    to_unsigned(1662115171,32),
    to_unsigned(1662245533,32),
    to_unsigned(1662375879,32),
    to_unsigned(1662506210,32),
    to_unsigned(1662636526,32),
    to_unsigned(1662766827,32),
    to_unsigned(1662897112,32),
    to_unsigned(1663027382,32),
    to_unsigned(1663157637,32),
    to_unsigned(1663287876,32),
    to_unsigned(1663418100,32),
    to_unsigned(1663548309,32),
    to_unsigned(1663678502,32),
    to_unsigned(1663808681,32),
    to_unsigned(1663938844,32),
    to_unsigned(1664068991,32),
    to_unsigned(1664199124,32),
    to_unsigned(1664329241,32),
    to_unsigned(1664459342,32),
    to_unsigned(1664589429,32),
    to_unsigned(1664719500,32),
    to_unsigned(1664849556,32),
    to_unsigned(1664979596,32),
    to_unsigned(1665109622,32),
    to_unsigned(1665239632,32),
    to_unsigned(1665369626,32),
    to_unsigned(1665499606,32),
    to_unsigned(1665629570,32),
    to_unsigned(1665759518,32),
    to_unsigned(1665889452,32),
    to_unsigned(1666019370,32),
    to_unsigned(1666149273,32),
    to_unsigned(1666279160,32),
    to_unsigned(1666409032,32),
    to_unsigned(1666538889,32),
    to_unsigned(1666668731,32),
    to_unsigned(1666798557,32),
    to_unsigned(1666928368,32),
    to_unsigned(1667058163,32),
    to_unsigned(1667187943,32),
    to_unsigned(1667317708,32),
    to_unsigned(1667447458,32),
    to_unsigned(1667577192,32),
    to_unsigned(1667706911,32),
    to_unsigned(1667836615,32),
    to_unsigned(1667966303,32),
    to_unsigned(1668095976,32),
    to_unsigned(1668225633,32),
    to_unsigned(1668355276,32),
    to_unsigned(1668484902,32),
    to_unsigned(1668614514,32),
    to_unsigned(1668744110,32),
    to_unsigned(1668873691,32),
    to_unsigned(1669003257,32),
    to_unsigned(1669132807,32),
    to_unsigned(1669262342,32),
    to_unsigned(1669391861,32),
    to_unsigned(1669521366,32),
    to_unsigned(1669650855,32),
    to_unsigned(1669780328,32),
    to_unsigned(1669909786,32),
    to_unsigned(1670039229,32),
    to_unsigned(1670168656,32),
    to_unsigned(1670298069,32),
    to_unsigned(1670427465,32),
    to_unsigned(1670556847,32),
    to_unsigned(1670686213,32),
    to_unsigned(1670815563,32),
    to_unsigned(1670944899,32),
    to_unsigned(1671074219,32),
    to_unsigned(1671203523,32),
    to_unsigned(1671332813,32),
    to_unsigned(1671462086,32),
    to_unsigned(1671591345,32),
    to_unsigned(1671720588,32),
    to_unsigned(1671849816,32),
    to_unsigned(1671979028,32),
    to_unsigned(1672108225,32),
    to_unsigned(1672237407,32),
    to_unsigned(1672366573,32),
    to_unsigned(1672495724,32),
    to_unsigned(1672624860,32),
    to_unsigned(1672753980,32),
    to_unsigned(1672883085,32),
    to_unsigned(1673012174,32),
    to_unsigned(1673141248,32),
    to_unsigned(1673270307,32),
    to_unsigned(1673399350,32),
    to_unsigned(1673528378,32),
    to_unsigned(1673657391,32),
    to_unsigned(1673786388,32),
    to_unsigned(1673915370,32),
    to_unsigned(1674044336,32),
    to_unsigned(1674173287,32),
    to_unsigned(1674302223,32),
    to_unsigned(1674431143,32),
    to_unsigned(1674560048,32),
    to_unsigned(1674688937,32),
    to_unsigned(1674817811,32),
    to_unsigned(1674946670,32),
    to_unsigned(1675075513,32),
    to_unsigned(1675204341,32),
    to_unsigned(1675333154,32),
    to_unsigned(1675461951,32),
    to_unsigned(1675590732,32),
    to_unsigned(1675719499,32),
    to_unsigned(1675848249,32),
    to_unsigned(1675976985,32),
    to_unsigned(1676105705,32),
    to_unsigned(1676234410,32),
    to_unsigned(1676363099,32),
    to_unsigned(1676491773,32),
    to_unsigned(1676620431,32),
    to_unsigned(1676749074,32),
    to_unsigned(1676877702,32),
    to_unsigned(1677006314,32),
    to_unsigned(1677134910,32),
    to_unsigned(1677263492,32),
    to_unsigned(1677392058,32),
    to_unsigned(1677520608,32),
    to_unsigned(1677649143,32),
    to_unsigned(1677777663,32),
    to_unsigned(1677906167,32),
    to_unsigned(1678034656,32),
    to_unsigned(1678163129,32),
    to_unsigned(1678291587,32),
    to_unsigned(1678420030,32),
    to_unsigned(1678548457,32),
    to_unsigned(1678676869,32),
    to_unsigned(1678805265,32),
    to_unsigned(1678933646,32),
    to_unsigned(1679062011,32),
    to_unsigned(1679190361,32),
    to_unsigned(1679318696,32),
    to_unsigned(1679447015,32),
    to_unsigned(1679575319,32),
    to_unsigned(1679703607,32),
    to_unsigned(1679831880,32),
    to_unsigned(1679960137,32),
    to_unsigned(1680088379,32),
    to_unsigned(1680216605,32),
    to_unsigned(1680344816,32),
    to_unsigned(1680473012,32),
    to_unsigned(1680601192,32),
    to_unsigned(1680729357,32),
    to_unsigned(1680857506,32),
    to_unsigned(1680985640,32),
    to_unsigned(1681113758,32),
    to_unsigned(1681241861,32),
    to_unsigned(1681369948,32),
    to_unsigned(1681498020,32),
    to_unsigned(1681626077,32),
    to_unsigned(1681754118,32),
    to_unsigned(1681882143,32),
    to_unsigned(1682010153,32),
    to_unsigned(1682138148,32),
    to_unsigned(1682266127,32),
    to_unsigned(1682394091,32),
    to_unsigned(1682522039,32),
    to_unsigned(1682649972,32),
    to_unsigned(1682777889,32),
    to_unsigned(1682905791,32),
    to_unsigned(1683033678,32),
    to_unsigned(1683161549,32),
    to_unsigned(1683289404,32),
    to_unsigned(1683417244,32),
    to_unsigned(1683545069,32),
    to_unsigned(1683672878,32),
    to_unsigned(1683800671,32),
    to_unsigned(1683928449,32),
    to_unsigned(1684056212,32),
    to_unsigned(1684183959,32),
    to_unsigned(1684311691,32),
    to_unsigned(1684439407,32),
    to_unsigned(1684567108,32),
    to_unsigned(1684694793,32),
    to_unsigned(1684822463,32),
    to_unsigned(1684950117,32),
    to_unsigned(1685077756,32),
    to_unsigned(1685205379,32),
    to_unsigned(1685332987,32),
    to_unsigned(1685460579,32),
    to_unsigned(1685588156,32),
    to_unsigned(1685715717,32),
    to_unsigned(1685843263,32),
    to_unsigned(1685970793,32),
    to_unsigned(1686098308,32),
    to_unsigned(1686225807,32),
    to_unsigned(1686353291,32),
    to_unsigned(1686480759,32),
    to_unsigned(1686608212,32),
    to_unsigned(1686735649,32),
    to_unsigned(1686863071,32),
    to_unsigned(1686990477,32),
    to_unsigned(1687117868,32),
    to_unsigned(1687245243,32),
    to_unsigned(1687372603,32),
    to_unsigned(1687499947,32),
    to_unsigned(1687627276,32),
    to_unsigned(1687754589,32),
    to_unsigned(1687881887,32),
    to_unsigned(1688009169,32),
    to_unsigned(1688136436,32),
    to_unsigned(1688263687,32),
    to_unsigned(1688390923,32),
    to_unsigned(1688518143,32),
    to_unsigned(1688645348,32),
    to_unsigned(1688772537,32),
    to_unsigned(1688899710,32),
    to_unsigned(1689026868,32),
    to_unsigned(1689154011,32),
    to_unsigned(1689281138,32),
    to_unsigned(1689408249,32),
    to_unsigned(1689535345,32),
    to_unsigned(1689662426,32),
    to_unsigned(1689789491,32),
    to_unsigned(1689916540,32),
    to_unsigned(1690043574,32),
    to_unsigned(1690170592,32),
    to_unsigned(1690297595,32),
    to_unsigned(1690424582,32),
    to_unsigned(1690551554,32),
    to_unsigned(1690678510,32),
    to_unsigned(1690805450,32),
    to_unsigned(1690932375,32),
    to_unsigned(1691059285,32),
    to_unsigned(1691186179,32),
    to_unsigned(1691313057,32),
    to_unsigned(1691439920,32),
    to_unsigned(1691566767,32),
    to_unsigned(1691693599,32),
    to_unsigned(1691820415,32),
    to_unsigned(1691947216,32),
    to_unsigned(1692074001,32),
    to_unsigned(1692200771,32),
    to_unsigned(1692327525,32),
    to_unsigned(1692454263,32),
    to_unsigned(1692580986,32),
    to_unsigned(1692707693,32),
    to_unsigned(1692834385,32),
    to_unsigned(1692961061,32),
    to_unsigned(1693087722,32),
    to_unsigned(1693214367,32),
    to_unsigned(1693340997,32),
    to_unsigned(1693467611,32),
    to_unsigned(1693594209,32),
    to_unsigned(1693720792,32),
    to_unsigned(1693847359,32),
    to_unsigned(1693973911,32),
    to_unsigned(1694100447,32),
    to_unsigned(1694226968,32),
    to_unsigned(1694353473,32),
    to_unsigned(1694479962,32),
    to_unsigned(1694606436,32),
    to_unsigned(1694732894,32),
    to_unsigned(1694859337,32),
    to_unsigned(1694985764,32),
    to_unsigned(1695112175,32),
    to_unsigned(1695238571,32),
    to_unsigned(1695364952,32),
    to_unsigned(1695491317,32),
    to_unsigned(1695617666,32),
    to_unsigned(1695743999,32),
    to_unsigned(1695870317,32),
    to_unsigned(1695996620,32),
    to_unsigned(1696122907,32),
    to_unsigned(1696249178,32),
    to_unsigned(1696375434,32),
    to_unsigned(1696501674,32),
    to_unsigned(1696627898,32),
    to_unsigned(1696754107,32),
    to_unsigned(1696880300,32),
    to_unsigned(1697006478,32),
    to_unsigned(1697132640,32),
    to_unsigned(1697258786,32),
    to_unsigned(1697384917,32),
    to_unsigned(1697511033,32),
    to_unsigned(1697637132,32),
    to_unsigned(1697763216,32),
    to_unsigned(1697889285,32),
    to_unsigned(1698015338,32),
    to_unsigned(1698141375,32),
    to_unsigned(1698267397,32),
    to_unsigned(1698393403,32),
    to_unsigned(1698519393,32),
    to_unsigned(1698645368,32),
    to_unsigned(1698771327,32),
    to_unsigned(1698897271,32),
    to_unsigned(1699023199,32),
    to_unsigned(1699149111,32),
    to_unsigned(1699275008,32),
    to_unsigned(1699400889,32),
    to_unsigned(1699526754,32),
    to_unsigned(1699652604,32),
    to_unsigned(1699778438,32),
    to_unsigned(1699904257,32),
    to_unsigned(1700030060,32),
    to_unsigned(1700155847,32),
    to_unsigned(1700281619,32),
    to_unsigned(1700407375,32),
    to_unsigned(1700533116,32),
    to_unsigned(1700658841,32),
    to_unsigned(1700784550,32),
    to_unsigned(1700910243,32),
    to_unsigned(1701035921,32),
    to_unsigned(1701161584,32),
    to_unsigned(1701287230,32),
    to_unsigned(1701412861,32),
    to_unsigned(1701538477,32),
    to_unsigned(1701664077,32),
    to_unsigned(1701789661,32),
    to_unsigned(1701915229,32),
    to_unsigned(1702040782,32),
    to_unsigned(1702166319,32),
    to_unsigned(1702291841,32),
    to_unsigned(1702417347,32),
    to_unsigned(1702542837,32),
    to_unsigned(1702668312,32),
    to_unsigned(1702793771,32),
    to_unsigned(1702919214,32),
    to_unsigned(1703044642,32),
    to_unsigned(1703170054,32),
    to_unsigned(1703295450,32),
    to_unsigned(1703420831,32),
    to_unsigned(1703546196,32),
    to_unsigned(1703671545,32),
    to_unsigned(1703796879,32),
    to_unsigned(1703922197,32),
    to_unsigned(1704047499,32),
    to_unsigned(1704172786,32),
    to_unsigned(1704298057,32),
    to_unsigned(1704423312,32),
    to_unsigned(1704548552,32),
    to_unsigned(1704673776,32),
    to_unsigned(1704798984,32),
    to_unsigned(1704924177,32),
    to_unsigned(1705049354,32),
    to_unsigned(1705174516,32),
    to_unsigned(1705299661,32),
    to_unsigned(1705424791,32),
    to_unsigned(1705549906,32),
    to_unsigned(1705675004,32),
    to_unsigned(1705800087,32),
    to_unsigned(1705925155,32),
    to_unsigned(1706050206,32),
    to_unsigned(1706175242,32),
    to_unsigned(1706300262,32),
    to_unsigned(1706425267,32),
    to_unsigned(1706550256,32),
    to_unsigned(1706675229,32),
    to_unsigned(1706800187,32),
    to_unsigned(1706925129,32),
    to_unsigned(1707050055,32),
    to_unsigned(1707174965,32),
    to_unsigned(1707299860,32),
    to_unsigned(1707424739,32),
    to_unsigned(1707549602,32),
    to_unsigned(1707674450,32),
    to_unsigned(1707799282,32),
    to_unsigned(1707924098,32),
    to_unsigned(1708048899,32),
    to_unsigned(1708173684,32),
    to_unsigned(1708298453,32),
    to_unsigned(1708423206,32),
    to_unsigned(1708547944,32),
    to_unsigned(1708672666,32),
    to_unsigned(1708797373,32),
    to_unsigned(1708922063,32),
    to_unsigned(1709046738,32),
    to_unsigned(1709171398,32),
    to_unsigned(1709296041,32),
    to_unsigned(1709420669,32),
    to_unsigned(1709545281,32),
    to_unsigned(1709669877,32),
    to_unsigned(1709794458,32),
    to_unsigned(1709919023,32),
    to_unsigned(1710043572,32),
    to_unsigned(1710168106,32),
    to_unsigned(1710292624,32),
    to_unsigned(1710417126,32),
    to_unsigned(1710541612,32),
    to_unsigned(1710666083,32),
    to_unsigned(1710790538,32),
    to_unsigned(1710914977,32),
    to_unsigned(1711039400,32),
    to_unsigned(1711163808,32),
    to_unsigned(1711288200,32),
    to_unsigned(1711412576,32),
    to_unsigned(1711536937,32),
    to_unsigned(1711661282,32),
    to_unsigned(1711785611,32),
    to_unsigned(1711909924,32),
    to_unsigned(1712034222,32),
    to_unsigned(1712158504,32),
    to_unsigned(1712282770,32),
    to_unsigned(1712407020,32),
    to_unsigned(1712531255,32),
    to_unsigned(1712655474,32),
    to_unsigned(1712779677,32),
    to_unsigned(1712903865,32),
    to_unsigned(1713028036,32),
    to_unsigned(1713152192,32),
    to_unsigned(1713276332,32),
    to_unsigned(1713400457,32),
    to_unsigned(1713524566,32),
    to_unsigned(1713648659,32),
    to_unsigned(1713772736,32),
    to_unsigned(1713896797,32),
    to_unsigned(1714020843,32),
    to_unsigned(1714144873,32),
    to_unsigned(1714268887,32),
    to_unsigned(1714392885,32),
    to_unsigned(1714516868,32),
    to_unsigned(1714640835,32),
    to_unsigned(1714764786,32),
    to_unsigned(1714888722,32),
    to_unsigned(1715012641,32),
    to_unsigned(1715136545,32),
    to_unsigned(1715260433,32),
    to_unsigned(1715384306,32),
    to_unsigned(1715508162,32),
    to_unsigned(1715632003,32),
    to_unsigned(1715755828,32),
    to_unsigned(1715879637,32),
    to_unsigned(1716003431,32),
    to_unsigned(1716127208,32),
    to_unsigned(1716250970,32),
    to_unsigned(1716374716,32),
    to_unsigned(1716498447,32),
    to_unsigned(1716622161,32),
    to_unsigned(1716745860,32),
    to_unsigned(1716869543,32),
    to_unsigned(1716993211,32),
    to_unsigned(1717116862,32),
    to_unsigned(1717240498,32),
    to_unsigned(1717364118,32),
    to_unsigned(1717487722,32),
    to_unsigned(1717611310,32),
    to_unsigned(1717734883,32),
    to_unsigned(1717858439,32),
    to_unsigned(1717981980,32),
    to_unsigned(1718105506,32),
    to_unsigned(1718229015,32),
    to_unsigned(1718352509,32),
    to_unsigned(1718475986,32),
    to_unsigned(1718599448,32),
    to_unsigned(1718722895,32),
    to_unsigned(1718846325,32),
    to_unsigned(1718969740,32),
    to_unsigned(1719093138,32),
    to_unsigned(1719216521,32),
    to_unsigned(1719339889,32),
    to_unsigned(1719463240,32),
    to_unsigned(1719586576,32),
    to_unsigned(1719709896,32),
    to_unsigned(1719833199,32),
    to_unsigned(1719956488,32),
    to_unsigned(1720079760,32),
    to_unsigned(1720203017,32),
    to_unsigned(1720326257,32),
    to_unsigned(1720449482,32),
    to_unsigned(1720572691,32),
    to_unsigned(1720695885,32),
    to_unsigned(1720819062,32),
    to_unsigned(1720942224,32),
    to_unsigned(1721065370,32),
    to_unsigned(1721188500,32),
    to_unsigned(1721311614,32),
    to_unsigned(1721434712,32),
    to_unsigned(1721557795,32),
    to_unsigned(1721680862,32),
    to_unsigned(1721803913,32),
    to_unsigned(1721926948,32),
    to_unsigned(1722049967,32),
    to_unsigned(1722172970,32),
    to_unsigned(1722295958,32),
    to_unsigned(1722418930,32),
    to_unsigned(1722541886,32),
    to_unsigned(1722664826,32),
    to_unsigned(1722787750,32),
    to_unsigned(1722910659,32),
    to_unsigned(1723033551,32),
    to_unsigned(1723156428,32),
    to_unsigned(1723279289,32),
    to_unsigned(1723402134,32),
    to_unsigned(1723524963,32),
    to_unsigned(1723647777,32),
    to_unsigned(1723770574,32),
    to_unsigned(1723893356,32),
    to_unsigned(1724016122,32),
    to_unsigned(1724138872,32),
    to_unsigned(1724261606,32),
    to_unsigned(1724384324,32),
    to_unsigned(1724507027,32),
    to_unsigned(1724629713,32),
    to_unsigned(1724752384,32),
    to_unsigned(1724875039,32),
    to_unsigned(1724997678,32),
    to_unsigned(1725120301,32),
    to_unsigned(1725242909,32),
    to_unsigned(1725365500,32),
    to_unsigned(1725488076,32),
    to_unsigned(1725610636,32),
    to_unsigned(1725733179,32),
    to_unsigned(1725855707,32),
    to_unsigned(1725978220,32),
    to_unsigned(1726100716,32),
    to_unsigned(1726223196,32),
    to_unsigned(1726345661,32),
    to_unsigned(1726468110,32),
    to_unsigned(1726590543,32),
    to_unsigned(1726712960,32),
    to_unsigned(1726835361,32),
    to_unsigned(1726957746,32),
    to_unsigned(1727080115,32),
    to_unsigned(1727202469,32),
    to_unsigned(1727324806,32),
    to_unsigned(1727447128,32),
    to_unsigned(1727569434,32),
    to_unsigned(1727691724,32),
    to_unsigned(1727813998,32),
    to_unsigned(1727936256,32),
    to_unsigned(1728058499,32),
    to_unsigned(1728180725,32),
    to_unsigned(1728302936,32),
    to_unsigned(1728425130,32),
    to_unsigned(1728547309,32),
    to_unsigned(1728669472,32),
    to_unsigned(1728791619,32),
    to_unsigned(1728913750,32),
    to_unsigned(1729035865,32),
    to_unsigned(1729157965,32),
    to_unsigned(1729280048,32),
    to_unsigned(1729402116,32),
    to_unsigned(1729524167,32),
    to_unsigned(1729646203,32),
    to_unsigned(1729768223,32),
    to_unsigned(1729890227,32),
    to_unsigned(1730012215,32),
    to_unsigned(1730134187,32),
    to_unsigned(1730256143,32),
    to_unsigned(1730378084,32),
    to_unsigned(1730500008,32),
    to_unsigned(1730621917,32),
    to_unsigned(1730743809,32),
    to_unsigned(1730865686,32),
    to_unsigned(1730987547,32),
    to_unsigned(1731109392,32),
    to_unsigned(1731231221,32),
    to_unsigned(1731353034,32),
    to_unsigned(1731474831,32),
    to_unsigned(1731596612,32),
    to_unsigned(1731718377,32),
    to_unsigned(1731840127,32),
    to_unsigned(1731961860,32),
    to_unsigned(1732083578,32),
    to_unsigned(1732205280,32),
    to_unsigned(1732326965,32),
    to_unsigned(1732448635,32),
    to_unsigned(1732570289,32),
    to_unsigned(1732691927,32),
    to_unsigned(1732813549,32),
    to_unsigned(1732935155,32),
    to_unsigned(1733056745,32),
    to_unsigned(1733178319,32),
    to_unsigned(1733299878,32),
    to_unsigned(1733421420,32),
    to_unsigned(1733542947,32),
    to_unsigned(1733664457,32),
    to_unsigned(1733785952,32),
    to_unsigned(1733907430,32),
    to_unsigned(1734028893,32),
    to_unsigned(1734150340,32),
    to_unsigned(1734271771,32),
    to_unsigned(1734393185,32),
    to_unsigned(1734514584,32),
    to_unsigned(1734635967,32),
    to_unsigned(1734757334,32),
    to_unsigned(1734878685,32),
    to_unsigned(1735000021,32),
    to_unsigned(1735121340,32),
    to_unsigned(1735242643,32),
    to_unsigned(1735363930,32),
    to_unsigned(1735485202,32),
    to_unsigned(1735606457,32),
    to_unsigned(1735727697,32),
    to_unsigned(1735848920,32),
    to_unsigned(1735970128,32),
    to_unsigned(1736091319,32),
    to_unsigned(1736212495,32),
    to_unsigned(1736333655,32),
    to_unsigned(1736454798,32),
    to_unsigned(1736575926,32),
    to_unsigned(1736697038,32),
    to_unsigned(1736818134,32),
    to_unsigned(1736939213,32),
    to_unsigned(1737060277,32),
    to_unsigned(1737181325,32),
    to_unsigned(1737302357,32),
    to_unsigned(1737423373,32),
    to_unsigned(1737544373,32),
    to_unsigned(1737665357,32),
    to_unsigned(1737786325,32),
    to_unsigned(1737907277,32),
    to_unsigned(1738028214,32),
    to_unsigned(1738149134,32),
    to_unsigned(1738270038,32),
    to_unsigned(1738390926,32),
    to_unsigned(1738511798,32),
    to_unsigned(1738632655,32),
    to_unsigned(1738753495,32),
    to_unsigned(1738874319,32),
    to_unsigned(1738995127,32),
    to_unsigned(1739115920,32),
    to_unsigned(1739236696,32),
    to_unsigned(1739357456,32),
    to_unsigned(1739478201,32),
    to_unsigned(1739598929,32),
    to_unsigned(1739719641,32),
    to_unsigned(1739840338,32),
    to_unsigned(1739961018,32),
    to_unsigned(1740081683,32),
    to_unsigned(1740202331,32),
    to_unsigned(1740322963,32),
    to_unsigned(1740443580,32),
    to_unsigned(1740564180,32),
    to_unsigned(1740684765,32),
    to_unsigned(1740805333,32),
    to_unsigned(1740925885,32),
    to_unsigned(1741046422,32),
    to_unsigned(1741166942,32),
    to_unsigned(1741287447,32),
    to_unsigned(1741407935,32),
    to_unsigned(1741528407,32),
    to_unsigned(1741648864,32),
    to_unsigned(1741769304,32),
    to_unsigned(1741889729,32),
    to_unsigned(1742010137,32),
    to_unsigned(1742130529,32),
    to_unsigned(1742250906,32),
    to_unsigned(1742371266,32),
    to_unsigned(1742491610,32),
    to_unsigned(1742611938,32),
    to_unsigned(1742732251,32),
    to_unsigned(1742852547,32),
    to_unsigned(1742972827,32),
    to_unsigned(1743093091,32),
    to_unsigned(1743213340,32),
    to_unsigned(1743333572,32),
    to_unsigned(1743453788,32),
    to_unsigned(1743573988,32),
    to_unsigned(1743694172,32),
    to_unsigned(1743814340,32),
    to_unsigned(1743934492,32),
    to_unsigned(1744054628,32),
    to_unsigned(1744174748,32),
    to_unsigned(1744294852,32),
    to_unsigned(1744414940,32),
    to_unsigned(1744535012,32),
    to_unsigned(1744655068,32),
    to_unsigned(1744775107,32),
    to_unsigned(1744895131,32),
    to_unsigned(1745015139,32),
    to_unsigned(1745135130,32),
    to_unsigned(1745255106,32),
    to_unsigned(1745375066,32),
    to_unsigned(1745495009,32),
    to_unsigned(1745614937,32),
    to_unsigned(1745734848,32),
    to_unsigned(1745854744,32),
    to_unsigned(1745974623,32),
    to_unsigned(1746094486,32),
    to_unsigned(1746214334,32),
    to_unsigned(1746334165,32),
    to_unsigned(1746453980,32),
    to_unsigned(1746573779,32),
    to_unsigned(1746693562,32),
    to_unsigned(1746813329,32),
    to_unsigned(1746933080,32),
    to_unsigned(1747052815,32),
    to_unsigned(1747172534,32),
    to_unsigned(1747292236,32),
    to_unsigned(1747411923,32),
    to_unsigned(1747531594,32),
    to_unsigned(1747651248,32),
    to_unsigned(1747770887,32),
    to_unsigned(1747890509,32),
    to_unsigned(1748010116,32),
    to_unsigned(1748129706,32),
    to_unsigned(1748249280,32),
    to_unsigned(1748368839,32),
    to_unsigned(1748488381,32),
    to_unsigned(1748607907,32),
    to_unsigned(1748727417,32),
    to_unsigned(1748846911,32),
    to_unsigned(1748966388,32),
    to_unsigned(1749085850,32),
    to_unsigned(1749205296,32),
    to_unsigned(1749324725,32),
    to_unsigned(1749444139,32),
    to_unsigned(1749563536,32),
    to_unsigned(1749682918,32),
    to_unsigned(1749802283,32),
    to_unsigned(1749921632,32),
    to_unsigned(1750040965,32),
    to_unsigned(1750160282,32),
    to_unsigned(1750279583,32),
    to_unsigned(1750398868,32),
    to_unsigned(1750518137,32),
    to_unsigned(1750637389,32),
    to_unsigned(1750756626,32),
    to_unsigned(1750875846,32),
    to_unsigned(1750995051,32),
    to_unsigned(1751114239,32),
    to_unsigned(1751233411,32),
    to_unsigned(1751352567,32),
    to_unsigned(1751471707,32),
    to_unsigned(1751590831,32),
    to_unsigned(1751709939,32),
    to_unsigned(1751829031,32),
    to_unsigned(1751948106,32),
    to_unsigned(1752067166,32),
    to_unsigned(1752186209,32),
    to_unsigned(1752305236,32),
    to_unsigned(1752424247,32),
    to_unsigned(1752543243,32),
    to_unsigned(1752662221,32),
    to_unsigned(1752781184,32),
    to_unsigned(1752900131,32),
    to_unsigned(1753019062,32),
    to_unsigned(1753137976,32),
    to_unsigned(1753256875,32),
    to_unsigned(1753375757,32),
    to_unsigned(1753494623,32),
    to_unsigned(1753613473,32),
    to_unsigned(1753732307,32),
    to_unsigned(1753851125,32),
    to_unsigned(1753969926,32),
    to_unsigned(1754088712,32),
    to_unsigned(1754207481,32),
    to_unsigned(1754326235,32),
    to_unsigned(1754444972,32),
    to_unsigned(1754563693,32),
    to_unsigned(1754682398,32),
    to_unsigned(1754801087,32),
    to_unsigned(1754919759,32),
    to_unsigned(1755038416,32),
    to_unsigned(1755157056,32),
    to_unsigned(1755275681,32),
    to_unsigned(1755394289,32),
    to_unsigned(1755512881,32),
    to_unsigned(1755631457,32),
    to_unsigned(1755750016,32),
    to_unsigned(1755868560,32),
    to_unsigned(1755987087,32),
    to_unsigned(1756105599,32),
    to_unsigned(1756224094,32),
    to_unsigned(1756342573,32),
    to_unsigned(1756461036,32),
    to_unsigned(1756579482,32),
    to_unsigned(1756697913,32),
    to_unsigned(1756816327,32),
    to_unsigned(1756934726,32),
    to_unsigned(1757053108,32),
    to_unsigned(1757171474,32),
    to_unsigned(1757289824,32),
    to_unsigned(1757408157,32),
    to_unsigned(1757526475,32),
    to_unsigned(1757644776,32),
    to_unsigned(1757763062,32),
    to_unsigned(1757881331,32),
    to_unsigned(1757999584,32),
    to_unsigned(1758117820,32),
    to_unsigned(1758236041,32),
    to_unsigned(1758354245,32),
    to_unsigned(1758472434,32),
    to_unsigned(1758590606,32),
    to_unsigned(1758708762,32),
    to_unsigned(1758826901,32),
    to_unsigned(1758945025,32),
    to_unsigned(1759063133,32),
    to_unsigned(1759181224,32),
    to_unsigned(1759299299,32),
    to_unsigned(1759417358,32),
    to_unsigned(1759535401,32),
    to_unsigned(1759653427,32),
    to_unsigned(1759771438,32),
    to_unsigned(1759889432,32),
    to_unsigned(1760007410,32),
    to_unsigned(1760125372,32),
    to_unsigned(1760243317,32),
    to_unsigned(1760361247,32),
    to_unsigned(1760479160,32),
    to_unsigned(1760597057,32),
    to_unsigned(1760714938,32),
    to_unsigned(1760832803,32),
    to_unsigned(1760950652,32),
    to_unsigned(1761068484,32),
    to_unsigned(1761186301,32),
    to_unsigned(1761304101,32),
    to_unsigned(1761421884,32),
    to_unsigned(1761539652,32),
    to_unsigned(1761657404,32),
    to_unsigned(1761775139,32),
    to_unsigned(1761892858,32),
    to_unsigned(1762010561,32),
    to_unsigned(1762128248,32),
    to_unsigned(1762245918,32),
    to_unsigned(1762363572,32),
    to_unsigned(1762481210,32),
    to_unsigned(1762598832,32),
    to_unsigned(1762716438,32),
    to_unsigned(1762834028,32),
    to_unsigned(1762951601,32),
    to_unsigned(1763069158,32),
    to_unsigned(1763186699,32),
    to_unsigned(1763304223,32),
    to_unsigned(1763421732,32),
    to_unsigned(1763539224,32),
    to_unsigned(1763656700,32),
    to_unsigned(1763774160,32),
    to_unsigned(1763891604,32),
    to_unsigned(1764009031,32),
    to_unsigned(1764126442,32),
    to_unsigned(1764243837,32),
    to_unsigned(1764361216,32),
    to_unsigned(1764478579,32),
    to_unsigned(1764595925,32),
    to_unsigned(1764713255,32),
    to_unsigned(1764830569,32),
    to_unsigned(1764947867,32),
    to_unsigned(1765065148,32),
    to_unsigned(1765182413,32),
    to_unsigned(1765299662,32),
    to_unsigned(1765416895,32),
    to_unsigned(1765534112,32),
    to_unsigned(1765651312,32),
    to_unsigned(1765768496,32),
    to_unsigned(1765885664,32),
    to_unsigned(1766002815,32),
    to_unsigned(1766119951,32),
    to_unsigned(1766237070,32),
    to_unsigned(1766354173,32),
    to_unsigned(1766471260,32),
    to_unsigned(1766588330,32),
    to_unsigned(1766705384,32),
    to_unsigned(1766822422,32),
    to_unsigned(1766939444,32),
    to_unsigned(1767056449,32),
    to_unsigned(1767173439,32),
    to_unsigned(1767290412,32),
    to_unsigned(1767407368,32),
    to_unsigned(1767524309,32),
    to_unsigned(1767641233,32),
    to_unsigned(1767758141,32),
    to_unsigned(1767875033,32),
    to_unsigned(1767991909,32),
    to_unsigned(1768108768,32),
    to_unsigned(1768225611,32),
    to_unsigned(1768342438,32),
    to_unsigned(1768459248,32),
    to_unsigned(1768576042,32),
    to_unsigned(1768692820,32),
    to_unsigned(1768809582,32),
    to_unsigned(1768926328,32),
    to_unsigned(1769043057,32),
    to_unsigned(1769159770,32),
    to_unsigned(1769276466,32),
    to_unsigned(1769393147,32),
    to_unsigned(1769509811,32),
    to_unsigned(1769626459,32),
    to_unsigned(1769743091,32),
    to_unsigned(1769859706,32),
    to_unsigned(1769976305,32),
    to_unsigned(1770092888,32),
    to_unsigned(1770209454,32),
    to_unsigned(1770326005,32),
    to_unsigned(1770442539,32),
    to_unsigned(1770559057,32),
    to_unsigned(1770675558,32),
    to_unsigned(1770792043,32),
    to_unsigned(1770908512,32),
    to_unsigned(1771024965,32),
    to_unsigned(1771141401,32),
    to_unsigned(1771257821,32),
    to_unsigned(1771374225,32),
    to_unsigned(1771490613,32),
    to_unsigned(1771606984,32),
    to_unsigned(1771723339,32),
    to_unsigned(1771839677,32),
    to_unsigned(1771956000,32),
    to_unsigned(1772072306,32),
    to_unsigned(1772188596,32),
    to_unsigned(1772304869,32),
    to_unsigned(1772421126,32),
    to_unsigned(1772537367,32),
    to_unsigned(1772653592,32),
    to_unsigned(1772769800,32),
    to_unsigned(1772885992,32),
    to_unsigned(1773002168,32),
    to_unsigned(1773118328,32),
    to_unsigned(1773234471,32),
    to_unsigned(1773350598,32),
    to_unsigned(1773466708,32),
    to_unsigned(1773582803,32),
    to_unsigned(1773698880,32),
    to_unsigned(1773814942,32),
    to_unsigned(1773930987,32),
    to_unsigned(1774047017,32),
    to_unsigned(1774163029,32),
    to_unsigned(1774279026,32),
    to_unsigned(1774395006,32),
    to_unsigned(1774510970,32),
    to_unsigned(1774626917,32),
    to_unsigned(1774742848,32),
    to_unsigned(1774858763,32),
    to_unsigned(1774974662,32),
    to_unsigned(1775090544,32),
    to_unsigned(1775206410,32),
    to_unsigned(1775322260,32),
    to_unsigned(1775438093,32),
    to_unsigned(1775553910,32),
    to_unsigned(1775669710,32),
    to_unsigned(1775785495,32),
    to_unsigned(1775901263,32),
    to_unsigned(1776017015,32),
    to_unsigned(1776132750,32),
    to_unsigned(1776248469,32),
    to_unsigned(1776364172,32),
    to_unsigned(1776479858,32),
    to_unsigned(1776595528,32),
    to_unsigned(1776711182,32),
    to_unsigned(1776826819,32),
    to_unsigned(1776942440,32),
    to_unsigned(1777058045,32),
    to_unsigned(1777173633,32),
    to_unsigned(1777289205,32),
    to_unsigned(1777404761,32),
    to_unsigned(1777520301,32),
    to_unsigned(1777635824,32),
    to_unsigned(1777751330,32),
    to_unsigned(1777866821,32),
    to_unsigned(1777982295,32),
    to_unsigned(1778097752,32),
    to_unsigned(1778213194,32),
    to_unsigned(1778328619,32),
    to_unsigned(1778444027,32),
    to_unsigned(1778559420,32),
    to_unsigned(1778674796,32),
    to_unsigned(1778790155,32),
    to_unsigned(1778905498,32),
    to_unsigned(1779020825,32),
    to_unsigned(1779136136,32),
    to_unsigned(1779251430,32),
    to_unsigned(1779366708,32),
    to_unsigned(1779481969,32),
    to_unsigned(1779597214,32),
    to_unsigned(1779712443,32),
    to_unsigned(1779827656,32),
    to_unsigned(1779942852,32),
    to_unsigned(1780058031,32),
    to_unsigned(1780173195,32),
    to_unsigned(1780288342,32),
    to_unsigned(1780403472,32),
    to_unsigned(1780518587,32),
    to_unsigned(1780633684,32),
    to_unsigned(1780748766,32),
    to_unsigned(1780863831,32),
    to_unsigned(1780978880,32),
    to_unsigned(1781093912,32),
    to_unsigned(1781208928,32),
    to_unsigned(1781323928,32),
    to_unsigned(1781438911,32),
    to_unsigned(1781553878,32),
    to_unsigned(1781668829,32),
    to_unsigned(1781783763,32),
    to_unsigned(1781898680,32),
    to_unsigned(1782013582,32),
    to_unsigned(1782128467,32),
    to_unsigned(1782243336,32),
    to_unsigned(1782358188,32),
    to_unsigned(1782473024,32),
    to_unsigned(1782587843,32),
    to_unsigned(1782702646,32),
    to_unsigned(1782817433,32),
    to_unsigned(1782932203,32),
    to_unsigned(1783046957,32),
    to_unsigned(1783161695,32),
    to_unsigned(1783276416,32),
    to_unsigned(1783391121,32),
    to_unsigned(1783505809,32),
    to_unsigned(1783620481,32),
    to_unsigned(1783735137,32),
    to_unsigned(1783849776,32),
    to_unsigned(1783964399,32),
    to_unsigned(1784079005,32),
    to_unsigned(1784193595,32),
    to_unsigned(1784308169,32),
    to_unsigned(1784422726,32),
    to_unsigned(1784537267,32),
    to_unsigned(1784651791,32),
    to_unsigned(1784766299,32),
    to_unsigned(1784880790,32),
    to_unsigned(1784995266,32),
    to_unsigned(1785109724,32),
    to_unsigned(1785224167,32),
    to_unsigned(1785338593,32),
    to_unsigned(1785453002,32),
    to_unsigned(1785567395,32),
    to_unsigned(1785681772,32),
    to_unsigned(1785796132,32),
    to_unsigned(1785910476,32),
    to_unsigned(1786024804,32),
    to_unsigned(1786139115,32),
    to_unsigned(1786253409,32),
    to_unsigned(1786367688,32),
    to_unsigned(1786481949,32),
    to_unsigned(1786596195,32),
    to_unsigned(1786710424,32),
    to_unsigned(1786824636,32),
    to_unsigned(1786938832,32),
    to_unsigned(1787053012,32),
    to_unsigned(1787167175,32),
    to_unsigned(1787281322,32),
    to_unsigned(1787395453,32),
    to_unsigned(1787509567,32),
    to_unsigned(1787623664,32),
    to_unsigned(1787737745,32),
    to_unsigned(1787851810,32),
    to_unsigned(1787965858,32),
    to_unsigned(1788079890,32),
    to_unsigned(1788193905,32),
    to_unsigned(1788307904,32),
    to_unsigned(1788421887,32),
    to_unsigned(1788535853,32),
    to_unsigned(1788649802,32),
    to_unsigned(1788763736,32),
    to_unsigned(1788877652,32),
    to_unsigned(1788991553,32),
    to_unsigned(1789105436,32),
    to_unsigned(1789219304,32),
    to_unsigned(1789333155,32),
    to_unsigned(1789446989,32),
    to_unsigned(1789560807,32),
    to_unsigned(1789674609,32),
    to_unsigned(1789788394,32),
    to_unsigned(1789902163,32),
    to_unsigned(1790015915,32),
    to_unsigned(1790129651,32),
    to_unsigned(1790243370,32),
    to_unsigned(1790357073,32),
    to_unsigned(1790470760,32),
    to_unsigned(1790584430,32),
    to_unsigned(1790698083,32),
    to_unsigned(1790811720,32),
    to_unsigned(1790925341,32),
    to_unsigned(1791038945,32),
    to_unsigned(1791152533,32),
    to_unsigned(1791266104,32),
    to_unsigned(1791379659,32),
    to_unsigned(1791493197,32),
    to_unsigned(1791606719,32),
    to_unsigned(1791720224,32),
    to_unsigned(1791833713,32),
    to_unsigned(1791947185,32),
    to_unsigned(1792060641,32),
    to_unsigned(1792174081,32),
    to_unsigned(1792287504,32),
    to_unsigned(1792400910,32),
    to_unsigned(1792514300,32),
    to_unsigned(1792627674,32),
    to_unsigned(1792741031,32),
    to_unsigned(1792854372,32),
    to_unsigned(1792967696,32),
    to_unsigned(1793081003,32),
    to_unsigned(1793194294,32),
    to_unsigned(1793307569,32),
    to_unsigned(1793420827,32),
    to_unsigned(1793534069,32),
    to_unsigned(1793647294,32),
    to_unsigned(1793760503,32),
    to_unsigned(1793873695,32),
    to_unsigned(1793986871,32),
    to_unsigned(1794100030,32),
    to_unsigned(1794213173,32),
    to_unsigned(1794326299,32),
    to_unsigned(1794439409,32),
    to_unsigned(1794552503,32),
    to_unsigned(1794665579,32),
    to_unsigned(1794778640,32),
    to_unsigned(1794891683,32),
    to_unsigned(1795004711,32),
    to_unsigned(1795117722,32),
    to_unsigned(1795230716,32),
    to_unsigned(1795343694,32),
    to_unsigned(1795456655,32),
    to_unsigned(1795569600,32),
    to_unsigned(1795682528,32),
    to_unsigned(1795795440,32),
    to_unsigned(1795908335,32),
    to_unsigned(1796021214,32),
    to_unsigned(1796134076,32),
    to_unsigned(1796246922,32),
    to_unsigned(1796359751,32),
    to_unsigned(1796472564,32),
    to_unsigned(1796585360,32),
    to_unsigned(1796698140,32),
    to_unsigned(1796810903,32),
    to_unsigned(1796923650,32),
    to_unsigned(1797036380,32),
    to_unsigned(1797149094,32),
    to_unsigned(1797261791,32),
    to_unsigned(1797374472,32),
    to_unsigned(1797487136,32),
    to_unsigned(1797599783,32),
    to_unsigned(1797712414,32),
    to_unsigned(1797825029,32),
    to_unsigned(1797937627,32),
    to_unsigned(1798050208,32),
    to_unsigned(1798162773,32),
    to_unsigned(1798275322,32),
    to_unsigned(1798387854,32),
    to_unsigned(1798500369,32),
    to_unsigned(1798612868,32),
    to_unsigned(1798725350,32),
    to_unsigned(1798837816,32),
    to_unsigned(1798950265,32),
    to_unsigned(1799062698,32),
    to_unsigned(1799175114,32),
    to_unsigned(1799287514,32),
    to_unsigned(1799399897,32),
    to_unsigned(1799512263,32),
    to_unsigned(1799624613,32),
    to_unsigned(1799736947,32),
    to_unsigned(1799849263,32),
    to_unsigned(1799961564,32),
    to_unsigned(1800073848,32),
    to_unsigned(1800186115,32),
    to_unsigned(1800298366,32),
    to_unsigned(1800410600,32),
    to_unsigned(1800522818,32),
    to_unsigned(1800635019,32),
    to_unsigned(1800747203,32),
    to_unsigned(1800859371,32),
    to_unsigned(1800971523,32),
    to_unsigned(1801083657,32),
    to_unsigned(1801195776,32),
    to_unsigned(1801307878,32),
    to_unsigned(1801419963,32),
    to_unsigned(1801532031,32),
    to_unsigned(1801644083,32),
    to_unsigned(1801756119,32),
    to_unsigned(1801868138,32),
    to_unsigned(1801980140,32),
    to_unsigned(1802092126,32),
    to_unsigned(1802204095,32),
    to_unsigned(1802316048,32),
    to_unsigned(1802427984,32),
    to_unsigned(1802539904,32),
    to_unsigned(1802651807,32),
    to_unsigned(1802763693,32),
    to_unsigned(1802875563,32),
    to_unsigned(1802987417,32),
    to_unsigned(1803099253,32),
    to_unsigned(1803211073,32),
    to_unsigned(1803322877,32),
    to_unsigned(1803434664,32),
    to_unsigned(1803546434,32),
    to_unsigned(1803658188,32),
    to_unsigned(1803769926,32),
    to_unsigned(1803881646,32),
    to_unsigned(1803993350,32),
    to_unsigned(1804105038,32),
    to_unsigned(1804216709,32),
    to_unsigned(1804328363,32),
    to_unsigned(1804440001,32),
    to_unsigned(1804551622,32),
    to_unsigned(1804663227,32),
    to_unsigned(1804774815,32),
    to_unsigned(1804886386,32),
    to_unsigned(1804997941,32),
    to_unsigned(1805109479,32),
    to_unsigned(1805221001,32),
    to_unsigned(1805332506,32),
    to_unsigned(1805443994,32),
    to_unsigned(1805555466,32),
    to_unsigned(1805666922,32),
    to_unsigned(1805778360,32),
    to_unsigned(1805889782,32),
    to_unsigned(1806001188,32),
    to_unsigned(1806112577,32),
    to_unsigned(1806223949,32),
    to_unsigned(1806335305,32),
    to_unsigned(1806446644,32),
    to_unsigned(1806557966,32),
    to_unsigned(1806669272,32),
    to_unsigned(1806780561,32),
    to_unsigned(1806891834,32),
    to_unsigned(1807003090,32),
    to_unsigned(1807114329,32),
    to_unsigned(1807225552,32),
    to_unsigned(1807336758,32),
    to_unsigned(1807447948,32),
    to_unsigned(1807559121,32),
    to_unsigned(1807670277,32),
    to_unsigned(1807781417,32),
    to_unsigned(1807892540,32),
    to_unsigned(1808003647,32),
    to_unsigned(1808114737,32),
    to_unsigned(1808225810,32),
    to_unsigned(1808336866,32),
    to_unsigned(1808447906,32),
    to_unsigned(1808558930,32),
    to_unsigned(1808669937,32),
    to_unsigned(1808780927,32),
    to_unsigned(1808891900,32),
    to_unsigned(1809002857,32),
    to_unsigned(1809113798,32),
    to_unsigned(1809224721,32),
    to_unsigned(1809335628,32),
    to_unsigned(1809446519,32),
    to_unsigned(1809557392,32),
    to_unsigned(1809668249,32),
    to_unsigned(1809779090,32),
    to_unsigned(1809889914,32),
    to_unsigned(1810000721,32),
    to_unsigned(1810111512,32),
    to_unsigned(1810222286,32),
    to_unsigned(1810333043,32),
    to_unsigned(1810443784,32),
    to_unsigned(1810554508,32),
    to_unsigned(1810665215,32),
    to_unsigned(1810775906,32),
    to_unsigned(1810886580,32),
    to_unsigned(1810997237,32),
    to_unsigned(1811107878,32),
    to_unsigned(1811218502,32),
    to_unsigned(1811329110,32),
    to_unsigned(1811439700,32),
    to_unsigned(1811550275,32),
    to_unsigned(1811660832,32),
    to_unsigned(1811771373,32),
    to_unsigned(1811881897,32),
    to_unsigned(1811992405,32),
    to_unsigned(1812102896,32),
    to_unsigned(1812213370,32),
    to_unsigned(1812323828,32),
    to_unsigned(1812434269,32),
    to_unsigned(1812544693,32),
    to_unsigned(1812655101,32),
    to_unsigned(1812765492,32),
    to_unsigned(1812875866,32),
    to_unsigned(1812986224,32),
    to_unsigned(1813096565,32),
    to_unsigned(1813206889,32),
    to_unsigned(1813317197,32),
    to_unsigned(1813427488,32),
    to_unsigned(1813537762,32),
    to_unsigned(1813648020,32),
    to_unsigned(1813758261,32),
    to_unsigned(1813868485,32),
    to_unsigned(1813978693,32),
    to_unsigned(1814088884,32),
    to_unsigned(1814199058,32),
    to_unsigned(1814309215,32),
    to_unsigned(1814419356,32),
    to_unsigned(1814529481,32),
    to_unsigned(1814639588,32),
    to_unsigned(1814749679,32),
    to_unsigned(1814859753,32),
    to_unsigned(1814969811,32),
    to_unsigned(1815079852,32),
    to_unsigned(1815189876,32),
    to_unsigned(1815299883,32),
    to_unsigned(1815409874,32),
    to_unsigned(1815519848,32),
    to_unsigned(1815629806,32),
    to_unsigned(1815739747,32),
    to_unsigned(1815849671,32),
    to_unsigned(1815959578,32),
    to_unsigned(1816069469,32),
    to_unsigned(1816179343,32),
    to_unsigned(1816289200,32),
    to_unsigned(1816399040,32),
    to_unsigned(1816508864,32),
    to_unsigned(1816618672,32),
    to_unsigned(1816728462,32),
    to_unsigned(1816838236,32),
    to_unsigned(1816947993,32),
    to_unsigned(1817057733,32),
    to_unsigned(1817167457,32),
    to_unsigned(1817277164,32),
    to_unsigned(1817386854,32),
    to_unsigned(1817496528,32),
    to_unsigned(1817606185,32),
    to_unsigned(1817715825,32),
    to_unsigned(1817825448,32),
    to_unsigned(1817935055,32),
    to_unsigned(1818044645,32),
    to_unsigned(1818154218,32),
    to_unsigned(1818263775,32),
    to_unsigned(1818373315,32),
    to_unsigned(1818482838,32),
    to_unsigned(1818592345,32),
    to_unsigned(1818701834,32),
    to_unsigned(1818811307,32),
    to_unsigned(1818920764,32),
    to_unsigned(1819030203,32),
    to_unsigned(1819139626,32),
    to_unsigned(1819249032,32),
    to_unsigned(1819358422,32),
    to_unsigned(1819467795,32),
    to_unsigned(1819577151,32),
    to_unsigned(1819686490,32),
    to_unsigned(1819795812,32),
    to_unsigned(1819905118,32),
    to_unsigned(1820014407,32),
    to_unsigned(1820123680,32),
    to_unsigned(1820232935,32),
    to_unsigned(1820342174,32),
    to_unsigned(1820451396,32),
    to_unsigned(1820560602,32),
    to_unsigned(1820669790,32),
    to_unsigned(1820778962,32),
    to_unsigned(1820888118,32),
    to_unsigned(1820997256,32),
    to_unsigned(1821106378,32),
    to_unsigned(1821215483,32),
    to_unsigned(1821324571,32),
    to_unsigned(1821433643,32),
    to_unsigned(1821542697,32),
    to_unsigned(1821651736,32),
    to_unsigned(1821760757,32),
    to_unsigned(1821869761,32),
    to_unsigned(1821978749,32),
    to_unsigned(1822087720,32),
    to_unsigned(1822196675,32),
    to_unsigned(1822305612,32),
    to_unsigned(1822414533,32),
    to_unsigned(1822523437,32),
    to_unsigned(1822632324,32),
    to_unsigned(1822741195,32),
    to_unsigned(1822850049,32),
    to_unsigned(1822958886,32),
    to_unsigned(1823067706,32),
    to_unsigned(1823176510,32),
    to_unsigned(1823285296,32),
    to_unsigned(1823394066,32),
    to_unsigned(1823502820,32),
    to_unsigned(1823611556,32),
    to_unsigned(1823720276,32),
    to_unsigned(1823828979,32),
    to_unsigned(1823937665,32),
    to_unsigned(1824046334,32),
    to_unsigned(1824154987,32),
    to_unsigned(1824263623,32),
    to_unsigned(1824372242,32),
    to_unsigned(1824480844,32),
    to_unsigned(1824589430,32),
    to_unsigned(1824697999,32),
    to_unsigned(1824806551,32),
    to_unsigned(1824915086,32),
    to_unsigned(1825023605,32),
    to_unsigned(1825132106,32),
    to_unsigned(1825240591,32),
    to_unsigned(1825349060,32),
    to_unsigned(1825457511,32),
    to_unsigned(1825565946,32),
    to_unsigned(1825674363,32),
    to_unsigned(1825782765,32),
    to_unsigned(1825891149,32),
    to_unsigned(1825999516,32),
    to_unsigned(1826107867,32),
    to_unsigned(1826216201,32),
    to_unsigned(1826324518,32),
    to_unsigned(1826432818,32),
    to_unsigned(1826541102,32),
    to_unsigned(1826649369,32),
    to_unsigned(1826757619,32),
    to_unsigned(1826865852,32),
    to_unsigned(1826974068,32),
    to_unsigned(1827082268,32),
    to_unsigned(1827190451,32),
    to_unsigned(1827298617,32),
    to_unsigned(1827406766,32),
    to_unsigned(1827514898,32),
    to_unsigned(1827623014,32),
    to_unsigned(1827731113,32),
    to_unsigned(1827839195,32),
    to_unsigned(1827947260,32),
    to_unsigned(1828055309,32),
    to_unsigned(1828163340,32),
    to_unsigned(1828271355,32),
    to_unsigned(1828379353,32),
    to_unsigned(1828487334,32),
    to_unsigned(1828595299,32),
    to_unsigned(1828703246,32),
    to_unsigned(1828811177,32),
    to_unsigned(1828919091,32),
    to_unsigned(1829026988,32),
    to_unsigned(1829134868,32),
    to_unsigned(1829242732,32),
    to_unsigned(1829350579,32),
    to_unsigned(1829458409,32),
    to_unsigned(1829566222,32),
    to_unsigned(1829674018,32),
    to_unsigned(1829781797,32),
    to_unsigned(1829889560,32),
    to_unsigned(1829997306,32),
    to_unsigned(1830105035,32),
    to_unsigned(1830212747,32),
    to_unsigned(1830320442,32),
    to_unsigned(1830428121,32),
    to_unsigned(1830535783,32),
    to_unsigned(1830643428,32),
    to_unsigned(1830751056,32),
    to_unsigned(1830858667,32),
    to_unsigned(1830966261,32),
    to_unsigned(1831073839,32),
    to_unsigned(1831181399,32),
    to_unsigned(1831288943,32),
    to_unsigned(1831396470,32),
    to_unsigned(1831503981,32),
    to_unsigned(1831611474,32),
    to_unsigned(1831718951,32),
    to_unsigned(1831826410,32),
    to_unsigned(1831933853,32),
    to_unsigned(1832041279,32),
    to_unsigned(1832148688,32),
    to_unsigned(1832256081,32),
    to_unsigned(1832363456,32),
    to_unsigned(1832470815,32),
    to_unsigned(1832578157,32),
    to_unsigned(1832685482,32),
    to_unsigned(1832792790,32),
    to_unsigned(1832900081,32),
    to_unsigned(1833007356,32),
    to_unsigned(1833114613,32),
    to_unsigned(1833221854,32),
    to_unsigned(1833329078,32),
    to_unsigned(1833436285,32),
    to_unsigned(1833543475,32),
    to_unsigned(1833650649,32),
    to_unsigned(1833757805,32),
    to_unsigned(1833864945,32),
    to_unsigned(1833972068,32),
    to_unsigned(1834079174,32),
    to_unsigned(1834186263,32),
    to_unsigned(1834293335,32),
    to_unsigned(1834400390,32),
    to_unsigned(1834507429,32),
    to_unsigned(1834614450,32),
    to_unsigned(1834721455,32),
    to_unsigned(1834828443,32),
    to_unsigned(1834935414,32),
    to_unsigned(1835042368,32),
    to_unsigned(1835149305,32),
    to_unsigned(1835256226,32),
    to_unsigned(1835363129,32),
    to_unsigned(1835470016,32),
    to_unsigned(1835576886,32),
    to_unsigned(1835683739,32),
    to_unsigned(1835790575,32),
    to_unsigned(1835897394,32),
    to_unsigned(1836004196,32),
    to_unsigned(1836110982,32),
    to_unsigned(1836217750,32),
    to_unsigned(1836324502,32),
    to_unsigned(1836431237,32),
    to_unsigned(1836537955,32),
    to_unsigned(1836644656,32),
    to_unsigned(1836751340,32),
    to_unsigned(1836858007,32),
    to_unsigned(1836964658,32),
    to_unsigned(1837071291,32),
    to_unsigned(1837177908,32),
    to_unsigned(1837284508,32),
    to_unsigned(1837391091,32),
    to_unsigned(1837497657,32),
    to_unsigned(1837604206,32),
    to_unsigned(1837710738,32),
    to_unsigned(1837817253,32),
    to_unsigned(1837923752,32),
    to_unsigned(1838030233,32),
    to_unsigned(1838136698,32),
    to_unsigned(1838243145,32),
    to_unsigned(1838349576,32),
    to_unsigned(1838455990,32),
    to_unsigned(1838562387,32),
    to_unsigned(1838668767,32),
    to_unsigned(1838775130,32),
    to_unsigned(1838881477,32),
    to_unsigned(1838987806,32),
    to_unsigned(1839094119,32),
    to_unsigned(1839200414,32),
    to_unsigned(1839306693,32),
    to_unsigned(1839412955,32),
    to_unsigned(1839519200,32),
    to_unsigned(1839625428,32),
    to_unsigned(1839731639,32),
    to_unsigned(1839837833,32),
    to_unsigned(1839944010,32),
    to_unsigned(1840050171,32),
    to_unsigned(1840156314,32),
    to_unsigned(1840262440,32),
    to_unsigned(1840368550,32),
    to_unsigned(1840474643,32),
    to_unsigned(1840580719,32),
    to_unsigned(1840686777,32),
    to_unsigned(1840792819,32),
    to_unsigned(1840898844,32),
    to_unsigned(1841004852,32),
    to_unsigned(1841110844,32),
    to_unsigned(1841216818,32),
    to_unsigned(1841322775,32),
    to_unsigned(1841428715,32),
    to_unsigned(1841534639,32),
    to_unsigned(1841640545,32),
    to_unsigned(1841746435,32),
    to_unsigned(1841852308,32),
    to_unsigned(1841958164,32),
    to_unsigned(1842064002,32),
    to_unsigned(1842169824,32),
    to_unsigned(1842275629,32),
    to_unsigned(1842381417,32),
    to_unsigned(1842487188,32),
    to_unsigned(1842592942,32),
    to_unsigned(1842698680,32),
    to_unsigned(1842804400,32),
    to_unsigned(1842910103,32),
    to_unsigned(1843015790,32),
    to_unsigned(1843121459,32),
    to_unsigned(1843227112,32),
    to_unsigned(1843332747,32),
    to_unsigned(1843438366,32),
    to_unsigned(1843543968,32),
    to_unsigned(1843649552,32),
    to_unsigned(1843755120,32),
    to_unsigned(1843860671,32),
    to_unsigned(1843966205,32),
    to_unsigned(1844071722,32),
    to_unsigned(1844177222,32),
    to_unsigned(1844282705,32),
    to_unsigned(1844388171,32),
    to_unsigned(1844493620,32),
    to_unsigned(1844599052,32),
    to_unsigned(1844704467,32),
    to_unsigned(1844809866,32),
    to_unsigned(1844915247,32),
    to_unsigned(1845020611,32),
    to_unsigned(1845125959,32),
    to_unsigned(1845231289,32),
    to_unsigned(1845336603,32),
    to_unsigned(1845441899,32),
    to_unsigned(1845547179,32),
    to_unsigned(1845652441,32),
    to_unsigned(1845757687,32),
    to_unsigned(1845862916,32),
    to_unsigned(1845968127,32),
    to_unsigned(1846073322,32),
    to_unsigned(1846178500,32),
    to_unsigned(1846283661,32),
    to_unsigned(1846388805,32),
    to_unsigned(1846493931,32),
    to_unsigned(1846599041,32),
    to_unsigned(1846704134,32),
    to_unsigned(1846809210,32),
    to_unsigned(1846914269,32),
    to_unsigned(1847019311,32),
    to_unsigned(1847124336,32),
    to_unsigned(1847229344,32),
    to_unsigned(1847334335,32),
    to_unsigned(1847439309,32),
    to_unsigned(1847544266,32),
    to_unsigned(1847649206,32),
    to_unsigned(1847754129,32),
    to_unsigned(1847859035,32),
    to_unsigned(1847963925,32),
    to_unsigned(1848068797,32),
    to_unsigned(1848173652,32),
    to_unsigned(1848278490,32),
    to_unsigned(1848383311,32),
    to_unsigned(1848488116,32),
    to_unsigned(1848592903,32),
    to_unsigned(1848697673,32),
    to_unsigned(1848802426,32),
    to_unsigned(1848907162,32),
    to_unsigned(1849011882,32),
    to_unsigned(1849116584,32),
    to_unsigned(1849221269,32),
    to_unsigned(1849325937,32),
    to_unsigned(1849430589,32),
    to_unsigned(1849535223,32),
    to_unsigned(1849639840,32),
    to_unsigned(1849744440,32),
    to_unsigned(1849849024,32),
    to_unsigned(1849953590,32),
    to_unsigned(1850058139,32),
    to_unsigned(1850162671,32),
    to_unsigned(1850267187,32),
    to_unsigned(1850371685,32),
    to_unsigned(1850476166,32),
    to_unsigned(1850580630,32),
    to_unsigned(1850685077,32),
    to_unsigned(1850789508,32),
    to_unsigned(1850893921,32),
    to_unsigned(1850998317,32),
    to_unsigned(1851102696,32),
    to_unsigned(1851207058,32),
    to_unsigned(1851311403,32),
    to_unsigned(1851415731,32),
    to_unsigned(1851520042,32),
    to_unsigned(1851624337,32),
    to_unsigned(1851728614,32),
    to_unsigned(1851832874,32),
    to_unsigned(1851937117,32),
    to_unsigned(1852041343,32),
    to_unsigned(1852145551,32),
    to_unsigned(1852249743,32),
    to_unsigned(1852353918,32),
    to_unsigned(1852458076,32),
    to_unsigned(1852562217,32),
    to_unsigned(1852666341,32),
    to_unsigned(1852770448,32),
    to_unsigned(1852874537,32),
    to_unsigned(1852978610,32),
    to_unsigned(1853082666,32),
    to_unsigned(1853186704,32),
    to_unsigned(1853290726,32),
    to_unsigned(1853394731,32),
    to_unsigned(1853498718,32),
    to_unsigned(1853602689,32),
    to_unsigned(1853706642,32),
    to_unsigned(1853810579,32),
    to_unsigned(1853914498,32),
    to_unsigned(1854018400,32),
    to_unsigned(1854122286,32),
    to_unsigned(1854226154,32),
    to_unsigned(1854330005,32),
    to_unsigned(1854433839,32),
    to_unsigned(1854537657,32),
    to_unsigned(1854641457,32),
    to_unsigned(1854745240,32),
    to_unsigned(1854849006,32),
    to_unsigned(1854952755,32),
    to_unsigned(1855056487,32),
    to_unsigned(1855160201,32),
    to_unsigned(1855263899,32),
    to_unsigned(1855367580,32),
    to_unsigned(1855471244,32),
    to_unsigned(1855574890,32),
    to_unsigned(1855678520,32),
    to_unsigned(1855782132,32),
    to_unsigned(1855885728,32),
    to_unsigned(1855989306,32),
    to_unsigned(1856092868,32),
    to_unsigned(1856196412,32),
    to_unsigned(1856299939,32),
    to_unsigned(1856403449,32),
    to_unsigned(1856506942,32),
    to_unsigned(1856610418,32),
    to_unsigned(1856713877,32),
    to_unsigned(1856817319,32),
    to_unsigned(1856920744,32),
    to_unsigned(1857024152,32),
    to_unsigned(1857127543,32),
    to_unsigned(1857230916,32),
    to_unsigned(1857334273,32),
    to_unsigned(1857437612,32),
    to_unsigned(1857540935,32),
    to_unsigned(1857644240,32),
    to_unsigned(1857747528,32),
    to_unsigned(1857850799,32),
    to_unsigned(1857954053,32),
    to_unsigned(1858057291,32),
    to_unsigned(1858160510,32),
    to_unsigned(1858263713,32),
    to_unsigned(1858366899,32),
    to_unsigned(1858470068,32),
    to_unsigned(1858573219,32),
    to_unsigned(1858676354,32),
    to_unsigned(1858779471,32),
    to_unsigned(1858882572,32),
    to_unsigned(1858985655,32),
    to_unsigned(1859088721,32),
    to_unsigned(1859191770,32),
    to_unsigned(1859294802,32),
    to_unsigned(1859397817,32),
    to_unsigned(1859500815,32),
    to_unsigned(1859603796,32),
    to_unsigned(1859706760,32),
    to_unsigned(1859809706,32),
    to_unsigned(1859912636,32),
    to_unsigned(1860015548,32),
    to_unsigned(1860118443,32),
    to_unsigned(1860221321,32),
    to_unsigned(1860324182,32),
    to_unsigned(1860427026,32),
    to_unsigned(1860529853,32),
    to_unsigned(1860632663,32),
    to_unsigned(1860735456,32),
    to_unsigned(1860838231,32),
    to_unsigned(1860940990,32),
    to_unsigned(1861043731,32),
    to_unsigned(1861146455,32),
    to_unsigned(1861249163,32),
    to_unsigned(1861351853,32),
    to_unsigned(1861454525,32),
    to_unsigned(1861557181,32),
    to_unsigned(1861659820,32),
    to_unsigned(1861762442,32),
    to_unsigned(1861865046,32),
    to_unsigned(1861967633,32),
    to_unsigned(1862070204,32),
    to_unsigned(1862172757,32),
    to_unsigned(1862275293,32),
    to_unsigned(1862377812,32),
    to_unsigned(1862480314,32),
    to_unsigned(1862582798,32),
    to_unsigned(1862685266,32),
    to_unsigned(1862787716,32),
    to_unsigned(1862890149,32),
    to_unsigned(1862992566,32),
    to_unsigned(1863094965,32),
    to_unsigned(1863197347,32),
    to_unsigned(1863299711,32),
    to_unsigned(1863402059,32),
    to_unsigned(1863504390,32),
    to_unsigned(1863606703,32),
    to_unsigned(1863708999,32),
    to_unsigned(1863811278,32),
    to_unsigned(1863913540,32),
    to_unsigned(1864015785,32),
    to_unsigned(1864118013,32),
    to_unsigned(1864220224,32),
    to_unsigned(1864322417,32),
    to_unsigned(1864424594,32),
    to_unsigned(1864526753,32),
    to_unsigned(1864628895,32),
    to_unsigned(1864731020,32),
    to_unsigned(1864833128,32),
    to_unsigned(1864935218,32),
    to_unsigned(1865037292,32),
    to_unsigned(1865139348,32),
    to_unsigned(1865241387,32),
    to_unsigned(1865343409,32),
    to_unsigned(1865445414,32),
    to_unsigned(1865547402,32),
    to_unsigned(1865649373,32),
    to_unsigned(1865751326,32),
    to_unsigned(1865853263,32),
    to_unsigned(1865955182,32),
    to_unsigned(1866057084,32),
    to_unsigned(1866158969,32),
    to_unsigned(1866260836,32),
    to_unsigned(1866362687,32),
    to_unsigned(1866464520,32),
    to_unsigned(1866566337,32),
    to_unsigned(1866668136,32),
    to_unsigned(1866769918,32),
    to_unsigned(1866871683,32),
    to_unsigned(1866973430,32),
    to_unsigned(1867075161,32),
    to_unsigned(1867176874,32),
    to_unsigned(1867278570,32),
    to_unsigned(1867380249,32),
    to_unsigned(1867481911,32),
    to_unsigned(1867583556,32),
    to_unsigned(1867685183,32),
    to_unsigned(1867786793,32),
    to_unsigned(1867888387,32),
    to_unsigned(1867989963,32),
    to_unsigned(1868091521,32),
    to_unsigned(1868193063,32),
    to_unsigned(1868294587,32),
    to_unsigned(1868396095,32),
    to_unsigned(1868497585,32),
    to_unsigned(1868599058,32),
    to_unsigned(1868700514,32),
    to_unsigned(1868801952,32),
    to_unsigned(1868903374,32),
    to_unsigned(1869004778,32),
    to_unsigned(1869106165,32),
    to_unsigned(1869207535,32),
    to_unsigned(1869308887,32),
    to_unsigned(1869410223,32),
    to_unsigned(1869511541,32),
    to_unsigned(1869612842,32),
    to_unsigned(1869714126,32),
    to_unsigned(1869815393,32),
    to_unsigned(1869916643,32),
    to_unsigned(1870017875,32),
    to_unsigned(1870119090,32),
    to_unsigned(1870220288,32),
    to_unsigned(1870321469,32),
    to_unsigned(1870422633,32),
    to_unsigned(1870523779,32),
    to_unsigned(1870624909,32),
    to_unsigned(1870726021,32),
    to_unsigned(1870827116,32),
    to_unsigned(1870928193,32),
    to_unsigned(1871029254,32),
    to_unsigned(1871130297,32),
    to_unsigned(1871231323,32),
    to_unsigned(1871332332,32),
    to_unsigned(1871433324,32),
    to_unsigned(1871534298,32),
    to_unsigned(1871635255,32),
    to_unsigned(1871736195,32),
    to_unsigned(1871837118,32),
    to_unsigned(1871938024,32),
    to_unsigned(1872038912,32),
    to_unsigned(1872139784,32),
    to_unsigned(1872240638,32),
    to_unsigned(1872341474,32),
    to_unsigned(1872442294,32),
    to_unsigned(1872543096,32),
    to_unsigned(1872643882,32),
    to_unsigned(1872744650,32),
    to_unsigned(1872845400,32),
    to_unsigned(1872946134,32),
    to_unsigned(1873046850,32),
    to_unsigned(1873147549,32),
    to_unsigned(1873248231,32),
    to_unsigned(1873348896,32),
    to_unsigned(1873449543,32),
    to_unsigned(1873550174,32),
    to_unsigned(1873650787,32),
    to_unsigned(1873751383,32),
    to_unsigned(1873851961,32),
    to_unsigned(1873952522,32),
    to_unsigned(1874053067,32),
    to_unsigned(1874153593,32),
    to_unsigned(1874254103,32),
    to_unsigned(1874354596,32),
    to_unsigned(1874455071,32),
    to_unsigned(1874555529,32),
    to_unsigned(1874655970,32),
    to_unsigned(1874756393,32),
    to_unsigned(1874856799,32),
    to_unsigned(1874957188,32),
    to_unsigned(1875057560,32),
    to_unsigned(1875157915,32),
    to_unsigned(1875258252,32),
    to_unsigned(1875358572,32),
    to_unsigned(1875458875,32),
    to_unsigned(1875559161,32),
    to_unsigned(1875659429,32),
    to_unsigned(1875759680,32),
    to_unsigned(1875859914,32),
    to_unsigned(1875960131,32),
    to_unsigned(1876060330,32),
    to_unsigned(1876160513,32),
    to_unsigned(1876260678,32),
    to_unsigned(1876360825,32),
    to_unsigned(1876460956,32),
    to_unsigned(1876561069,32),
    to_unsigned(1876661165,32),
    to_unsigned(1876761244,32),
    to_unsigned(1876861305,32),
    to_unsigned(1876961349,32),
    to_unsigned(1877061376,32),
    to_unsigned(1877161386,32),
    to_unsigned(1877261378,32),
    to_unsigned(1877361353,32),
    to_unsigned(1877461311,32),
    to_unsigned(1877561252,32),
    to_unsigned(1877661175,32),
    to_unsigned(1877761082,32),
    to_unsigned(1877860971,32),
    to_unsigned(1877960842,32),
    to_unsigned(1878060697,32),
    to_unsigned(1878160534,32),
    to_unsigned(1878260353,32),
    to_unsigned(1878360156,32),
    to_unsigned(1878459941,32),
    to_unsigned(1878559709,32),
    to_unsigned(1878659460,32),
    to_unsigned(1878759194,32),
    to_unsigned(1878858910,32),
    to_unsigned(1878958609,32),
    to_unsigned(1879058291,32),
    to_unsigned(1879157955,32),
    to_unsigned(1879257602,32),
    to_unsigned(1879357232,32),
    to_unsigned(1879456845,32),
    to_unsigned(1879556440,32),
    to_unsigned(1879656018,32),
    to_unsigned(1879755579,32),
    to_unsigned(1879855122,32),
    to_unsigned(1879954649,32),
    to_unsigned(1880054158,32),
    to_unsigned(1880153649,32),
    to_unsigned(1880253124,32),
    to_unsigned(1880352581,32),
    to_unsigned(1880452021,32),
    to_unsigned(1880551443,32),
    to_unsigned(1880650848,32),
    to_unsigned(1880750236,32),
    to_unsigned(1880849607,32),
    to_unsigned(1880948960,32),
    to_unsigned(1881048296,32),
    to_unsigned(1881147615,32),
    to_unsigned(1881246917,32),
    to_unsigned(1881346201,32),
    to_unsigned(1881445468,32),
    to_unsigned(1881544717,32),
    to_unsigned(1881643950,32),
    to_unsigned(1881743165,32),
    to_unsigned(1881842363,32),
    to_unsigned(1881941543,32),
    to_unsigned(1882040706,32),
    to_unsigned(1882139852,32),
    to_unsigned(1882238981,32),
    to_unsigned(1882338092,32),
    to_unsigned(1882437186,32),
    to_unsigned(1882536262,32),
    to_unsigned(1882635322,32),
    to_unsigned(1882734364,32),
    to_unsigned(1882833389,32),
    to_unsigned(1882932396,32),
    to_unsigned(1883031386,32),
    to_unsigned(1883130359,32),
    to_unsigned(1883229314,32),
    to_unsigned(1883328253,32),
    to_unsigned(1883427173,32),
    to_unsigned(1883526077,32),
    to_unsigned(1883624963,32),
    to_unsigned(1883723832,32),
    to_unsigned(1883822684,32),
    to_unsigned(1883921518,32),
    to_unsigned(1884020335,32),
    to_unsigned(1884119135,32),
    to_unsigned(1884217917,32),
    to_unsigned(1884316682,32),
    to_unsigned(1884415430,32),
    to_unsigned(1884514160,32),
    to_unsigned(1884612873,32),
    to_unsigned(1884711569,32),
    to_unsigned(1884810247,32),
    to_unsigned(1884908909,32),
    to_unsigned(1885007552,32),
    to_unsigned(1885106179,32),
    to_unsigned(1885204788,32),
    to_unsigned(1885303380,32),
    to_unsigned(1885401954,32),
    to_unsigned(1885500511,32),
    to_unsigned(1885599051,32),
    to_unsigned(1885697574,32),
    to_unsigned(1885796079,32),
    to_unsigned(1885894566,32),
    to_unsigned(1885993037,32),
    to_unsigned(1886091490,32),
    to_unsigned(1886189926,32),
    to_unsigned(1886288344,32),
    to_unsigned(1886386745,32),
    to_unsigned(1886485129,32),
    to_unsigned(1886583496,32),
    to_unsigned(1886681845,32),
    to_unsigned(1886780177,32),
    to_unsigned(1886878491,32),
    to_unsigned(1886976788,32),
    to_unsigned(1887075068,32),
    to_unsigned(1887173330,32),
    to_unsigned(1887271575,32),
    to_unsigned(1887369803,32),
    to_unsigned(1887468013,32),
    to_unsigned(1887566206,32),
    to_unsigned(1887664382,32),
    to_unsigned(1887762540,32),
    to_unsigned(1887860681,32),
    to_unsigned(1887958805,32),
    to_unsigned(1888056911,32),
    to_unsigned(1888155000,32),
    to_unsigned(1888253071,32),
    to_unsigned(1888351125,32),
    to_unsigned(1888449162,32),
    to_unsigned(1888547182,32),
    to_unsigned(1888645184,32),
    to_unsigned(1888743168,32),
    to_unsigned(1888841136,32),
    to_unsigned(1888939086,32),
    to_unsigned(1889037018,32),
    to_unsigned(1889134934,32),
    to_unsigned(1889232832,32),
    to_unsigned(1889330712,32),
    to_unsigned(1889428575,32),
    to_unsigned(1889526421,32),
    to_unsigned(1889624250,32),
    to_unsigned(1889722061,32),
    to_unsigned(1889819854,32),
    to_unsigned(1889917631,32),
    to_unsigned(1890015390,32),
    to_unsigned(1890113131,32),
    to_unsigned(1890210855,32),
    to_unsigned(1890308562,32),
    to_unsigned(1890406252,32),
    to_unsigned(1890503924,32),
    to_unsigned(1890601579,32),
    to_unsigned(1890699216,32),
    to_unsigned(1890796836,32),
    to_unsigned(1890894438,32),
    to_unsigned(1890992024,32),
    to_unsigned(1891089591,32),
    to_unsigned(1891187142,32),
    to_unsigned(1891284675,32),
    to_unsigned(1891382191,32),
    to_unsigned(1891479689,32),
    to_unsigned(1891577170,32),
    to_unsigned(1891674633,32),
    to_unsigned(1891772079,32),
    to_unsigned(1891869508,32),
    to_unsigned(1891966920,32),
    to_unsigned(1892064313,32),
    to_unsigned(1892161690,32),
    to_unsigned(1892259049,32),
    to_unsigned(1892356391,32),
    to_unsigned(1892453715,32),
    to_unsigned(1892551022,32),
    to_unsigned(1892648312,32),
    to_unsigned(1892745584,32),
    to_unsigned(1892842839,32),
    to_unsigned(1892940076,32),
    to_unsigned(1893037296,32),
    to_unsigned(1893134499,32),
    to_unsigned(1893231684,32),
    to_unsigned(1893328852,32),
    to_unsigned(1893426002,32),
    to_unsigned(1893523135,32),
    to_unsigned(1893620251,32),
    to_unsigned(1893717349,32),
    to_unsigned(1893814430,32),
    to_unsigned(1893911493,32),
    to_unsigned(1894008539,32),
    to_unsigned(1894105568,32),
    to_unsigned(1894202579,32),
    to_unsigned(1894299572,32),
    to_unsigned(1894396549,32),
    to_unsigned(1894493508,32),
    to_unsigned(1894590449,32),
    to_unsigned(1894687373,32),
    to_unsigned(1894784280,32),
    to_unsigned(1894881169,32),
    to_unsigned(1894978041,32),
    to_unsigned(1895074895,32),
    to_unsigned(1895171732,32),
    to_unsigned(1895268552,32),
    to_unsigned(1895365354,32),
    to_unsigned(1895462139,32),
    to_unsigned(1895558906,32),
    to_unsigned(1895655656,32),
    to_unsigned(1895752388,32),
    to_unsigned(1895849103,32),
    to_unsigned(1895945801,32),
    to_unsigned(1896042481,32),
    to_unsigned(1896139144,32),
    to_unsigned(1896235789,32),
    to_unsigned(1896332417,32),
    to_unsigned(1896429028,32),
    to_unsigned(1896525621,32),
    to_unsigned(1896622196,32),
    to_unsigned(1896718754,32),
    to_unsigned(1896815295,32),
    to_unsigned(1896911818,32),
    to_unsigned(1897008324,32),
    to_unsigned(1897104813,32),
    to_unsigned(1897201284,32),
    to_unsigned(1897297737,32),
    to_unsigned(1897394173,32),
    to_unsigned(1897490592,32),
    to_unsigned(1897586993,32),
    to_unsigned(1897683377,32),
    to_unsigned(1897779743,32),
    to_unsigned(1897876092,32),
    to_unsigned(1897972423,32),
    to_unsigned(1898068737,32),
    to_unsigned(1898165034,32),
    to_unsigned(1898261313,32),
    to_unsigned(1898357575,32),
    to_unsigned(1898453819,32),
    to_unsigned(1898550046,32),
    to_unsigned(1898646255,32),
    to_unsigned(1898742447,32),
    to_unsigned(1898838621,32),
    to_unsigned(1898934778,32),
    to_unsigned(1899030918,32),
    to_unsigned(1899127040,32),
    to_unsigned(1899223144,32),
    to_unsigned(1899319231,32),
    to_unsigned(1899415301,32),
    to_unsigned(1899511353,32),
    to_unsigned(1899607388,32),
    to_unsigned(1899703405,32),
    to_unsigned(1899799405,32),
    to_unsigned(1899895387,32),
    to_unsigned(1899991352,32),
    to_unsigned(1900087300,32),
    to_unsigned(1900183230,32),
    to_unsigned(1900279142,32),
    to_unsigned(1900375037,32),
    to_unsigned(1900470915,32),
    to_unsigned(1900566775,32),
    to_unsigned(1900662618,32),
    to_unsigned(1900758443,32),
    to_unsigned(1900854250,32),
    to_unsigned(1900950041,32),
    to_unsigned(1901045813,32),
    to_unsigned(1901141569,32),
    to_unsigned(1901237306,32),
    to_unsigned(1901333027,32),
    to_unsigned(1901428730,32),
    to_unsigned(1901524415,32),
    to_unsigned(1901620083,32),
    to_unsigned(1901715733,32),
    to_unsigned(1901811366,32),
    to_unsigned(1901906982,32),
    to_unsigned(1902002580,32),
    to_unsigned(1902098160,32),
    to_unsigned(1902193723,32),
    to_unsigned(1902289268,32),
    to_unsigned(1902384797,32),
    to_unsigned(1902480307,32),
    to_unsigned(1902575800,32),
    to_unsigned(1902671276,32),
    to_unsigned(1902766734,32),
    to_unsigned(1902862174,32),
    to_unsigned(1902957597,32),
    to_unsigned(1903053003,32),
    to_unsigned(1903148391,32),
    to_unsigned(1903243762,32),
    to_unsigned(1903339115,32),
    to_unsigned(1903434450,32),
    to_unsigned(1903529769,32),
    to_unsigned(1903625069,32),
    to_unsigned(1903720352,32),
    to_unsigned(1903815618,32),
    to_unsigned(1903910866,32),
    to_unsigned(1904006097,32),
    to_unsigned(1904101310,32),
    to_unsigned(1904196506,32),
    to_unsigned(1904291684,32),
    to_unsigned(1904386844,32),
    to_unsigned(1904481987,32),
    to_unsigned(1904577113,32),
    to_unsigned(1904672221,32),
    to_unsigned(1904767312,32),
    to_unsigned(1904862385,32),
    to_unsigned(1904957440,32),
    to_unsigned(1905052478,32),
    to_unsigned(1905147499,32),
    to_unsigned(1905242502,32),
    to_unsigned(1905337488,32),
    to_unsigned(1905432456,32),
    to_unsigned(1905527406,32),
    to_unsigned(1905622339,32),
    to_unsigned(1905717255,32),
    to_unsigned(1905812153,32),
    to_unsigned(1905907033,32),
    to_unsigned(1906001896,32),
    to_unsigned(1906096741,32),
    to_unsigned(1906191569,32),
    to_unsigned(1906286380,32),
    to_unsigned(1906381172,32),
    to_unsigned(1906475948,32),
    to_unsigned(1906570706,32),
    to_unsigned(1906665446,32),
    to_unsigned(1906760169,32),
    to_unsigned(1906854874,32),
    to_unsigned(1906949561,32),
    to_unsigned(1907044232,32),
    to_unsigned(1907138884,32),
    to_unsigned(1907233519,32),
    to_unsigned(1907328137,32),
    to_unsigned(1907422737,32),
    to_unsigned(1907517320,32),
    to_unsigned(1907611884,32),
    to_unsigned(1907706432,32),
    to_unsigned(1907800962,32),
    to_unsigned(1907895474,32),
    to_unsigned(1907989969,32),
    to_unsigned(1908084446,32),
    to_unsigned(1908178906,32),
    to_unsigned(1908273348,32),
    to_unsigned(1908367773,32),
    to_unsigned(1908462180,32),
    to_unsigned(1908556570,32),
    to_unsigned(1908650942,32),
    to_unsigned(1908745296,32),
    to_unsigned(1908839633,32),
    to_unsigned(1908933953,32),
    to_unsigned(1909028254,32),
    to_unsigned(1909122539,32),
    to_unsigned(1909216806,32),
    to_unsigned(1909311055,32),
    to_unsigned(1909405286,32),
    to_unsigned(1909499501,32),
    to_unsigned(1909593697,32),
    to_unsigned(1909687876,32),
    to_unsigned(1909782038,32),
    to_unsigned(1909876182,32),
    to_unsigned(1909970308,32),
    to_unsigned(1910064417,32),
    to_unsigned(1910158508,32),
    to_unsigned(1910252582,32),
    to_unsigned(1910346638,32),
    to_unsigned(1910440676,32),
    to_unsigned(1910534697,32),
    to_unsigned(1910628701,32),
    to_unsigned(1910722687,32),
    to_unsigned(1910816655,32),
    to_unsigned(1910910606,32),
    to_unsigned(1911004539,32),
    to_unsigned(1911098455,32),
    to_unsigned(1911192353,32),
    to_unsigned(1911286233,32),
    to_unsigned(1911380096,32),
    to_unsigned(1911473941,32),
    to_unsigned(1911567769,32),
    to_unsigned(1911661579,32),
    to_unsigned(1911755372,32),
    to_unsigned(1911849147,32),
    to_unsigned(1911942905,32),
    to_unsigned(1912036645,32),
    to_unsigned(1912130367,32),
    to_unsigned(1912224072,32),
    to_unsigned(1912317759,32),
    to_unsigned(1912411428,32),
    to_unsigned(1912505081,32),
    to_unsigned(1912598715,32),
    to_unsigned(1912692332,32),
    to_unsigned(1912785931,32),
    to_unsigned(1912879513,32),
    to_unsigned(1912973077,32),
    to_unsigned(1913066624,32),
    to_unsigned(1913160153,32),
    to_unsigned(1913253664,32),
    to_unsigned(1913347158,32),
    to_unsigned(1913440634,32),
    to_unsigned(1913534093,32),
    to_unsigned(1913627534,32),
    to_unsigned(1913720957,32),
    to_unsigned(1913814363,32),
    to_unsigned(1913907751,32),
    to_unsigned(1914001122,32),
    to_unsigned(1914094475,32),
    to_unsigned(1914187810,32),
    to_unsigned(1914281128,32),
    to_unsigned(1914374428,32),
    to_unsigned(1914467711,32),
    to_unsigned(1914560976,32),
    to_unsigned(1914654224,32),
    to_unsigned(1914747454,32),
    to_unsigned(1914840666,32),
    to_unsigned(1914933861,32),
    to_unsigned(1915027038,32),
    to_unsigned(1915120197,32),
    to_unsigned(1915213339,32),
    to_unsigned(1915306463,32),
    to_unsigned(1915399570,32),
    to_unsigned(1915492659,32),
    to_unsigned(1915585731,32),
    to_unsigned(1915678785,32),
    to_unsigned(1915771821,32),
    to_unsigned(1915864839,32),
    to_unsigned(1915957840,32),
    to_unsigned(1916050824,32),
    to_unsigned(1916143790,32),
    to_unsigned(1916236738,32),
    to_unsigned(1916329668,32),
    to_unsigned(1916422581,32),
    to_unsigned(1916515477,32),
    to_unsigned(1916608355,32),
    to_unsigned(1916701215,32),
    to_unsigned(1916794057,32),
    to_unsigned(1916886882,32),
    to_unsigned(1916979689,32),
    to_unsigned(1917072479,32),
    to_unsigned(1917165251,32),
    to_unsigned(1917258005,32),
    to_unsigned(1917350742,32),
    to_unsigned(1917443461,32),
    to_unsigned(1917536163,32),
    to_unsigned(1917628847,32),
    to_unsigned(1917721513,32),
    to_unsigned(1917814162,32),
    to_unsigned(1917906793,32),
    to_unsigned(1917999406,32),
    to_unsigned(1918092002,32),
    to_unsigned(1918184580,32),
    to_unsigned(1918277140,32),
    to_unsigned(1918369683,32),
    to_unsigned(1918462209,32),
    to_unsigned(1918554716,32),
    to_unsigned(1918647206,32),
    to_unsigned(1918739678,32),
    to_unsigned(1918832133,32),
    to_unsigned(1918924570,32),
    to_unsigned(1919016990,32),
    to_unsigned(1919109391,32),
    to_unsigned(1919201775,32),
    to_unsigned(1919294142,32),
    to_unsigned(1919386491,32),
    to_unsigned(1919478822,32),
    to_unsigned(1919571136,32),
    to_unsigned(1919663432,32),
    to_unsigned(1919755710,32),
    to_unsigned(1919847970,32),
    to_unsigned(1919940213,32),
    to_unsigned(1920032439,32),
    to_unsigned(1920124646,32),
    to_unsigned(1920216837,32),
    to_unsigned(1920309009,32),
    to_unsigned(1920401164,32),
    to_unsigned(1920493301,32),
    to_unsigned(1920585420,32),
    to_unsigned(1920677522,32),
    to_unsigned(1920769606,32),
    to_unsigned(1920861673,32),
    to_unsigned(1920953721,32),
    to_unsigned(1921045753,32),
    to_unsigned(1921137766,32),
    to_unsigned(1921229762,32),
    to_unsigned(1921321740,32),
    to_unsigned(1921413701,32),
    to_unsigned(1921505643,32),
    to_unsigned(1921597569,32),
    to_unsigned(1921689476,32),
    to_unsigned(1921781366,32),
    to_unsigned(1921873238,32),
    to_unsigned(1921965093,32),
    to_unsigned(1922056930,32),
    to_unsigned(1922148749,32),
    to_unsigned(1922240550,32),
    to_unsigned(1922332334,32),
    to_unsigned(1922424100,32),
    to_unsigned(1922515849,32),
    to_unsigned(1922607580,32),
    to_unsigned(1922699293,32),
    to_unsigned(1922790989,32),
    to_unsigned(1922882666,32),
    to_unsigned(1922974327,32),
    to_unsigned(1923065969,32),
    to_unsigned(1923157594,32),
    to_unsigned(1923249201,32),
    to_unsigned(1923340790,32),
    to_unsigned(1923432362,32),
    to_unsigned(1923523916,32),
    to_unsigned(1923615453,32),
    to_unsigned(1923706971,32),
    to_unsigned(1923798473,32),
    to_unsigned(1923889956,32),
    to_unsigned(1923981422,32),
    to_unsigned(1924072870,32),
    to_unsigned(1924164300,32),
    to_unsigned(1924255713,32),
    to_unsigned(1924347108,32),
    to_unsigned(1924438485,32),
    to_unsigned(1924529844,32),
    to_unsigned(1924621186,32),
    to_unsigned(1924712510,32),
    to_unsigned(1924803817,32),
    to_unsigned(1924895106,32),
    to_unsigned(1924986377,32),
    to_unsigned(1925077630,32),
    to_unsigned(1925168866,32),
    to_unsigned(1925260084,32),
    to_unsigned(1925351284,32),
    to_unsigned(1925442467,32),
    to_unsigned(1925533632,32),
    to_unsigned(1925624779,32),
    to_unsigned(1925715909,32),
    to_unsigned(1925807020,32),
    to_unsigned(1925898115,32),
    to_unsigned(1925989191,32),
    to_unsigned(1926080250,32),
    to_unsigned(1926171291,32),
    to_unsigned(1926262314,32),
    to_unsigned(1926353320,32),
    to_unsigned(1926444308,32),
    to_unsigned(1926535278,32),
    to_unsigned(1926626230,32),
    to_unsigned(1926717165,32),
    to_unsigned(1926808082,32),
    to_unsigned(1926898981,32),
    to_unsigned(1926989863,32),
    to_unsigned(1927080727,32),
    to_unsigned(1927171573,32),
    to_unsigned(1927262402,32),
    to_unsigned(1927353213,32),
    to_unsigned(1927444006,32),
    to_unsigned(1927534781,32),
    to_unsigned(1927625539,32),
    to_unsigned(1927716279,32),
    to_unsigned(1927807001,32),
    to_unsigned(1927897705,32),
    to_unsigned(1927988392,32),
    to_unsigned(1928079061,32),
    to_unsigned(1928169712,32),
    to_unsigned(1928260346,32),
    to_unsigned(1928350962,32),
    to_unsigned(1928441560,32),
    to_unsigned(1928532140,32),
    to_unsigned(1928622703,32),
    to_unsigned(1928713248,32),
    to_unsigned(1928803775,32),
    to_unsigned(1928894285,32),
    to_unsigned(1928984777,32),
    to_unsigned(1929075251,32),
    to_unsigned(1929165707,32),
    to_unsigned(1929256146,32),
    to_unsigned(1929346566,32),
    to_unsigned(1929436970,32),
    to_unsigned(1929527355,32),
    to_unsigned(1929617723,32),
    to_unsigned(1929708072,32),
    to_unsigned(1929798405,32),
    to_unsigned(1929888719,32),
    to_unsigned(1929979016,32),
    to_unsigned(1930069295,32),
    to_unsigned(1930159556,32),
    to_unsigned(1930249799,32),
    to_unsigned(1930340025,32),
    to_unsigned(1930430233,32),
    to_unsigned(1930520423,32),
    to_unsigned(1930610596,32),
    to_unsigned(1930700751,32),
    to_unsigned(1930790888,32),
    to_unsigned(1930881007,32),
    to_unsigned(1930971108,32),
    to_unsigned(1931061192,32),
    to_unsigned(1931151258,32),
    to_unsigned(1931241306,32),
    to_unsigned(1931331337,32),
    to_unsigned(1931421350,32),
    to_unsigned(1931511345,32),
    to_unsigned(1931601322,32),
    to_unsigned(1931691281,32),
    to_unsigned(1931781223,32),
    to_unsigned(1931871147,32),
    to_unsigned(1931961053,32),
    to_unsigned(1932050942,32),
    to_unsigned(1932140813,32),
    to_unsigned(1932230665,32),
    to_unsigned(1932320501,32),
    to_unsigned(1932410318,32),
    to_unsigned(1932500118,32),
    to_unsigned(1932589900,32),
    to_unsigned(1932679664,32),
    to_unsigned(1932769410,32),
    to_unsigned(1932859139,32),
    to_unsigned(1932948850,32),
    to_unsigned(1933038543,32),
    to_unsigned(1933128218,32),
    to_unsigned(1933217875,32),
    to_unsigned(1933307515,32),
    to_unsigned(1933397137,32),
    to_unsigned(1933486741,32),
    to_unsigned(1933576328,32),
    to_unsigned(1933665897,32),
    to_unsigned(1933755448,32),
    to_unsigned(1933844981,32),
    to_unsigned(1933934496,32),
    to_unsigned(1934023994,32),
    to_unsigned(1934113473,32),
    to_unsigned(1934202935,32),
    to_unsigned(1934292380,32),
    to_unsigned(1934381806,32),
    to_unsigned(1934471215,32),
    to_unsigned(1934560606,32),
    to_unsigned(1934649979,32),
    to_unsigned(1934739334,32),
    to_unsigned(1934828672,32),
    to_unsigned(1934917991,32),
    to_unsigned(1935007293,32),
    to_unsigned(1935096578,32),
    to_unsigned(1935185844,32),
    to_unsigned(1935275093,32),
    to_unsigned(1935364324,32),
    to_unsigned(1935453537,32),
    to_unsigned(1935542732,32),
    to_unsigned(1935631909,32),
    to_unsigned(1935721069,32),
    to_unsigned(1935810211,32),
    to_unsigned(1935899335,32),
    to_unsigned(1935988441,32),
    to_unsigned(1936077530,32),
    to_unsigned(1936166600,32),
    to_unsigned(1936255653,32),
    to_unsigned(1936344688,32),
    to_unsigned(1936433706,32),
    to_unsigned(1936522705,32),
    to_unsigned(1936611687,32),
    to_unsigned(1936700651,32),
    to_unsigned(1936789597,32),
    to_unsigned(1936878525,32),
    to_unsigned(1936967436,32),
    to_unsigned(1937056328,32),
    to_unsigned(1937145203,32),
    to_unsigned(1937234060,32),
    to_unsigned(1937322900,32),
    to_unsigned(1937411721,32),
    to_unsigned(1937500525,32),
    to_unsigned(1937589311,32),
    to_unsigned(1937678079,32),
    to_unsigned(1937766829,32),
    to_unsigned(1937855561,32),
    to_unsigned(1937944276,32),
    to_unsigned(1938032973,32),
    to_unsigned(1938121652,32),
    to_unsigned(1938210313,32),
    to_unsigned(1938298956,32),
    to_unsigned(1938387582,32),
    to_unsigned(1938476189,32),
    to_unsigned(1938564779,32),
    to_unsigned(1938653351,32),
    to_unsigned(1938741906,32),
    to_unsigned(1938830442,32),
    to_unsigned(1938918961,32),
    to_unsigned(1939007462,32),
    to_unsigned(1939095945,32),
    to_unsigned(1939184410,32),
    to_unsigned(1939272857,32),
    to_unsigned(1939361287,32),
    to_unsigned(1939449698,32),
    to_unsigned(1939538092,32),
    to_unsigned(1939626468,32),
    to_unsigned(1939714826,32),
    to_unsigned(1939803167,32),
    to_unsigned(1939891489,32),
    to_unsigned(1939979794,32),
    to_unsigned(1940068081,32),
    to_unsigned(1940156350,32),
    to_unsigned(1940244601,32),
    to_unsigned(1940332834,32),
    to_unsigned(1940421050,32),
    to_unsigned(1940509248,32),
    to_unsigned(1940597427,32),
    to_unsigned(1940685589,32),
    to_unsigned(1940773734,32),
    to_unsigned(1940861860,32),
    to_unsigned(1940949968,32),
    to_unsigned(1941038059,32),
    to_unsigned(1941126132,32),
    to_unsigned(1941214187,32),
    to_unsigned(1941302224,32),
    to_unsigned(1941390243,32),
    to_unsigned(1941478245,32),
    to_unsigned(1941566228,32),
    to_unsigned(1941654194,32),
    to_unsigned(1941742142,32),
    to_unsigned(1941830072,32),
    to_unsigned(1941917984,32),
    to_unsigned(1942005879,32),
    to_unsigned(1942093755,32),
    to_unsigned(1942181614,32),
    to_unsigned(1942269455,32),
    to_unsigned(1942357278,32),
    to_unsigned(1942445083,32),
    to_unsigned(1942532870,32),
    to_unsigned(1942620639,32),
    to_unsigned(1942708391,32),
    to_unsigned(1942796125,32),
    to_unsigned(1942883840,32),
    to_unsigned(1942971538,32),
    to_unsigned(1943059218,32),
    to_unsigned(1943146881,32),
    to_unsigned(1943234525,32),
    to_unsigned(1943322152,32),
    to_unsigned(1943409760,32),
    to_unsigned(1943497351,32),
    to_unsigned(1943584924,32),
    to_unsigned(1943672479,32),
    to_unsigned(1943760016,32),
    to_unsigned(1943847536,32),
    to_unsigned(1943935037,32),
    to_unsigned(1944022521,32),
    to_unsigned(1944109986,32),
    to_unsigned(1944197434,32),
    to_unsigned(1944284864,32),
    to_unsigned(1944372276,32),
    to_unsigned(1944459671,32),
    to_unsigned(1944547047,32),
    to_unsigned(1944634405,32),
    to_unsigned(1944721746,32),
    to_unsigned(1944809069,32),
    to_unsigned(1944896374,32),
    to_unsigned(1944983661,32),
    to_unsigned(1945070930,32),
    to_unsigned(1945158181,32),
    to_unsigned(1945245414,32),
    to_unsigned(1945332630,32),
    to_unsigned(1945419827,32),
    to_unsigned(1945507007,32),
    to_unsigned(1945594169,32),
    to_unsigned(1945681313,32),
    to_unsigned(1945768439,32),
    to_unsigned(1945855547,32),
    to_unsigned(1945942637,32),
    to_unsigned(1946029710,32),
    to_unsigned(1946116764,32),
    to_unsigned(1946203801,32),
    to_unsigned(1946290820,32),
    to_unsigned(1946377821,32),
    to_unsigned(1946464803,32),
    to_unsigned(1946551769,32),
    to_unsigned(1946638716,32),
    to_unsigned(1946725645,32),
    to_unsigned(1946812556,32),
    to_unsigned(1946899450,32),
    to_unsigned(1946986325,32),
    to_unsigned(1947073183,32),
    to_unsigned(1947160023,32),
    to_unsigned(1947246845,32),
    to_unsigned(1947333649,32),
    to_unsigned(1947420435,32),
    to_unsigned(1947507203,32),
    to_unsigned(1947593954,32),
    to_unsigned(1947680686,32),
    to_unsigned(1947767400,32),
    to_unsigned(1947854097,32),
    to_unsigned(1947940776,32),
    to_unsigned(1948027437,32),
    to_unsigned(1948114079,32),
    to_unsigned(1948200704,32),
    to_unsigned(1948287311,32),
    to_unsigned(1948373901,32),
    to_unsigned(1948460472,32),
    to_unsigned(1948547025,32),
    to_unsigned(1948633561,32),
    to_unsigned(1948720078,32),
    to_unsigned(1948806578,32),
    to_unsigned(1948893059,32),
    to_unsigned(1948979523,32),
    to_unsigned(1949065969,32),
    to_unsigned(1949152397,32),
    to_unsigned(1949238807,32),
    to_unsigned(1949325199,32),
    to_unsigned(1949411573,32),
    to_unsigned(1949497930,32),
    to_unsigned(1949584268,32),
    to_unsigned(1949670588,32),
    to_unsigned(1949756891,32),
    to_unsigned(1949843176,32),
    to_unsigned(1949929442,32),
    to_unsigned(1950015691,32),
    to_unsigned(1950101922,32),
    to_unsigned(1950188135,32),
    to_unsigned(1950274330,32),
    to_unsigned(1950360507,32),
    to_unsigned(1950446666,32),
    to_unsigned(1950532807,32),
    to_unsigned(1950618930,32),
    to_unsigned(1950705036,32),
    to_unsigned(1950791123,32),
    to_unsigned(1950877193,32),
    to_unsigned(1950963244,32),
    to_unsigned(1951049278,32),
    to_unsigned(1951135293,32),
    to_unsigned(1951221291,32),
    to_unsigned(1951307271,32),
    to_unsigned(1951393233,32),
    to_unsigned(1951479177,32),
    to_unsigned(1951565103,32),
    to_unsigned(1951651011,32),
    to_unsigned(1951736901,32),
    to_unsigned(1951822773,32),
    to_unsigned(1951908627,32),
    to_unsigned(1951994464,32),
    to_unsigned(1952080282,32),
    to_unsigned(1952166082,32),
    to_unsigned(1952251865,32),
    to_unsigned(1952337629,32),
    to_unsigned(1952423376,32),
    to_unsigned(1952509105,32),
    to_unsigned(1952594815,32),
    to_unsigned(1952680508,32),
    to_unsigned(1952766183,32),
    to_unsigned(1952851840,32),
    to_unsigned(1952937479,32),
    to_unsigned(1953023100,32),
    to_unsigned(1953108703,32),
    to_unsigned(1953194288,32),
    to_unsigned(1953279855,32),
    to_unsigned(1953365404,32),
    to_unsigned(1953450935,32),
    to_unsigned(1953536448,32),
    to_unsigned(1953621943,32),
    to_unsigned(1953707421,32),
    to_unsigned(1953792880,32),
    to_unsigned(1953878321,32),
    to_unsigned(1953963745,32),
    to_unsigned(1954049150,32),
    to_unsigned(1954134538,32),
    to_unsigned(1954219907,32),
    to_unsigned(1954305259,32),
    to_unsigned(1954390593,32),
    to_unsigned(1954475908,32),
    to_unsigned(1954561206,32),
    to_unsigned(1954646486,32),
    to_unsigned(1954731747,32),
    to_unsigned(1954816991,32),
    to_unsigned(1954902217,32),
    to_unsigned(1954987425,32),
    to_unsigned(1955072615,32),
    to_unsigned(1955157787,32),
    to_unsigned(1955242941,32),
    to_unsigned(1955328077,32),
    to_unsigned(1955413195,32),
    to_unsigned(1955498295,32),
    to_unsigned(1955583377,32),
    to_unsigned(1955668441,32),
    to_unsigned(1955753487,32),
    to_unsigned(1955838515,32),
    to_unsigned(1955923525,32),
    to_unsigned(1956008517,32),
    to_unsigned(1956093491,32),
    to_unsigned(1956178448,32),
    to_unsigned(1956263386,32),
    to_unsigned(1956348306,32),
    to_unsigned(1956433208,32),
    to_unsigned(1956518093,32),
    to_unsigned(1956602959,32),
    to_unsigned(1956687807,32),
    to_unsigned(1956772637,32),
    to_unsigned(1956857450,32),
    to_unsigned(1956942244,32),
    to_unsigned(1957027021,32),
    to_unsigned(1957111779,32),
    to_unsigned(1957196519,32),
    to_unsigned(1957281242,32),
    to_unsigned(1957365946,32),
    to_unsigned(1957450632,32),
    to_unsigned(1957535301,32),
    to_unsigned(1957619951,32),
    to_unsigned(1957704584,32),
    to_unsigned(1957789198,32),
    to_unsigned(1957873795,32),
    to_unsigned(1957958373,32),
    to_unsigned(1958042933,32),
    to_unsigned(1958127476,32),
    to_unsigned(1958212000,32),
    to_unsigned(1958296507,32),
    to_unsigned(1958380995,32),
    to_unsigned(1958465466,32),
    to_unsigned(1958549918,32),
    to_unsigned(1958634353,32),
    to_unsigned(1958718769,32),
    to_unsigned(1958803167,32),
    to_unsigned(1958887548,32),
    to_unsigned(1958971910,32),
    to_unsigned(1959056255,32),
    to_unsigned(1959140581,32),
    to_unsigned(1959224890,32),
    to_unsigned(1959309180,32),
    to_unsigned(1959393452,32),
    to_unsigned(1959477707,32),
    to_unsigned(1959561943,32),
    to_unsigned(1959646161,32),
    to_unsigned(1959730362,32),
    to_unsigned(1959814544,32),
    to_unsigned(1959898708,32),
    to_unsigned(1959982855,32),
    to_unsigned(1960066983,32),
    to_unsigned(1960151093,32),
    to_unsigned(1960235185,32),
    to_unsigned(1960319260,32),
    to_unsigned(1960403316,32),
    to_unsigned(1960487354,32),
    to_unsigned(1960571374,32),
    to_unsigned(1960655376,32),
    to_unsigned(1960739361,32),
    to_unsigned(1960823327,32),
    to_unsigned(1960907275,32),
    to_unsigned(1960991205,32),
    to_unsigned(1961075117,32),
    to_unsigned(1961159011,32),
    to_unsigned(1961242887,32),
    to_unsigned(1961326745,32),
    to_unsigned(1961410585,32),
    to_unsigned(1961494407,32),
    to_unsigned(1961578210,32),
    to_unsigned(1961661996,32),
    to_unsigned(1961745764,32),
    to_unsigned(1961829514,32),
    to_unsigned(1961913246,32),
    to_unsigned(1961996959,32),
    to_unsigned(1962080655,32),
    to_unsigned(1962164333,32),
    to_unsigned(1962247992,32),
    to_unsigned(1962331634,32),
    to_unsigned(1962415257,32),
    to_unsigned(1962498863,32),
    to_unsigned(1962582450,32),
    to_unsigned(1962666020,32),
    to_unsigned(1962749571,32),
    to_unsigned(1962833104,32),
    to_unsigned(1962916620,32),
    to_unsigned(1963000117,32),
    to_unsigned(1963083596,32),
    to_unsigned(1963167057,32),
    to_unsigned(1963250500,32),
    to_unsigned(1963333925,32),
    to_unsigned(1963417332,32),
    to_unsigned(1963500721,32),
    to_unsigned(1963584092,32),
    to_unsigned(1963667445,32),
    to_unsigned(1963750780,32),
    to_unsigned(1963834097,32),
    to_unsigned(1963917395,32),
    to_unsigned(1964000676,32),
    to_unsigned(1964083939,32),
    to_unsigned(1964167183,32),
    to_unsigned(1964250410,32),
    to_unsigned(1964333618,32),
    to_unsigned(1964416809,32),
    to_unsigned(1964499981,32),
    to_unsigned(1964583135,32),
    to_unsigned(1964666272,32),
    to_unsigned(1964749390,32),
    to_unsigned(1964832490,32),
    to_unsigned(1964915572,32),
    to_unsigned(1964998636,32),
    to_unsigned(1965081682,32),
    to_unsigned(1965164710,32),
    to_unsigned(1965247719,32),
    to_unsigned(1965330711,32),
    to_unsigned(1965413685,32),
    to_unsigned(1965496640,32),
    to_unsigned(1965579578,32),
    to_unsigned(1965662497,32),
    to_unsigned(1965745399,32),
    to_unsigned(1965828282,32),
    to_unsigned(1965911147,32),
    to_unsigned(1965993995,32),
    to_unsigned(1966076824,32),
    to_unsigned(1966159635,32),
    to_unsigned(1966242428,32),
    to_unsigned(1966325203,32),
    to_unsigned(1966407960,32),
    to_unsigned(1966490698,32),
    to_unsigned(1966573419,32),
    to_unsigned(1966656122,32),
    to_unsigned(1966738806,32),
    to_unsigned(1966821473,32),
    to_unsigned(1966904121,32),
    to_unsigned(1966986751,32),
    to_unsigned(1967069363,32),
    to_unsigned(1967151958,32),
    to_unsigned(1967234534,32),
    to_unsigned(1967317092,32),
    to_unsigned(1967399631,32),
    to_unsigned(1967482153,32),
    to_unsigned(1967564657,32),
    to_unsigned(1967647143,32),
    to_unsigned(1967729610,32),
    to_unsigned(1967812060,32),
    to_unsigned(1967894491,32),
    to_unsigned(1967976904,32),
    to_unsigned(1968059299,32),
    to_unsigned(1968141677,32),
    to_unsigned(1968224036,32),
    to_unsigned(1968306377,32),
    to_unsigned(1968388699,32),
    to_unsigned(1968471004,32),
    to_unsigned(1968553291,32),
    to_unsigned(1968635559,32),
    to_unsigned(1968717810,32),
    to_unsigned(1968800042,32),
    to_unsigned(1968882256,32),
    to_unsigned(1968964453,32),
    to_unsigned(1969046631,32),
    to_unsigned(1969128791,32),
    to_unsigned(1969210932,32),
    to_unsigned(1969293056,32),
    to_unsigned(1969375162,32),
    to_unsigned(1969457249,32),
    to_unsigned(1969539319,32),
    to_unsigned(1969621370,32),
    to_unsigned(1969703403,32),
    to_unsigned(1969785419,32),
    to_unsigned(1969867416,32),
    to_unsigned(1969949395,32),
    to_unsigned(1970031355,32),
    to_unsigned(1970113298,32),
    to_unsigned(1970195223,32),
    to_unsigned(1970277129,32),
    to_unsigned(1970359018,32),
    to_unsigned(1970440888,32),
    to_unsigned(1970522740,32),
    to_unsigned(1970604574,32),
    to_unsigned(1970686390,32),
    to_unsigned(1970768188,32),
    to_unsigned(1970849968,32),
    to_unsigned(1970931729,32),
    to_unsigned(1971013473,32),
    to_unsigned(1971095198,32),
    to_unsigned(1971176905,32),
    to_unsigned(1971258594,32),
    to_unsigned(1971340265,32),
    to_unsigned(1971421918,32),
    to_unsigned(1971503553,32),
    to_unsigned(1971585170,32),
    to_unsigned(1971666768,32),
    to_unsigned(1971748349,32),
    to_unsigned(1971829911,32),
    to_unsigned(1971911455,32),
    to_unsigned(1971992981,32),
    to_unsigned(1972074489,32),
    to_unsigned(1972155979,32),
    to_unsigned(1972237450,32),
    to_unsigned(1972318904,32),
    to_unsigned(1972400339,32),
    to_unsigned(1972481756,32),
    to_unsigned(1972563156,32),
    to_unsigned(1972644537,32),
    to_unsigned(1972725899,32),
    to_unsigned(1972807244,32),
    to_unsigned(1972888571,32),
    to_unsigned(1972969879,32),
    to_unsigned(1973051170,32),
    to_unsigned(1973132442,32),
    to_unsigned(1973213696,32),
    to_unsigned(1973294932,32),
    to_unsigned(1973376149,32),
    to_unsigned(1973457349,32),
    to_unsigned(1973538531,32),
    to_unsigned(1973619694,32),
    to_unsigned(1973700839,32),
    to_unsigned(1973781966,32),
    to_unsigned(1973863075,32),
    to_unsigned(1973944166,32),
    to_unsigned(1974025239,32),
    to_unsigned(1974106293,32),
    to_unsigned(1974187329,32),
    to_unsigned(1974268348,32),
    to_unsigned(1974349348,32),
    to_unsigned(1974430330,32),
    to_unsigned(1974511293,32),
    to_unsigned(1974592239,32),
    to_unsigned(1974673166,32),
    to_unsigned(1974754076,32),
    to_unsigned(1974834967,32),
    to_unsigned(1974915840,32),
    to_unsigned(1974996695,32),
    to_unsigned(1975077532,32),
    to_unsigned(1975158350,32),
    to_unsigned(1975239150,32),
    to_unsigned(1975319933,32),
    to_unsigned(1975400697,32),
    to_unsigned(1975481443,32),
    to_unsigned(1975562170,32),
    to_unsigned(1975642880,32),
    to_unsigned(1975723572,32),
    to_unsigned(1975804245,32),
    to_unsigned(1975884900,32),
    to_unsigned(1975965537,32),
    to_unsigned(1976046156,32),
    to_unsigned(1976126756,32),
    to_unsigned(1976207339,32),
    to_unsigned(1976287903,32),
    to_unsigned(1976368449,32),
    to_unsigned(1976448977,32),
    to_unsigned(1976529487,32),
    to_unsigned(1976609979,32),
    to_unsigned(1976690452,32),
    to_unsigned(1976770907,32),
    to_unsigned(1976851345,32),
    to_unsigned(1976931764,32),
    to_unsigned(1977012164,32),
    to_unsigned(1977092547,32),
    to_unsigned(1977172911,32),
    to_unsigned(1977253258,32),
    to_unsigned(1977333586,32),
    to_unsigned(1977413896,32),
    to_unsigned(1977494187,32),
    to_unsigned(1977574461,32),
    to_unsigned(1977654716,32),
    to_unsigned(1977734954,32),
    to_unsigned(1977815173,32),
    to_unsigned(1977895374,32),
    to_unsigned(1977975556,32),
    to_unsigned(1978055721,32),
    to_unsigned(1978135867,32),
    to_unsigned(1978215995,32),
    to_unsigned(1978296105,32),
    to_unsigned(1978376197,32),
    to_unsigned(1978456270,32),
    to_unsigned(1978536326,32),
    to_unsigned(1978616363,32),
    to_unsigned(1978696382,32),
    to_unsigned(1978776383,32),
    to_unsigned(1978856366,32),
    to_unsigned(1978936330,32),
    to_unsigned(1979016276,32),
    to_unsigned(1979096204,32),
    to_unsigned(1979176114,32),
    to_unsigned(1979256006,32),
    to_unsigned(1979335879,32),
    to_unsigned(1979415735,32),
    to_unsigned(1979495572,32),
    to_unsigned(1979575391,32),
    to_unsigned(1979655191,32),
    to_unsigned(1979734974,32),
    to_unsigned(1979814738,32),
    to_unsigned(1979894484,32),
    to_unsigned(1979974212,32),
    to_unsigned(1980053922,32),
    to_unsigned(1980133614,32),
    to_unsigned(1980213287,32),
    to_unsigned(1980292942,32),
    to_unsigned(1980372579,32),
    to_unsigned(1980452198,32),
    to_unsigned(1980531798,32),
    to_unsigned(1980611380,32),
    to_unsigned(1980690945,32),
    to_unsigned(1980770490,32),
    to_unsigned(1980850018,32),
    to_unsigned(1980929528,32),
    to_unsigned(1981009019,32),
    to_unsigned(1981088492,32),
    to_unsigned(1981167947,32),
    to_unsigned(1981247383,32),
    to_unsigned(1981326802,32),
    to_unsigned(1981406202,32),
    to_unsigned(1981485584,32),
    to_unsigned(1981564948,32),
    to_unsigned(1981644294,32),
    to_unsigned(1981723621,32),
    to_unsigned(1981802930,32),
    to_unsigned(1981882221,32),
    to_unsigned(1981961494,32),
    to_unsigned(1982040748,32),
    to_unsigned(1982119985,32),
    to_unsigned(1982199203,32),
    to_unsigned(1982278402,32),
    to_unsigned(1982357584,32),
    to_unsigned(1982436747,32),
    to_unsigned(1982515893,32),
    to_unsigned(1982595020,32),
    to_unsigned(1982674128,32),
    to_unsigned(1982753219,32),
    to_unsigned(1982832291,32),
    to_unsigned(1982911345,32),
    to_unsigned(1982990381,32),
    to_unsigned(1983069399,32),
    to_unsigned(1983148398,32),
    to_unsigned(1983227379,32),
    to_unsigned(1983306342,32),
    to_unsigned(1983385287,32),
    to_unsigned(1983464213,32),
    to_unsigned(1983543121,32),
    to_unsigned(1983622011,32),
    to_unsigned(1983700883,32),
    to_unsigned(1983779737,32),
    to_unsigned(1983858572,32),
    to_unsigned(1983937389,32),
    to_unsigned(1984016188,32),
    to_unsigned(1984094968,32),
    to_unsigned(1984173731,32),
    to_unsigned(1984252475,32),
    to_unsigned(1984331201,32),
    to_unsigned(1984409908,32),
    to_unsigned(1984488598,32),
    to_unsigned(1984567269,32),
    to_unsigned(1984645922,32),
    to_unsigned(1984724557,32),
    to_unsigned(1984803173,32),
    to_unsigned(1984881771,32),
    to_unsigned(1984960351,32),
    to_unsigned(1985038913,32),
    to_unsigned(1985117456,32),
    to_unsigned(1985195981,32),
    to_unsigned(1985274488,32),
    to_unsigned(1985352977,32),
    to_unsigned(1985431447,32),
    to_unsigned(1985509900,32),
    to_unsigned(1985588334,32),
    to_unsigned(1985666749,32),
    to_unsigned(1985745147,32),
    to_unsigned(1985823526,32),
    to_unsigned(1985901887,32),
    to_unsigned(1985980230,32),
    to_unsigned(1986058554,32),
    to_unsigned(1986136860,32),
    to_unsigned(1986215148,32),
    to_unsigned(1986293418,32),
    to_unsigned(1986371669,32),
    to_unsigned(1986449902,32),
    to_unsigned(1986528117,32),
    to_unsigned(1986606314,32),
    to_unsigned(1986684492,32),
    to_unsigned(1986762652,32),
    to_unsigned(1986840794,32),
    to_unsigned(1986918918,32),
    to_unsigned(1986997023,32),
    to_unsigned(1987075110,32),
    to_unsigned(1987153179,32),
    to_unsigned(1987231229,32),
    to_unsigned(1987309262,32),
    to_unsigned(1987387276,32),
    to_unsigned(1987465271,32),
    to_unsigned(1987543249,32),
    to_unsigned(1987621208,32),
    to_unsigned(1987699149,32),
    to_unsigned(1987777072,32),
    to_unsigned(1987854976,32),
    to_unsigned(1987932862,32),
    to_unsigned(1988010730,32),
    to_unsigned(1988088580,32),
    to_unsigned(1988166411,32),
    to_unsigned(1988244224,32),
    to_unsigned(1988322019,32),
    to_unsigned(1988399795,32),
    to_unsigned(1988477553,32),
    to_unsigned(1988555293,32),
    to_unsigned(1988633015,32),
    to_unsigned(1988710718,32),
    to_unsigned(1988788403,32),
    to_unsigned(1988866070,32),
    to_unsigned(1988943718,32),
    to_unsigned(1989021349,32),
    to_unsigned(1989098961,32),
    to_unsigned(1989176554,32),
    to_unsigned(1989254130,32),
    to_unsigned(1989331687,32),
    to_unsigned(1989409226,32),
    to_unsigned(1989486746,32),
    to_unsigned(1989564248,32),
    to_unsigned(1989641732,32),
    to_unsigned(1989719198,32),
    to_unsigned(1989796645,32),
    to_unsigned(1989874074,32),
    to_unsigned(1989951485,32),
    to_unsigned(1990028878,32),
    to_unsigned(1990106252,32),
    to_unsigned(1990183608,32),
    to_unsigned(1990260945,32),
    to_unsigned(1990338265,32),
    to_unsigned(1990415566,32),
    to_unsigned(1990492848,32),
    to_unsigned(1990570113,32),
    to_unsigned(1990647359,32),
    to_unsigned(1990724587,32),
    to_unsigned(1990801796,32),
    to_unsigned(1990878988,32),
    to_unsigned(1990956161,32),
    to_unsigned(1991033315,32),
    to_unsigned(1991110452,32),
    to_unsigned(1991187570,32),
    to_unsigned(1991264669,32),
    to_unsigned(1991341751,32),
    to_unsigned(1991418814,32),
    to_unsigned(1991495859,32),
    to_unsigned(1991572885,32),
    to_unsigned(1991649893,32),
    to_unsigned(1991726883,32),
    to_unsigned(1991803855,32),
    to_unsigned(1991880808,32),
    to_unsigned(1991957743,32),
    to_unsigned(1992034660,32),
    to_unsigned(1992111558,32),
    to_unsigned(1992188438,32),
    to_unsigned(1992265300,32),
    to_unsigned(1992342143,32),
    to_unsigned(1992418969,32),
    to_unsigned(1992495775,32),
    to_unsigned(1992572564,32),
    to_unsigned(1992649334,32),
    to_unsigned(1992726086,32),
    to_unsigned(1992802819,32),
    to_unsigned(1992879535,32),
    to_unsigned(1992956232,32),
    to_unsigned(1993032910,32),
    to_unsigned(1993109570,32),
    to_unsigned(1993186212,32),
    to_unsigned(1993262836,32),
    to_unsigned(1993339441,32),
    to_unsigned(1993416028,32),
    to_unsigned(1993492597,32),
    to_unsigned(1993569147,32),
    to_unsigned(1993645679,32),
    to_unsigned(1993722193,32),
    to_unsigned(1993798688,32),
    to_unsigned(1993875165,32),
    to_unsigned(1993951624,32),
    to_unsigned(1994028064,32),
    to_unsigned(1994104486,32),
    to_unsigned(1994180890,32),
    to_unsigned(1994257275,32),
    to_unsigned(1994333643,32),
    to_unsigned(1994409991,32),
    to_unsigned(1994486322,32),
    to_unsigned(1994562634,32),
    to_unsigned(1994638927,32),
    to_unsigned(1994715203,32),
    to_unsigned(1994791460,32),
    to_unsigned(1994867699,32),
    to_unsigned(1994943919,32),
    to_unsigned(1995020121,32),
    to_unsigned(1995096305,32),
    to_unsigned(1995172470,32),
    to_unsigned(1995248617,32),
    to_unsigned(1995324746,32),
    to_unsigned(1995400856,32),
    to_unsigned(1995476948,32),
    to_unsigned(1995553022,32),
    to_unsigned(1995629077,32),
    to_unsigned(1995705114,32),
    to_unsigned(1995781133,32),
    to_unsigned(1995857133,32),
    to_unsigned(1995933115,32),
    to_unsigned(1996009079,32),
    to_unsigned(1996085024,32),
    to_unsigned(1996160951,32),
    to_unsigned(1996236859,32),
    to_unsigned(1996312750,32),
    to_unsigned(1996388621,32),
    to_unsigned(1996464475,32),
    to_unsigned(1996540310,32),
    to_unsigned(1996616127,32),
    to_unsigned(1996691925,32),
    to_unsigned(1996767705,32),
    to_unsigned(1996843467,32),
    to_unsigned(1996919211,32),
    to_unsigned(1996994936,32),
    to_unsigned(1997070642,32),
    to_unsigned(1997146331,32),
    to_unsigned(1997222001,32),
    to_unsigned(1997297652,32),
    to_unsigned(1997373285,32),
    to_unsigned(1997448900,32),
    to_unsigned(1997524497,32),
    to_unsigned(1997600075,32),
    to_unsigned(1997675635,32),
    to_unsigned(1997751176,32),
    to_unsigned(1997826699,32),
    to_unsigned(1997902204,32),
    to_unsigned(1997977690,32),
    to_unsigned(1998053158,32),
    to_unsigned(1998128608,32),
    to_unsigned(1998204039,32),
    to_unsigned(1998279452,32),
    to_unsigned(1998354847,32),
    to_unsigned(1998430223,32),
    to_unsigned(1998505581,32),
    to_unsigned(1998580920,32),
    to_unsigned(1998656241,32),
    to_unsigned(1998731544,32),
    to_unsigned(1998806828,32),
    to_unsigned(1998882094,32),
    to_unsigned(1998957342,32),
    to_unsigned(1999032571,32),
    to_unsigned(1999107782,32),
    to_unsigned(1999182974,32),
    to_unsigned(1999258148,32),
    to_unsigned(1999333304,32),
    to_unsigned(1999408441,32),
    to_unsigned(1999483560,32),
    to_unsigned(1999558660,32),
    to_unsigned(1999633743,32),
    to_unsigned(1999708806,32),
    to_unsigned(1999783852,32),
    to_unsigned(1999858879,32),
    to_unsigned(1999933888,32),
    to_unsigned(2000008878,32),
    to_unsigned(2000083850,32),
    to_unsigned(2000158803,32),
    to_unsigned(2000233738,32),
    to_unsigned(2000308655,32),
    to_unsigned(2000383553,32),
    to_unsigned(2000458433,32),
    to_unsigned(2000533295,32),
    to_unsigned(2000608138,32),
    to_unsigned(2000682963,32),
    to_unsigned(2000757769,32),
    to_unsigned(2000832557,32),
    to_unsigned(2000907327,32),
    to_unsigned(2000982078,32),
    to_unsigned(2001056811,32),
    to_unsigned(2001131525,32),
    to_unsigned(2001206221,32),
    to_unsigned(2001280899,32),
    to_unsigned(2001355558,32),
    to_unsigned(2001430199,32),
    to_unsigned(2001504821,32),
    to_unsigned(2001579425,32),
    to_unsigned(2001654011,32),
    to_unsigned(2001728578,32),
    to_unsigned(2001803127,32),
    to_unsigned(2001877658,32),
    to_unsigned(2001952170,32),
    to_unsigned(2002026663,32),
    to_unsigned(2002101139,32),
    to_unsigned(2002175596,32),
    to_unsigned(2002250034,32),
    to_unsigned(2002324454,32),
    to_unsigned(2002398856,32),
    to_unsigned(2002473239,32),
    to_unsigned(2002547604,32),
    to_unsigned(2002621950,32),
    to_unsigned(2002696278,32),
    to_unsigned(2002770588,32),
    to_unsigned(2002844879,32),
    to_unsigned(2002919152,32),
    to_unsigned(2002993406,32),
    to_unsigned(2003067642,32),
    to_unsigned(2003141860,32),
    to_unsigned(2003216059,32),
    to_unsigned(2003290240,32),
    to_unsigned(2003364402,32),
    to_unsigned(2003438546,32),
    to_unsigned(2003512671,32),
    to_unsigned(2003586778,32),
    to_unsigned(2003660867,32),
    to_unsigned(2003734937,32),
    to_unsigned(2003808989,32),
    to_unsigned(2003883022,32),
    to_unsigned(2003957037,32),
    to_unsigned(2004031034,32),
    to_unsigned(2004105012,32),
    to_unsigned(2004178972,32),
    to_unsigned(2004252913,32),
    to_unsigned(2004326836,32),
    to_unsigned(2004400740,32),
    to_unsigned(2004474626,32),
    to_unsigned(2004548494,32),
    to_unsigned(2004622343,32),
    to_unsigned(2004696174,32),
    to_unsigned(2004769986,32),
    to_unsigned(2004843780,32),
    to_unsigned(2004917556,32),
    to_unsigned(2004991313,32),
    to_unsigned(2005065051,32),
    to_unsigned(2005138771,32),
    to_unsigned(2005212473,32),
    to_unsigned(2005286156,32),
    to_unsigned(2005359821,32),
    to_unsigned(2005433468,32),
    to_unsigned(2005507096,32),
    to_unsigned(2005580705,32),
    to_unsigned(2005654297,32),
    to_unsigned(2005727869,32),
    to_unsigned(2005801424,32),
    to_unsigned(2005874959,32),
    to_unsigned(2005948477,32),
    to_unsigned(2006021976,32),
    to_unsigned(2006095456,32),
    to_unsigned(2006168918,32),
    to_unsigned(2006242362,32),
    to_unsigned(2006315787,32),
    to_unsigned(2006389194,32),
    to_unsigned(2006462582,32),
    to_unsigned(2006535952,32),
    to_unsigned(2006609304,32),
    to_unsigned(2006682637,32),
    to_unsigned(2006755951,32),
    to_unsigned(2006829247,32),
    to_unsigned(2006902525,32),
    to_unsigned(2006975784,32),
    to_unsigned(2007049025,32),
    to_unsigned(2007122247,32),
    to_unsigned(2007195451,32),
    to_unsigned(2007268636,32),
    to_unsigned(2007341803,32),
    to_unsigned(2007414952,32),
    to_unsigned(2007488082,32),
    to_unsigned(2007561194,32),
    to_unsigned(2007634287,32),
    to_unsigned(2007707361,32),
    to_unsigned(2007780418,32),
    to_unsigned(2007853455,32),
    to_unsigned(2007926475,32),
    to_unsigned(2007999476,32),
    to_unsigned(2008072458,32),
    to_unsigned(2008145422,32),
    to_unsigned(2008218367,32),
    to_unsigned(2008291295,32),
    to_unsigned(2008364203,32),
    to_unsigned(2008437093,32),
    to_unsigned(2008509965,32),
    to_unsigned(2008582818,32),
    to_unsigned(2008655653,32),
    to_unsigned(2008728469,32),
    to_unsigned(2008801267,32),
    to_unsigned(2008874046,32),
    to_unsigned(2008946807,32),
    to_unsigned(2009019550,32),
    to_unsigned(2009092274,32),
    to_unsigned(2009164979,32),
    to_unsigned(2009237666,32),
    to_unsigned(2009310335,32),
    to_unsigned(2009382985,32),
    to_unsigned(2009455616,32),
    to_unsigned(2009528229,32),
    to_unsigned(2009600824,32),
    to_unsigned(2009673400,32),
    to_unsigned(2009745958,32),
    to_unsigned(2009818497,32),
    to_unsigned(2009891018,32),
    to_unsigned(2009963520,32),
    to_unsigned(2010036004,32),
    to_unsigned(2010108469,32),
    to_unsigned(2010180916,32),
    to_unsigned(2010253345,32),
    to_unsigned(2010325755,32),
    to_unsigned(2010398146,32),
    to_unsigned(2010470519,32),
    to_unsigned(2010542873,32),
    to_unsigned(2010615209,32),
    to_unsigned(2010687527,32),
    to_unsigned(2010759826,32),
    to_unsigned(2010832107,32),
    to_unsigned(2010904369,32),
    to_unsigned(2010976612,32),
    to_unsigned(2011048837,32),
    to_unsigned(2011121044,32),
    to_unsigned(2011193232,32),
    to_unsigned(2011265402,32),
    to_unsigned(2011337553,32),
    to_unsigned(2011409686,32),
    to_unsigned(2011481800,32),
    to_unsigned(2011553895,32),
    to_unsigned(2011625973,32),
    to_unsigned(2011698031,32),
    to_unsigned(2011770072,32),
    to_unsigned(2011842093,32),
    to_unsigned(2011914097,32),
    to_unsigned(2011986081,32),
    to_unsigned(2012058048,32),
    to_unsigned(2012129995,32),
    to_unsigned(2012201925,32),
    to_unsigned(2012273835,32),
    to_unsigned(2012345728,32),
    to_unsigned(2012417601,32),
    to_unsigned(2012489457,32),
    to_unsigned(2012561293,32),
    to_unsigned(2012633112,32),
    to_unsigned(2012704911,32),
    to_unsigned(2012776693,32),
    to_unsigned(2012848456,32),
    to_unsigned(2012920200,32),
    to_unsigned(2012991926,32),
    to_unsigned(2013063633,32),
    to_unsigned(2013135322,32),
    to_unsigned(2013206992,32),
    to_unsigned(2013278644,32),
    to_unsigned(2013350277,32),
    to_unsigned(2013421892,32),
    to_unsigned(2013493488,32),
    to_unsigned(2013565066,32),
    to_unsigned(2013636625,32),
    to_unsigned(2013708165,32),
    to_unsigned(2013779688,32),
    to_unsigned(2013851191,32),
    to_unsigned(2013922677,32),
    to_unsigned(2013994143,32),
    to_unsigned(2014065591,32),
    to_unsigned(2014137021,32),
    to_unsigned(2014208432,32),
    to_unsigned(2014279825,32),
    to_unsigned(2014351199,32),
    to_unsigned(2014422554,32),
    to_unsigned(2014493892,32),
    to_unsigned(2014565210,32),
    to_unsigned(2014636510,32),
    to_unsigned(2014707792,32),
    to_unsigned(2014779055,32),
    to_unsigned(2014850299,32),
    to_unsigned(2014921525,32),
    to_unsigned(2014992733,32),
    to_unsigned(2015063921,32),
    to_unsigned(2015135092,32),
    to_unsigned(2015206244,32),
    to_unsigned(2015277377,32),
    to_unsigned(2015348492,32),
    to_unsigned(2015419588,32),
    to_unsigned(2015490666,32),
    to_unsigned(2015561725,32),
    to_unsigned(2015632766,32),
    to_unsigned(2015703788,32),
    to_unsigned(2015774792,32),
    to_unsigned(2015845777,32),
    to_unsigned(2015916744,32),
    to_unsigned(2015987692,32),
    to_unsigned(2016058621,32),
    to_unsigned(2016129532,32),
    to_unsigned(2016200425,32),
    to_unsigned(2016271299,32),
    to_unsigned(2016342154,32),
    to_unsigned(2016412991,32),
    to_unsigned(2016483809,32),
    to_unsigned(2016554609,32),
    to_unsigned(2016625390,32),
    to_unsigned(2016696153,32),
    to_unsigned(2016766897,32),
    to_unsigned(2016837623,32),
    to_unsigned(2016908330,32),
    to_unsigned(2016979019,32),
    to_unsigned(2017049689,32),
    to_unsigned(2017120340,32),
    to_unsigned(2017190973,32),
    to_unsigned(2017261588,32),
    to_unsigned(2017332184,32),
    to_unsigned(2017402761,32),
    to_unsigned(2017473320,32),
    to_unsigned(2017543860,32),
    to_unsigned(2017614382,32),
    to_unsigned(2017684885,32),
    to_unsigned(2017755369,32),
    to_unsigned(2017825836,32),
    to_unsigned(2017896283,32),
    to_unsigned(2017966712,32),
    to_unsigned(2018037122,32),
    to_unsigned(2018107514,32),
    to_unsigned(2018177888,32),
    to_unsigned(2018248242,32),
    to_unsigned(2018318579,32),
    to_unsigned(2018388896,32),
    to_unsigned(2018459195,32),
    to_unsigned(2018529476,32),
    to_unsigned(2018599738,32),
    to_unsigned(2018669982,32),
    to_unsigned(2018740206,32),
    to_unsigned(2018810413,32),
    to_unsigned(2018880601,32),
    to_unsigned(2018950770,32),
    to_unsigned(2019020921,32),
    to_unsigned(2019091053,32),
    to_unsigned(2019161166,32),
    to_unsigned(2019231261,32),
    to_unsigned(2019301338,32),
    to_unsigned(2019371396,32),
    to_unsigned(2019441435,32),
    to_unsigned(2019511456,32),
    to_unsigned(2019581458,32),
    to_unsigned(2019651441,32),
    to_unsigned(2019721407,32),
    to_unsigned(2019791353,32),
    to_unsigned(2019861281,32),
    to_unsigned(2019931190,32),
    to_unsigned(2020001081,32),
    to_unsigned(2020070953,32),
    to_unsigned(2020140807,32),
    to_unsigned(2020210642,32),
    to_unsigned(2020280459,32),
    to_unsigned(2020350257,32),
    to_unsigned(2020420036,32),
    to_unsigned(2020489797,32),
    to_unsigned(2020559539,32),
    to_unsigned(2020629263,32),
    to_unsigned(2020698968,32),
    to_unsigned(2020768654,32),
    to_unsigned(2020838322,32),
    to_unsigned(2020907972,32),
    to_unsigned(2020977602,32),
    to_unsigned(2021047215,32),
    to_unsigned(2021116808,32),
    to_unsigned(2021186383,32),
    to_unsigned(2021255940,32),
    to_unsigned(2021325478,32),
    to_unsigned(2021394997,32),
    to_unsigned(2021464498,32),
    to_unsigned(2021533980,32),
    to_unsigned(2021603444,32),
    to_unsigned(2021672889,32),
    to_unsigned(2021742315,32),
    to_unsigned(2021811723,32),
    to_unsigned(2021881112,32),
    to_unsigned(2021950483,32),
    to_unsigned(2022019835,32),
    to_unsigned(2022089169,32),
    to_unsigned(2022158483,32),
    to_unsigned(2022227780,32),
    to_unsigned(2022297057,32),
    to_unsigned(2022366317,32),
    to_unsigned(2022435557,32),
    to_unsigned(2022504779,32),
    to_unsigned(2022573983,32),
    to_unsigned(2022643167,32),
    to_unsigned(2022712334,32),
    to_unsigned(2022781481,32),
    to_unsigned(2022850610,32),
    to_unsigned(2022919721,32),
    to_unsigned(2022988812,32),
    to_unsigned(2023057886,32),
    to_unsigned(2023126940,32),
    to_unsigned(2023195976,32),
    to_unsigned(2023264994,32),
    to_unsigned(2023333993,32),
    to_unsigned(2023402973,32),
    to_unsigned(2023471935,32),
    to_unsigned(2023540878,32),
    to_unsigned(2023609802,32),
    to_unsigned(2023678708,32),
    to_unsigned(2023747595,32),
    to_unsigned(2023816464,32),
    to_unsigned(2023885314,32),
    to_unsigned(2023954145,32),
    to_unsigned(2024022958,32),
    to_unsigned(2024091752,32),
    to_unsigned(2024160528,32),
    to_unsigned(2024229285,32),
    to_unsigned(2024298023,32),
    to_unsigned(2024366743,32),
    to_unsigned(2024435444,32),
    to_unsigned(2024504127,32),
    to_unsigned(2024572791,32),
    to_unsigned(2024641436,32),
    to_unsigned(2024710063,32),
    to_unsigned(2024778671,32),
    to_unsigned(2024847261,32),
    to_unsigned(2024915832,32),
    to_unsigned(2024984384,32),
    to_unsigned(2025052918,32),
    to_unsigned(2025121433,32),
    to_unsigned(2025189929,32),
    to_unsigned(2025258407,32),
    to_unsigned(2025326866,32),
    to_unsigned(2025395307,32),
    to_unsigned(2025463729,32),
    to_unsigned(2025532132,32),
    to_unsigned(2025600517,32),
    to_unsigned(2025668883,32),
    to_unsigned(2025737231,32),
    to_unsigned(2025805560,32),
    to_unsigned(2025873870,32),
    to_unsigned(2025942162,32),
    to_unsigned(2026010435,32),
    to_unsigned(2026078689,32),
    to_unsigned(2026146925,32),
    to_unsigned(2026215142,32),
    to_unsigned(2026283341,32),
    to_unsigned(2026351521,32),
    to_unsigned(2026419682,32),
    to_unsigned(2026487825,32),
    to_unsigned(2026555949,32),
    to_unsigned(2026624054,32),
    to_unsigned(2026692141,32),
    to_unsigned(2026760209,32),
    to_unsigned(2026828259,32),
    to_unsigned(2026896290,32),
    to_unsigned(2026964302,32),
    to_unsigned(2027032296,32),
    to_unsigned(2027100271,32),
    to_unsigned(2027168227,32),
    to_unsigned(2027236165,32),
    to_unsigned(2027304084,32),
    to_unsigned(2027371984,32),
    to_unsigned(2027439866,32),
    to_unsigned(2027507729,32),
    to_unsigned(2027575574,32),
    to_unsigned(2027643400,32),
    to_unsigned(2027711207,32),
    to_unsigned(2027778996,32),
    to_unsigned(2027846766,32),
    to_unsigned(2027914517,32),
    to_unsigned(2027982250,32),
    to_unsigned(2028049964,32),
    to_unsigned(2028117660,32),
    to_unsigned(2028185336,32),
    to_unsigned(2028252995,32),
    to_unsigned(2028320634,32),
    to_unsigned(2028388255,32),
    to_unsigned(2028455857,32),
    to_unsigned(2028523441,32),
    to_unsigned(2028591006,32),
    to_unsigned(2028658552,32),
    to_unsigned(2028726080,32),
    to_unsigned(2028793589,32),
    to_unsigned(2028861079,32),
    to_unsigned(2028928551,32),
    to_unsigned(2028996004,32),
    to_unsigned(2029063438,32),
    to_unsigned(2029130854,32),
    to_unsigned(2029198251,32),
    to_unsigned(2029265630,32),
    to_unsigned(2029332990,32),
    to_unsigned(2029400331,32),
    to_unsigned(2029467653,32),
    to_unsigned(2029534957,32),
    to_unsigned(2029602242,32),
    to_unsigned(2029669509,32),
    to_unsigned(2029736757,32),
    to_unsigned(2029803986,32),
    to_unsigned(2029871196,32),
    to_unsigned(2029938388,32),
    to_unsigned(2030005562,32),
    to_unsigned(2030072716,32),
    to_unsigned(2030139852,32),
    to_unsigned(2030206969,32),
    to_unsigned(2030274068,32),
    to_unsigned(2030341148,32),
    to_unsigned(2030408209,32),
    to_unsigned(2030475252,32),
    to_unsigned(2030542276,32),
    to_unsigned(2030609281,32),
    to_unsigned(2030676268,32),
    to_unsigned(2030743236,32),
    to_unsigned(2030810185,32),
    to_unsigned(2030877116,32),
    to_unsigned(2030944028,32),
    to_unsigned(2031010921,32),
    to_unsigned(2031077796,32),
    to_unsigned(2031144651,32),
    to_unsigned(2031211489,32),
    to_unsigned(2031278307,32),
    to_unsigned(2031345107,32),
    to_unsigned(2031411889,32),
    to_unsigned(2031478651,32),
    to_unsigned(2031545395,32),
    to_unsigned(2031612120,32),
    to_unsigned(2031678827,32),
    to_unsigned(2031745515,32),
    to_unsigned(2031812184,32),
    to_unsigned(2031878835,32),
    to_unsigned(2031945467,32),
    to_unsigned(2032012080,32),
    to_unsigned(2032078674,32),
    to_unsigned(2032145250,32),
    to_unsigned(2032211807,32),
    to_unsigned(2032278346,32),
    to_unsigned(2032344866,32),
    to_unsigned(2032411367,32),
    to_unsigned(2032477849,32),
    to_unsigned(2032544313,32),
    to_unsigned(2032610758,32),
    to_unsigned(2032677184,32),
    to_unsigned(2032743592,32),
    to_unsigned(2032809981,32),
    to_unsigned(2032876351,32),
    to_unsigned(2032942703,32),
    to_unsigned(2033009036,32),
    to_unsigned(2033075350,32),
    to_unsigned(2033141646,32),
    to_unsigned(2033207923,32),
    to_unsigned(2033274181,32),
    to_unsigned(2033340421,32),
    to_unsigned(2033406641,32),
    to_unsigned(2033472844,32),
    to_unsigned(2033539027,32),
    to_unsigned(2033605192,32),
    to_unsigned(2033671338,32),
    to_unsigned(2033737465,32),
    to_unsigned(2033803574,32),
    to_unsigned(2033869664,32),
    to_unsigned(2033935735,32),
    to_unsigned(2034001788,32),
    to_unsigned(2034067822,32),
    to_unsigned(2034133837,32),
    to_unsigned(2034199833,32),
    to_unsigned(2034265811,32),
    to_unsigned(2034331770,32),
    to_unsigned(2034397711,32),
    to_unsigned(2034463632,32),
    to_unsigned(2034529535,32),
    to_unsigned(2034595420,32),
    to_unsigned(2034661285,32),
    to_unsigned(2034727132,32),
    to_unsigned(2034792961,32),
    to_unsigned(2034858770,32),
    to_unsigned(2034924561,32),
    to_unsigned(2034990333,32),
    to_unsigned(2035056086,32),
    to_unsigned(2035121821,32),
    to_unsigned(2035187537,32),
    to_unsigned(2035253234,32),
    to_unsigned(2035318913,32),
    to_unsigned(2035384573,32),
    to_unsigned(2035450214,32),
    to_unsigned(2035515836,32),
    to_unsigned(2035581440,32),
    to_unsigned(2035647025,32),
    to_unsigned(2035712591,32),
    to_unsigned(2035778139,32),
    to_unsigned(2035843668,32),
    to_unsigned(2035909178,32),
    to_unsigned(2035974669,32),
    to_unsigned(2036040142,32),
    to_unsigned(2036105596,32),
    to_unsigned(2036171031,32),
    to_unsigned(2036236448,32),
    to_unsigned(2036301846,32),
    to_unsigned(2036367225,32),
    to_unsigned(2036432586,32),
    to_unsigned(2036497927,32),
    to_unsigned(2036563250,32),
    to_unsigned(2036628555,32),
    to_unsigned(2036693840,32),
    to_unsigned(2036759107,32),
    to_unsigned(2036824355,32),
    to_unsigned(2036889584,32),
    to_unsigned(2036954795,32),
    to_unsigned(2037019987,32),
    to_unsigned(2037085160,32),
    to_unsigned(2037150315,32),
    to_unsigned(2037215451,32),
    to_unsigned(2037280568,32),
    to_unsigned(2037345666,32),
    to_unsigned(2037410746,32),
    to_unsigned(2037475806,32),
    to_unsigned(2037540849,32),
    to_unsigned(2037605872,32),
    to_unsigned(2037670877,32),
    to_unsigned(2037735863,32),
    to_unsigned(2037800830,32),
    to_unsigned(2037865778,32),
    to_unsigned(2037930708,32),
    to_unsigned(2037995619,32),
    to_unsigned(2038060512,32),
    to_unsigned(2038125385,32),
    to_unsigned(2038190240,32),
    to_unsigned(2038255076,32),
    to_unsigned(2038319893,32),
    to_unsigned(2038384692,32),
    to_unsigned(2038449472,32),
    to_unsigned(2038514233,32),
    to_unsigned(2038578975,32),
    to_unsigned(2038643699,32),
    to_unsigned(2038708404,32),
    to_unsigned(2038773090,32),
    to_unsigned(2038837758,32),
    to_unsigned(2038902406,32),
    to_unsigned(2038967036,32),
    to_unsigned(2039031648,32),
    to_unsigned(2039096240,32),
    to_unsigned(2039160814,32),
    to_unsigned(2039225369,32),
    to_unsigned(2039289905,32),
    to_unsigned(2039354423,32),
    to_unsigned(2039418922,32),
    to_unsigned(2039483402,32),
    to_unsigned(2039547863,32),
    to_unsigned(2039612305,32),
    to_unsigned(2039676729,32),
    to_unsigned(2039741134,32),
    to_unsigned(2039805520,32),
    to_unsigned(2039869888,32),
    to_unsigned(2039934237,32),
    to_unsigned(2039998567,32),
    to_unsigned(2040062878,32),
    to_unsigned(2040127171,32),
    to_unsigned(2040191444,32),
    to_unsigned(2040255699,32),
    to_unsigned(2040319936,32),
    to_unsigned(2040384153,32),
    to_unsigned(2040448352,32),
    to_unsigned(2040512532,32),
    to_unsigned(2040576693,32),
    to_unsigned(2040640836,32),
    to_unsigned(2040704960,32),
    to_unsigned(2040769065,32),
    to_unsigned(2040833151,32),
    to_unsigned(2040897218,32),
    to_unsigned(2040961267,32),
    to_unsigned(2041025297,32),
    to_unsigned(2041089308,32),
    to_unsigned(2041153301,32),
    to_unsigned(2041217274,32),
    to_unsigned(2041281229,32),
    to_unsigned(2041345165,32),
    to_unsigned(2041409083,32),
    to_unsigned(2041472981,32),
    to_unsigned(2041536861,32),
    to_unsigned(2041600722,32),
    to_unsigned(2041664564,32),
    to_unsigned(2041728388,32),
    to_unsigned(2041792193,32),
    to_unsigned(2041855979,32),
    to_unsigned(2041919746,32),
    to_unsigned(2041983495,32),
    to_unsigned(2042047224,32),
    to_unsigned(2042110935,32),
    to_unsigned(2042174627,32),
    to_unsigned(2042238301,32),
    to_unsigned(2042301955,32),
    to_unsigned(2042365591,32),
    to_unsigned(2042429208,32),
    to_unsigned(2042492807,32),
    to_unsigned(2042556386,32),
    to_unsigned(2042619947,32),
    to_unsigned(2042683489,32),
    to_unsigned(2042747012,32),
    to_unsigned(2042810516,32),
    to_unsigned(2042874002,32),
    to_unsigned(2042937469,32),
    to_unsigned(2043000917,32),
    to_unsigned(2043064346,32),
    to_unsigned(2043127757,32),
    to_unsigned(2043191149,32),
    to_unsigned(2043254522,32),
    to_unsigned(2043317876,32),
    to_unsigned(2043381211,32),
    to_unsigned(2043444528,32),
    to_unsigned(2043507826,32),
    to_unsigned(2043571105,32),
    to_unsigned(2043634365,32),
    to_unsigned(2043697607,32),
    to_unsigned(2043760829,32),
    to_unsigned(2043824033,32),
    to_unsigned(2043887218,32),
    to_unsigned(2043950385,32),
    to_unsigned(2044013532,32),
    to_unsigned(2044076661,32),
    to_unsigned(2044139771,32),
    to_unsigned(2044202862,32),
    to_unsigned(2044265935,32),
    to_unsigned(2044328988,32),
    to_unsigned(2044392023,32),
    to_unsigned(2044455039,32),
    to_unsigned(2044518036,32),
    to_unsigned(2044581015,32),
    to_unsigned(2044643975,32),
    to_unsigned(2044706915,32),
    to_unsigned(2044769837,32),
    to_unsigned(2044832741,32),
    to_unsigned(2044895625,32),
    to_unsigned(2044958491,32),
    to_unsigned(2045021338,32),
    to_unsigned(2045084166,32),
    to_unsigned(2045146975,32),
    to_unsigned(2045209766,32),
    to_unsigned(2045272537,32),
    to_unsigned(2045335290,32),
    to_unsigned(2045398024,32),
    to_unsigned(2045460740,32),
    to_unsigned(2045523436,32),
    to_unsigned(2045586114,32),
    to_unsigned(2045648773,32),
    to_unsigned(2045711413,32),
    to_unsigned(2045774034,32),
    to_unsigned(2045836636,32),
    to_unsigned(2045899220,32),
    to_unsigned(2045961785,32),
    to_unsigned(2046024331,32),
    to_unsigned(2046086858,32),
    to_unsigned(2046149367,32),
    to_unsigned(2046211856,32),
    to_unsigned(2046274327,32),
    to_unsigned(2046336779,32),
    to_unsigned(2046399212,32),
    to_unsigned(2046461627,32),
    to_unsigned(2046524022,32),
    to_unsigned(2046586399,32),
    to_unsigned(2046648757,32),
    to_unsigned(2046711096,32),
    to_unsigned(2046773417,32),
    to_unsigned(2046835718,32),
    to_unsigned(2046898001,32),
    to_unsigned(2046960265,32),
    to_unsigned(2047022510,32),
    to_unsigned(2047084736,32),
    to_unsigned(2047146944,32),
    to_unsigned(2047209132,32),
    to_unsigned(2047271302,32),
    to_unsigned(2047333453,32),
    to_unsigned(2047395585,32),
    to_unsigned(2047457699,32),
    to_unsigned(2047519793,32),
    to_unsigned(2047581869,32),
    to_unsigned(2047643926,32),
    to_unsigned(2047705964,32),
    to_unsigned(2047767983,32),
    to_unsigned(2047829984,32),
    to_unsigned(2047891965,32),
    to_unsigned(2047953928,32),
    to_unsigned(2048015872,32),
    to_unsigned(2048077797,32),
    to_unsigned(2048139703,32),
    to_unsigned(2048201591,32),
    to_unsigned(2048263459,32),
    to_unsigned(2048325309,32),
    to_unsigned(2048387140,32),
    to_unsigned(2048448952,32),
    to_unsigned(2048510746,32),
    to_unsigned(2048572520,32),
    to_unsigned(2048634276,32),
    to_unsigned(2048696013,32),
    to_unsigned(2048757731,32),
    to_unsigned(2048819430,32),
    to_unsigned(2048881110,32),
    to_unsigned(2048942772,32),
    to_unsigned(2049004415,32),
    to_unsigned(2049066039,32),
    to_unsigned(2049127644,32),
    to_unsigned(2049189230,32),
    to_unsigned(2049250797,32),
    to_unsigned(2049312346,32),
    to_unsigned(2049373875,32),
    to_unsigned(2049435386,32),
    to_unsigned(2049496878,32),
    to_unsigned(2049558351,32),
    to_unsigned(2049619806,32),
    to_unsigned(2049681241,32),
    to_unsigned(2049742658,32),
    to_unsigned(2049804056,32),
    to_unsigned(2049865435,32),
    to_unsigned(2049926795,32),
    to_unsigned(2049988136,32),
    to_unsigned(2050049458,32),
    to_unsigned(2050110762,32),
    to_unsigned(2050172047,32),
    to_unsigned(2050233313,32),
    to_unsigned(2050294560,32),
    to_unsigned(2050355788,32),
    to_unsigned(2050416997,32),
    to_unsigned(2050478188,32),
    to_unsigned(2050539360,32),
    to_unsigned(2050600512,32),
    to_unsigned(2050661646,32),
    to_unsigned(2050722761,32),
    to_unsigned(2050783858,32),
    to_unsigned(2050844935,32),
    to_unsigned(2050905994,32),
    to_unsigned(2050967033,32),
    to_unsigned(2051028054,32),
    to_unsigned(2051089056,32),
    to_unsigned(2051150040,32),
    to_unsigned(2051211004,32),
    to_unsigned(2051271949,32),
    to_unsigned(2051332876,32),
    to_unsigned(2051393784,32),
    to_unsigned(2051454673,32),
    to_unsigned(2051515543,32),
    to_unsigned(2051576394,32),
    to_unsigned(2051637226,32),
    to_unsigned(2051698040,32),
    to_unsigned(2051758834,32),
    to_unsigned(2051819610,32),
    to_unsigned(2051880367,32),
    to_unsigned(2051941105,32),
    to_unsigned(2052001824,32),
    to_unsigned(2052062524,32),
    to_unsigned(2052123206,32),
    to_unsigned(2052183868,32),
    to_unsigned(2052244512,32),
    to_unsigned(2052305137,32),
    to_unsigned(2052365743,32),
    to_unsigned(2052426330,32),
    to_unsigned(2052486898,32),
    to_unsigned(2052547448,32),
    to_unsigned(2052607978,32),
    to_unsigned(2052668490,32),
    to_unsigned(2052728983,32),
    to_unsigned(2052789457,32),
    to_unsigned(2052849912,32),
    to_unsigned(2052910348,32),
    to_unsigned(2052970765,32),
    to_unsigned(2053031163,32),
    to_unsigned(2053091543,32),
    to_unsigned(2053151904,32),
    to_unsigned(2053212246,32),
    to_unsigned(2053272569,32),
    to_unsigned(2053332873,32),
    to_unsigned(2053393158,32),
    to_unsigned(2053453424,32),
    to_unsigned(2053513672,32),
    to_unsigned(2053573900,32),
    to_unsigned(2053634110,32),
    to_unsigned(2053694301,32),
    to_unsigned(2053754473,32),
    to_unsigned(2053814626,32),
    to_unsigned(2053874760,32),
    to_unsigned(2053934875,32),
    to_unsigned(2053994972,32),
    to_unsigned(2054055049,32),
    to_unsigned(2054115108,32),
    to_unsigned(2054175148,32),
    to_unsigned(2054235169,32),
    to_unsigned(2054295171,32),
    to_unsigned(2054355154,32),
    to_unsigned(2054415118,32),
    to_unsigned(2054475064,32),
    to_unsigned(2054534990,32),
    to_unsigned(2054594898,32),
    to_unsigned(2054654786,32),
    to_unsigned(2054714656,32),
    to_unsigned(2054774507,32),
    to_unsigned(2054834339,32),
    to_unsigned(2054894152,32),
    to_unsigned(2054953947,32),
    to_unsigned(2055013722,32),
    to_unsigned(2055073479,32),
    to_unsigned(2055133216,32),
    to_unsigned(2055192935,32),
    to_unsigned(2055252635,32),
    to_unsigned(2055312316,32),
    to_unsigned(2055371978,32),
    to_unsigned(2055431621,32),
    to_unsigned(2055491245,32),
    to_unsigned(2055550851,32),
    to_unsigned(2055610437,32),
    to_unsigned(2055670005,32),
    to_unsigned(2055729554,32),
    to_unsigned(2055789083,32),
    to_unsigned(2055848594,32),
    to_unsigned(2055908086,32),
    to_unsigned(2055967559,32),
    to_unsigned(2056027014,32),
    to_unsigned(2056086449,32),
    to_unsigned(2056145865,32),
    to_unsigned(2056205263,32),
    to_unsigned(2056264641,32),
    to_unsigned(2056324001,32),
    to_unsigned(2056383342,32),
    to_unsigned(2056442664,32),
    to_unsigned(2056501967,32),
    to_unsigned(2056561251,32),
    to_unsigned(2056620516,32),
    to_unsigned(2056679762,32),
    to_unsigned(2056738990,32),
    to_unsigned(2056798198,32),
    to_unsigned(2056857388,32),
    to_unsigned(2056916559,32),
    to_unsigned(2056975710,32),
    to_unsigned(2057034843,32),
    to_unsigned(2057093957,32),
    to_unsigned(2057153052,32),
    to_unsigned(2057212128,32),
    to_unsigned(2057271186,32),
    to_unsigned(2057330224,32),
    to_unsigned(2057389243,32),
    to_unsigned(2057448244,32),
    to_unsigned(2057507225,32),
    to_unsigned(2057566188,32),
    to_unsigned(2057625132,32),
    to_unsigned(2057684057,32),
    to_unsigned(2057742963,32),
    to_unsigned(2057801850,32),
    to_unsigned(2057860718,32),
    to_unsigned(2057919567,32),
    to_unsigned(2057978397,32),
    to_unsigned(2058037209,32),
    to_unsigned(2058096001,32),
    to_unsigned(2058154775,32),
    to_unsigned(2058213529,32),
    to_unsigned(2058272265,32),
    to_unsigned(2058330982,32),
    to_unsigned(2058389680,32),
    to_unsigned(2058448358,32),
    to_unsigned(2058507018,32),
    to_unsigned(2058565660,32),
    to_unsigned(2058624282,32),
    to_unsigned(2058682885,32),
    to_unsigned(2058741469,32),
    to_unsigned(2058800035,32),
    to_unsigned(2058858581,32),
    to_unsigned(2058917109,32),
    to_unsigned(2058975617,32),
    to_unsigned(2059034107,32),
    to_unsigned(2059092578,32),
    to_unsigned(2059151030,32),
    to_unsigned(2059209463,32),
    to_unsigned(2059267877,32),
    to_unsigned(2059326272,32),
    to_unsigned(2059384648,32),
    to_unsigned(2059443005,32),
    to_unsigned(2059501343,32),
    to_unsigned(2059559663,32),
    to_unsigned(2059617963,32),
    to_unsigned(2059676244,32),
    to_unsigned(2059734507,32),
    to_unsigned(2059792751,32),
    to_unsigned(2059850975,32),
    to_unsigned(2059909181,32),
    to_unsigned(2059967368,32),
    to_unsigned(2060025536,32),
    to_unsigned(2060083685,32),
    to_unsigned(2060141815,32),
    to_unsigned(2060199926,32),
    to_unsigned(2060258018,32),
    to_unsigned(2060316091,32),
    to_unsigned(2060374145,32),
    to_unsigned(2060432181,32),
    to_unsigned(2060490197,32),
    to_unsigned(2060548194,32),
    to_unsigned(2060606173,32),
    to_unsigned(2060664132,32),
    to_unsigned(2060722073,32),
    to_unsigned(2060779995,32),
    to_unsigned(2060837897,32),
    to_unsigned(2060895781,32),
    to_unsigned(2060953646,32),
    to_unsigned(2061011492,32),
    to_unsigned(2061069319,32),
    to_unsigned(2061127127,32),
    to_unsigned(2061184916,32),
    to_unsigned(2061242686,32),
    to_unsigned(2061300437,32),
    to_unsigned(2061358170,32),
    to_unsigned(2061415883,32),
    to_unsigned(2061473577,32),
    to_unsigned(2061531253,32),
    to_unsigned(2061588909,32),
    to_unsigned(2061646547,32),
    to_unsigned(2061704165,32),
    to_unsigned(2061761765,32),
    to_unsigned(2061819345,32),
    to_unsigned(2061876907,32),
    to_unsigned(2061934450,32),
    to_unsigned(2061991973,32),
    to_unsigned(2062049478,32),
    to_unsigned(2062106964,32),
    to_unsigned(2062164431,32),
    to_unsigned(2062221879,32),
    to_unsigned(2062279308,32),
    to_unsigned(2062336718,32),
    to_unsigned(2062394109,32),
    to_unsigned(2062451481,32),
    to_unsigned(2062508835,32),
    to_unsigned(2062566169,32),
    to_unsigned(2062623484,32),
    to_unsigned(2062680780,32),
    to_unsigned(2062738058,32),
    to_unsigned(2062795316,32),
    to_unsigned(2062852555,32),
    to_unsigned(2062909776,32),
    to_unsigned(2062966977,32),
    to_unsigned(2063024160,32),
    to_unsigned(2063081324,32),
    to_unsigned(2063138468,32),
    to_unsigned(2063195594,32),
    to_unsigned(2063252700,32),
    to_unsigned(2063309788,32),
    to_unsigned(2063366857,32),
    to_unsigned(2063423907,32),
    to_unsigned(2063480938,32),
    to_unsigned(2063537949,32),
    to_unsigned(2063594942,32),
    to_unsigned(2063651916,32),
    to_unsigned(2063708871,32),
    to_unsigned(2063765807,32),
    to_unsigned(2063822724,32),
    to_unsigned(2063879622,32),
    to_unsigned(2063936501,32),
    to_unsigned(2063993361,32),
    to_unsigned(2064050202,32),
    to_unsigned(2064107025,32),
    to_unsigned(2064163828,32),
    to_unsigned(2064220612,32),
    to_unsigned(2064277377,32),
    to_unsigned(2064334123,32),
    to_unsigned(2064390851,32),
    to_unsigned(2064447559,32),
    to_unsigned(2064504248,32),
    to_unsigned(2064560919,32),
    to_unsigned(2064617570,32),
    to_unsigned(2064674203,32),
    to_unsigned(2064730816,32),
    to_unsigned(2064787410,32),
    to_unsigned(2064843986,32),
    to_unsigned(2064900542,32),
    to_unsigned(2064957080,32),
    to_unsigned(2065013598,32),
    to_unsigned(2065070098,32),
    to_unsigned(2065126578,32),
    to_unsigned(2065183040,32),
    to_unsigned(2065239483,32),
    to_unsigned(2065295906,32),
    to_unsigned(2065352311,32),
    to_unsigned(2065408697,32),
    to_unsigned(2065465063,32),
    to_unsigned(2065521411,32),
    to_unsigned(2065577740,32),
    to_unsigned(2065634049,32),
    to_unsigned(2065690340,32),
    to_unsigned(2065746612,32),
    to_unsigned(2065802864,32),
    to_unsigned(2065859098,32),
    to_unsigned(2065915313,32),
    to_unsigned(2065971509,32),
    to_unsigned(2066027686,32),
    to_unsigned(2066083843,32),
    to_unsigned(2066139982,32),
    to_unsigned(2066196102,32),
    to_unsigned(2066252203,32),
    to_unsigned(2066308285,32),
    to_unsigned(2066364347,32),
    to_unsigned(2066420391,32),
    to_unsigned(2066476416,32),
    to_unsigned(2066532422,32),
    to_unsigned(2066588409,32),
    to_unsigned(2066644377,32),
    to_unsigned(2066700325,32),
    to_unsigned(2066756255,32),
    to_unsigned(2066812166,32),
    to_unsigned(2066868058,32),
    to_unsigned(2066923931,32),
    to_unsigned(2066979785,32),
    to_unsigned(2067035620,32),
    to_unsigned(2067091436,32),
    to_unsigned(2067147232,32),
    to_unsigned(2067203010,32),
    to_unsigned(2067258769,32),
    to_unsigned(2067314509,32),
    to_unsigned(2067370230,32),
    to_unsigned(2067425932,32),
    to_unsigned(2067481615,32),
    to_unsigned(2067537279,32),
    to_unsigned(2067592923,32),
    to_unsigned(2067648549,32),
    to_unsigned(2067704156,32),
    to_unsigned(2067759744,32),
    to_unsigned(2067815313,32),
    to_unsigned(2067870863,32),
    to_unsigned(2067926393,32),
    to_unsigned(2067981905,32),
    to_unsigned(2068037398,32),
    to_unsigned(2068092872,32),
    to_unsigned(2068148327,32),
    to_unsigned(2068203762,32),
    to_unsigned(2068259179,32),
    to_unsigned(2068314577,32),
    to_unsigned(2068369956,32),
    to_unsigned(2068425315,32),
    to_unsigned(2068480656,32),
    to_unsigned(2068535978,32),
    to_unsigned(2068591280,32),
    to_unsigned(2068646564,32),
    to_unsigned(2068701829,32),
    to_unsigned(2068757074,32),
    to_unsigned(2068812301,32),
    to_unsigned(2068867509,32),
    to_unsigned(2068922697,32),
    to_unsigned(2068977867,32),
    to_unsigned(2069033017,32),
    to_unsigned(2069088149,32),
    to_unsigned(2069143262,32),
    to_unsigned(2069198355,32),
    to_unsigned(2069253430,32),
    to_unsigned(2069308485,32),
    to_unsigned(2069363521,32),
    to_unsigned(2069418539,32),
    to_unsigned(2069473537,32),
    to_unsigned(2069528517,32),
    to_unsigned(2069583477,32),
    to_unsigned(2069638418,32),
    to_unsigned(2069693341,32),
    to_unsigned(2069748244,32),
    to_unsigned(2069803128,32),
    to_unsigned(2069857993,32),
    to_unsigned(2069912840,32),
    to_unsigned(2069967667,32),
    to_unsigned(2070022475,32),
    to_unsigned(2070077264,32),
    to_unsigned(2070132034,32),
    to_unsigned(2070186785,32),
    to_unsigned(2070241517,32),
    to_unsigned(2070296230,32),
    to_unsigned(2070350924,32),
    to_unsigned(2070405599,32),
    to_unsigned(2070460255,32),
    to_unsigned(2070514892,32),
    to_unsigned(2070569510,32),
    to_unsigned(2070624109,32),
    to_unsigned(2070678689,32),
    to_unsigned(2070733249,32),
    to_unsigned(2070787791,32),
    to_unsigned(2070842314,32),
    to_unsigned(2070896818,32),
    to_unsigned(2070951302,32),
    to_unsigned(2071005768,32),
    to_unsigned(2071060214,32),
    to_unsigned(2071114642,32),
    to_unsigned(2071169050,32),
    to_unsigned(2071223440,32),
    to_unsigned(2071277810,32),
    to_unsigned(2071332162,32),
    to_unsigned(2071386494,32),
    to_unsigned(2071440807,32),
    to_unsigned(2071495101,32),
    to_unsigned(2071549377,32),
    to_unsigned(2071603633,32),
    to_unsigned(2071657870,32),
    to_unsigned(2071712088,32),
    to_unsigned(2071766287,32),
    to_unsigned(2071820467,32),
    to_unsigned(2071874628,32),
    to_unsigned(2071928770,32),
    to_unsigned(2071982893,32),
    to_unsigned(2072036997,32),
    to_unsigned(2072091081,32),
    to_unsigned(2072145147,32),
    to_unsigned(2072199194,32),
    to_unsigned(2072253221,32),
    to_unsigned(2072307230,32),
    to_unsigned(2072361220,32),
    to_unsigned(2072415190,32),
    to_unsigned(2072469141,32),
    to_unsigned(2072523074,32),
    to_unsigned(2072576987,32),
    to_unsigned(2072630881,32),
    to_unsigned(2072684757,32),
    to_unsigned(2072738613,32),
    to_unsigned(2072792450,32),
    to_unsigned(2072846268,32),
    to_unsigned(2072900067,32),
    to_unsigned(2072953847,32),
    to_unsigned(2073007608,32),
    to_unsigned(2073061350,32),
    to_unsigned(2073115073,32),
    to_unsigned(2073168776,32),
    to_unsigned(2073222461,32),
    to_unsigned(2073276127,32),
    to_unsigned(2073329773,32),
    to_unsigned(2073383401,32),
    to_unsigned(2073437009,32),
    to_unsigned(2073490599,32),
    to_unsigned(2073544169,32),
    to_unsigned(2073597720,32),
    to_unsigned(2073651253,32),
    to_unsigned(2073704766,32),
    to_unsigned(2073758260,32),
    to_unsigned(2073811735,32),
    to_unsigned(2073865191,32),
    to_unsigned(2073918628,32),
    to_unsigned(2073972046,32),
    to_unsigned(2074025445,32),
    to_unsigned(2074078824,32),
    to_unsigned(2074132185,32),
    to_unsigned(2074185527,32),
    to_unsigned(2074238849,32),
    to_unsigned(2074292153,32),
    to_unsigned(2074345437,32),
    to_unsigned(2074398702,32),
    to_unsigned(2074451949,32),
    to_unsigned(2074505176,32),
    to_unsigned(2074558384,32),
    to_unsigned(2074611573,32),
    to_unsigned(2074664743,32),
    to_unsigned(2074717894,32),
    to_unsigned(2074771026,32),
    to_unsigned(2074824139,32),
    to_unsigned(2074877232,32),
    to_unsigned(2074930307,32),
    to_unsigned(2074983363,32),
    to_unsigned(2075036399,32),
    to_unsigned(2075089416,32),
    to_unsigned(2075142415,32),
    to_unsigned(2075195394,32),
    to_unsigned(2075248354,32),
    to_unsigned(2075301295,32),
    to_unsigned(2075354217,32),
    to_unsigned(2075407120,32),
    to_unsigned(2075460004,32),
    to_unsigned(2075512869,32),
    to_unsigned(2075565715,32),
    to_unsigned(2075618542,32),
    to_unsigned(2075671349,32),
    to_unsigned(2075724138,32),
    to_unsigned(2075776907,32),
    to_unsigned(2075829657,32),
    to_unsigned(2075882389,32),
    to_unsigned(2075935101,32),
    to_unsigned(2075987794,32),
    to_unsigned(2076040468,32),
    to_unsigned(2076093123,32),
    to_unsigned(2076145759,32),
    to_unsigned(2076198376,32),
    to_unsigned(2076250973,32),
    to_unsigned(2076303552,32),
    to_unsigned(2076356111,32),
    to_unsigned(2076408652,32),
    to_unsigned(2076461173,32),
    to_unsigned(2076513675,32),
    to_unsigned(2076566159,32),
    to_unsigned(2076618623,32),
    to_unsigned(2076671068,32),
    to_unsigned(2076723494,32),
    to_unsigned(2076775900,32),
    to_unsigned(2076828288,32),
    to_unsigned(2076880657,32),
    to_unsigned(2076933006,32),
    to_unsigned(2076985337,32),
    to_unsigned(2077037648,32),
    to_unsigned(2077089940,32),
    to_unsigned(2077142214,32),
    to_unsigned(2077194468,32),
    to_unsigned(2077246703,32),
    to_unsigned(2077298919,32),
    to_unsigned(2077351115,32),
    to_unsigned(2077403293,32),
    to_unsigned(2077455452,32),
    to_unsigned(2077507591,32),
    to_unsigned(2077559712,32),
    to_unsigned(2077611813,32),
    to_unsigned(2077663895,32),
    to_unsigned(2077715959,32),
    to_unsigned(2077768003,32),
    to_unsigned(2077820028,32),
    to_unsigned(2077872033,32),
    to_unsigned(2077924020,32),
    to_unsigned(2077975988,32),
    to_unsigned(2078027936,32),
    to_unsigned(2078079866,32),
    to_unsigned(2078131776,32),
    to_unsigned(2078183667,32),
    to_unsigned(2078235539,32),
    to_unsigned(2078287393,32),
    to_unsigned(2078339226,32),
    to_unsigned(2078391041,32),
    to_unsigned(2078442837,32),
    to_unsigned(2078494614,32),
    to_unsigned(2078546371,32),
    to_unsigned(2078598110,32),
    to_unsigned(2078649829,32),
    to_unsigned(2078701529,32),
    to_unsigned(2078753210,32),
    to_unsigned(2078804872,32),
    to_unsigned(2078856515,32),
    to_unsigned(2078908139,32),
    to_unsigned(2078959743,32),
    to_unsigned(2079011329,32),
    to_unsigned(2079062895,32),
    to_unsigned(2079114443,32),
    to_unsigned(2079165971,32),
    to_unsigned(2079217480,32),
    to_unsigned(2079268970,32),
    to_unsigned(2079320441,32),
    to_unsigned(2079371893,32),
    to_unsigned(2079423325,32),
    to_unsigned(2079474739,32),
    to_unsigned(2079526133,32),
    to_unsigned(2079577509,32),
    to_unsigned(2079628865,32),
    to_unsigned(2079680202,32),
    to_unsigned(2079731520,32),
    to_unsigned(2079782819,32),
    to_unsigned(2079834099,32),
    to_unsigned(2079885359,32),
    to_unsigned(2079936601,32),
    to_unsigned(2079987823,32),
    to_unsigned(2080039026,32),
    to_unsigned(2080090211,32),
    to_unsigned(2080141376,32),
    to_unsigned(2080192521,32),
    to_unsigned(2080243648,32),
    to_unsigned(2080294756,32),
    to_unsigned(2080345844,32),
    to_unsigned(2080396914,32),
    to_unsigned(2080447964,32),
    to_unsigned(2080498995,32),
    to_unsigned(2080550007,32),
    to_unsigned(2080601000,32),
    to_unsigned(2080651974,32),
    to_unsigned(2080702929,32),
    to_unsigned(2080753864,32),
    to_unsigned(2080804781,32),
    to_unsigned(2080855678,32),
    to_unsigned(2080906556,32),
    to_unsigned(2080957415,32),
    to_unsigned(2081008255,32),
    to_unsigned(2081059076,32),
    to_unsigned(2081109878,32),
    to_unsigned(2081160660,32),
    to_unsigned(2081211424,32),
    to_unsigned(2081262168,32),
    to_unsigned(2081312893,32),
    to_unsigned(2081363599,32),
    to_unsigned(2081414286,32),
    to_unsigned(2081464954,32),
    to_unsigned(2081515602,32),
    to_unsigned(2081566232,32),
    to_unsigned(2081616842,32),
    to_unsigned(2081667433,32),
    to_unsigned(2081718005,32),
    to_unsigned(2081768558,32),
    to_unsigned(2081819092,32),
    to_unsigned(2081869607,32),
    to_unsigned(2081920102,32),
    to_unsigned(2081970579,32),
    to_unsigned(2082021036,32),
    to_unsigned(2082071474,32),
    to_unsigned(2082121893,32),
    to_unsigned(2082172293,32),
    to_unsigned(2082222674,32),
    to_unsigned(2082273035,32),
    to_unsigned(2082323378,32),
    to_unsigned(2082373701,32),
    to_unsigned(2082424005,32),
    to_unsigned(2082474290,32),
    to_unsigned(2082524556,32),
    to_unsigned(2082574803,32),
    to_unsigned(2082625030,32),
    to_unsigned(2082675239,32),
    to_unsigned(2082725428,32),
    to_unsigned(2082775598,32),
    to_unsigned(2082825749,32),
    to_unsigned(2082875881,32),
    to_unsigned(2082925994,32),
    to_unsigned(2082976087,32),
    to_unsigned(2083026162,32),
    to_unsigned(2083076217,32),
    to_unsigned(2083126253,32),
    to_unsigned(2083176270,32),
    to_unsigned(2083226268,32),
    to_unsigned(2083276247,32),
    to_unsigned(2083326206,32),
    to_unsigned(2083376147,32),
    to_unsigned(2083426068,32),
    to_unsigned(2083475970,32),
    to_unsigned(2083525853,32),
    to_unsigned(2083575717,32),
    to_unsigned(2083625561,32),
    to_unsigned(2083675387,32),
    to_unsigned(2083725193,32),
    to_unsigned(2083774980,32),
    to_unsigned(2083824748,32),
    to_unsigned(2083874497,32),
    to_unsigned(2083924227,32),
    to_unsigned(2083973938,32),
    to_unsigned(2084023629,32),
    to_unsigned(2084073301,32),
    to_unsigned(2084122954,32),
    to_unsigned(2084172588,32),
    to_unsigned(2084222203,32),
    to_unsigned(2084271799,32),
    to_unsigned(2084321375,32),
    to_unsigned(2084370933,32),
    to_unsigned(2084420471,32),
    to_unsigned(2084469990,32),
    to_unsigned(2084519489,32),
    to_unsigned(2084568970,32),
    to_unsigned(2084618432,32),
    to_unsigned(2084667874,32),
    to_unsigned(2084717297,32),
    to_unsigned(2084766701,32),
    to_unsigned(2084816086,32),
    to_unsigned(2084865452,32),
    to_unsigned(2084914798,32),
    to_unsigned(2084964126,32),
    to_unsigned(2085013434,32),
    to_unsigned(2085062723,32),
    to_unsigned(2085111993,32),
    to_unsigned(2085161243,32),
    to_unsigned(2085210475,32),
    to_unsigned(2085259687,32),
    to_unsigned(2085308881,32),
    to_unsigned(2085358055,32),
    to_unsigned(2085407209,32),
    to_unsigned(2085456345,32),
    to_unsigned(2085505462,32),
    to_unsigned(2085554559,32),
    to_unsigned(2085603637,32),
    to_unsigned(2085652696,32),
    to_unsigned(2085701736,32),
    to_unsigned(2085750757,32),
    to_unsigned(2085799758,32),
    to_unsigned(2085848741,32),
    to_unsigned(2085897704,32),
    to_unsigned(2085946648,32),
    to_unsigned(2085995573,32),
    to_unsigned(2086044478,32),
    to_unsigned(2086093365,32),
    to_unsigned(2086142232,32),
    to_unsigned(2086191080,32),
    to_unsigned(2086239909,32),
    to_unsigned(2086288719,32),
    to_unsigned(2086337509,32),
    to_unsigned(2086386281,32),
    to_unsigned(2086435033,32),
    to_unsigned(2086483766,32),
    to_unsigned(2086532480,32),
    to_unsigned(2086581175,32),
    to_unsigned(2086629850,32),
    to_unsigned(2086678507,32),
    to_unsigned(2086727144,32),
    to_unsigned(2086775762,32),
    to_unsigned(2086824361,32),
    to_unsigned(2086872940,32),
    to_unsigned(2086921501,32),
    to_unsigned(2086970042,32),
    to_unsigned(2087018564,32),
    to_unsigned(2087067067,32),
    to_unsigned(2087115551,32),
    to_unsigned(2087164015,32),
    to_unsigned(2087212460,32),
    to_unsigned(2087260887,32),
    to_unsigned(2087309293,32),
    to_unsigned(2087357681,32),
    to_unsigned(2087406050,32),
    to_unsigned(2087454399,32),
    to_unsigned(2087502729,32),
    to_unsigned(2087551040,32),
    to_unsigned(2087599332,32),
    to_unsigned(2087647605,32),
    to_unsigned(2087695858,32),
    to_unsigned(2087744093,32),
    to_unsigned(2087792308,32),
    to_unsigned(2087840504,32),
    to_unsigned(2087888680,32),
    to_unsigned(2087936838,32),
    to_unsigned(2087984976,32),
    to_unsigned(2088033095,32),
    to_unsigned(2088081195,32),
    to_unsigned(2088129276,32),
    to_unsigned(2088177338,32),
    to_unsigned(2088225380,32),
    to_unsigned(2088273403,32),
    to_unsigned(2088321407,32),
    to_unsigned(2088369392,32),
    to_unsigned(2088417357,32),
    to_unsigned(2088465304,32),
    to_unsigned(2088513231,32),
    to_unsigned(2088561139,32),
    to_unsigned(2088609028,32),
    to_unsigned(2088656897,32),
    to_unsigned(2088704748,32),
    to_unsigned(2088752579,32),
    to_unsigned(2088800391,32),
    to_unsigned(2088848184,32),
    to_unsigned(2088895957,32),
    to_unsigned(2088943712,32),
    to_unsigned(2088991447,32),
    to_unsigned(2089039163,32),
    to_unsigned(2089086859,32),
    to_unsigned(2089134537,32),
    to_unsigned(2089182195,32),
    to_unsigned(2089229835,32),
    to_unsigned(2089277455,32),
    to_unsigned(2089325055,32),
    to_unsigned(2089372637,32),
    to_unsigned(2089420199,32),
    to_unsigned(2089467742,32),
    to_unsigned(2089515266,32),
    to_unsigned(2089562771,32),
    to_unsigned(2089610257,32),
    to_unsigned(2089657723,32),
    to_unsigned(2089705170,32),
    to_unsigned(2089752598,32),
    to_unsigned(2089800007,32),
    to_unsigned(2089847396,32),
    to_unsigned(2089894766,32),
    to_unsigned(2089942117,32),
    to_unsigned(2089989449,32),
    to_unsigned(2090036762,32),
    to_unsigned(2090084055,32),
    to_unsigned(2090131330,32),
    to_unsigned(2090178585,32),
    to_unsigned(2090225820,32),
    to_unsigned(2090273037,32),
    to_unsigned(2090320234,32),
    to_unsigned(2090367413,32),
    to_unsigned(2090414572,32),
    to_unsigned(2090461711,32),
    to_unsigned(2090508832,32),
    to_unsigned(2090555933,32),
    to_unsigned(2090603015,32),
    to_unsigned(2090650078,32),
    to_unsigned(2090697122,32),
    to_unsigned(2090744146,32),
    to_unsigned(2090791151,32),
    to_unsigned(2090838137,32),
    to_unsigned(2090885104,32),
    to_unsigned(2090932052,32),
    to_unsigned(2090978980,32),
    to_unsigned(2091025889,32),
    to_unsigned(2091072779,32),
    to_unsigned(2091119650,32),
    to_unsigned(2091166501,32),
    to_unsigned(2091213333,32),
    to_unsigned(2091260146,32),
    to_unsigned(2091306940,32),
    to_unsigned(2091353715,32),
    to_unsigned(2091400470,32),
    to_unsigned(2091447206,32),
    to_unsigned(2091493923,32),
    to_unsigned(2091540621,32),
    to_unsigned(2091587299,32),
    to_unsigned(2091633959,32),
    to_unsigned(2091680599,32),
    to_unsigned(2091727219,32),
    to_unsigned(2091773821,32),
    to_unsigned(2091820403,32),
    to_unsigned(2091866966,32),
    to_unsigned(2091913510,32),
    to_unsigned(2091960035,32),
    to_unsigned(2092006540,32),
    to_unsigned(2092053026,32),
    to_unsigned(2092099493,32),
    to_unsigned(2092145941,32),
    to_unsigned(2092192370,32),
    to_unsigned(2092238779,32),
    to_unsigned(2092285169,32),
    to_unsigned(2092331540,32),
    to_unsigned(2092377891,32),
    to_unsigned(2092424223,32),
    to_unsigned(2092470537,32),
    to_unsigned(2092516830,32),
    to_unsigned(2092563105,32),
    to_unsigned(2092609360,32),
    to_unsigned(2092655597,32),
    to_unsigned(2092701814,32),
    to_unsigned(2092748011,32),
    to_unsigned(2092794190,32),
    to_unsigned(2092840349,32),
    to_unsigned(2092886489,32),
    to_unsigned(2092932610,32),
    to_unsigned(2092978711,32),
    to_unsigned(2093024793,32),
    to_unsigned(2093070856,32),
    to_unsigned(2093116900,32),
    to_unsigned(2093162925,32),
    to_unsigned(2093208930,32),
    to_unsigned(2093254916,32),
    to_unsigned(2093300883,32),
    to_unsigned(2093346831,32),
    to_unsigned(2093392759,32),
    to_unsigned(2093438668,32),
    to_unsigned(2093484558,32),
    to_unsigned(2093530428,32),
    to_unsigned(2093576280,32),
    to_unsigned(2093622112,32),
    to_unsigned(2093667925,32),
    to_unsigned(2093713718,32),
    to_unsigned(2093759493,32),
    to_unsigned(2093805248,32),
    to_unsigned(2093850984,32),
    to_unsigned(2093896701,32),
    to_unsigned(2093942398,32),
    to_unsigned(2093988076,32),
    to_unsigned(2094033735,32),
    to_unsigned(2094079375,32),
    to_unsigned(2094124995,32),
    to_unsigned(2094170596,32),
    to_unsigned(2094216178,32),
    to_unsigned(2094261741,32),
    to_unsigned(2094307284,32),
    to_unsigned(2094352809,32),
    to_unsigned(2094398313,32),
    to_unsigned(2094443799,32),
    to_unsigned(2094489266,32),
    to_unsigned(2094534713,32),
    to_unsigned(2094580141,32),
    to_unsigned(2094625549,32),
    to_unsigned(2094670939,32),
    to_unsigned(2094716309,32),
    to_unsigned(2094761660,32),
    to_unsigned(2094806991,32),
    to_unsigned(2094852304,32),
    to_unsigned(2094897597,32),
    to_unsigned(2094942871,32),
    to_unsigned(2094988125,32),
    to_unsigned(2095033361,32),
    to_unsigned(2095078577,32),
    to_unsigned(2095123774,32),
    to_unsigned(2095168951,32),
    to_unsigned(2095214110,32),
    to_unsigned(2095259249,32),
    to_unsigned(2095304369,32),
    to_unsigned(2095349469,32),
    to_unsigned(2095394550,32),
    to_unsigned(2095439612,32),
    to_unsigned(2095484655,32),
    to_unsigned(2095529679,32),
    to_unsigned(2095574683,32),
    to_unsigned(2095619668,32),
    to_unsigned(2095664634,32),
    to_unsigned(2095709580,32),
    to_unsigned(2095754507,32),
    to_unsigned(2095799415,32),
    to_unsigned(2095844304,32),
    to_unsigned(2095889173,32),
    to_unsigned(2095934024,32),
    to_unsigned(2095978854,32),
    to_unsigned(2096023666,32),
    to_unsigned(2096068458,32),
    to_unsigned(2096113232,32),
    to_unsigned(2096157985,32),
    to_unsigned(2096202720,32),
    to_unsigned(2096247435,32),
    to_unsigned(2096292131,32),
    to_unsigned(2096336808,32),
    to_unsigned(2096381465,32),
    to_unsigned(2096426104,32),
    to_unsigned(2096470723,32),
    to_unsigned(2096515322,32),
    to_unsigned(2096559903,32),
    to_unsigned(2096604464,32),
    to_unsigned(2096649006,32),
    to_unsigned(2096693528,32),
    to_unsigned(2096738031,32),
    to_unsigned(2096782515,32),
    to_unsigned(2096826980,32),
    to_unsigned(2096871426,32),
    to_unsigned(2096915852,32),
    to_unsigned(2096960259,32),
    to_unsigned(2097004647,32),
    to_unsigned(2097049015,32),
    to_unsigned(2097093364,32),
    to_unsigned(2097137694,32),
    to_unsigned(2097182004,32),
    to_unsigned(2097226296,32),
    to_unsigned(2097270568,32),
    to_unsigned(2097314820,32),
    to_unsigned(2097359054,32),
    to_unsigned(2097403268,32),
    to_unsigned(2097447463,32),
    to_unsigned(2097491639,32),
    to_unsigned(2097535795,32),
    to_unsigned(2097579932,32),
    to_unsigned(2097624050,32),
    to_unsigned(2097668148,32),
    to_unsigned(2097712227,32),
    to_unsigned(2097756287,32),
    to_unsigned(2097800328,32),
    to_unsigned(2097844349,32),
    to_unsigned(2097888351,32),
    to_unsigned(2097932334,32),
    to_unsigned(2097976298,32),
    to_unsigned(2098020242,32),
    to_unsigned(2098064167,32),
    to_unsigned(2098108073,32),
    to_unsigned(2098151959,32),
    to_unsigned(2098195826,32),
    to_unsigned(2098239674,32),
    to_unsigned(2098283502,32),
    to_unsigned(2098327312,32),
    to_unsigned(2098371102,32),
    to_unsigned(2098414872,32),
    to_unsigned(2098458624,32),
    to_unsigned(2098502356,32),
    to_unsigned(2098546068,32),
    to_unsigned(2098589762,32),
    to_unsigned(2098633436,32),
    to_unsigned(2098677091,32),
    to_unsigned(2098720727,32),
    to_unsigned(2098764343,32),
    to_unsigned(2098807940,32),
    to_unsigned(2098851518,32),
    to_unsigned(2098895076,32),
    to_unsigned(2098938616,32),
    to_unsigned(2098982135,32),
    to_unsigned(2099025636,32),
    to_unsigned(2099069117,32),
    to_unsigned(2099112579,32),
    to_unsigned(2099156022,32),
    to_unsigned(2099199445,32),
    to_unsigned(2099242849,32),
    to_unsigned(2099286234,32),
    to_unsigned(2099329600,32),
    to_unsigned(2099372946,32),
    to_unsigned(2099416273,32),
    to_unsigned(2099459581,32),
    to_unsigned(2099502869,32),
    to_unsigned(2099546138,32),
    to_unsigned(2099589388,32),
    to_unsigned(2099632618,32),
    to_unsigned(2099675829,32),
    to_unsigned(2099719021,32),
    to_unsigned(2099762194,32),
    to_unsigned(2099805347,32),
    to_unsigned(2099848481,32),
    to_unsigned(2099891595,32),
    to_unsigned(2099934691,32),
    to_unsigned(2099977767,32),
    to_unsigned(2100020824,32),
    to_unsigned(2100063861,32),
    to_unsigned(2100106879,32),
    to_unsigned(2100149878,32),
    to_unsigned(2100192857,32),
    to_unsigned(2100235818,32),
    to_unsigned(2100278759,32),
    to_unsigned(2100321680,32),
    to_unsigned(2100364582,32),
    to_unsigned(2100407465,32),
    to_unsigned(2100450329,32),
    to_unsigned(2100493173,32),
    to_unsigned(2100535999,32),
    to_unsigned(2100578804,32),
    to_unsigned(2100621591,32),
    to_unsigned(2100664358,32),
    to_unsigned(2100707106,32),
    to_unsigned(2100749834,32),
    to_unsigned(2100792543,32),
    to_unsigned(2100835233,32),
    to_unsigned(2100877904,32),
    to_unsigned(2100920555,32),
    to_unsigned(2100963187,32),
    to_unsigned(2101005800,32),
    to_unsigned(2101048393,32),
    to_unsigned(2101090967,32),
    to_unsigned(2101133522,32),
    to_unsigned(2101176057,32),
    to_unsigned(2101218573,32),
    to_unsigned(2101261070,32),
    to_unsigned(2101303548,32),
    to_unsigned(2101346006,32),
    to_unsigned(2101388445,32),
    to_unsigned(2101430864,32),
    to_unsigned(2101473264,32),
    to_unsigned(2101515645,32),
    to_unsigned(2101558007,32),
    to_unsigned(2101600349,32),
    to_unsigned(2101642672,32),
    to_unsigned(2101684976,32),
    to_unsigned(2101727260,32),
    to_unsigned(2101769525,32),
    to_unsigned(2101811771,32),
    to_unsigned(2101853997,32),
    to_unsigned(2101896204,32),
    to_unsigned(2101938392,32),
    to_unsigned(2101980560,32),
    to_unsigned(2102022709,32),
    to_unsigned(2102064839,32),
    to_unsigned(2102106949,32),
    to_unsigned(2102149040,32),
    to_unsigned(2102191112,32),
    to_unsigned(2102233165,32),
    to_unsigned(2102275198,32),
    to_unsigned(2102317212,32),
    to_unsigned(2102359206,32),
    to_unsigned(2102401181,32),
    to_unsigned(2102443137,32),
    to_unsigned(2102485074,32),
    to_unsigned(2102526991,32),
    to_unsigned(2102568889,32),
    to_unsigned(2102610767,32),
    to_unsigned(2102652626,32),
    to_unsigned(2102694466,32),
    to_unsigned(2102736287,32),
    to_unsigned(2102778088,32),
    to_unsigned(2102819870,32),
    to_unsigned(2102861632,32),
    to_unsigned(2102903376,32),
    to_unsigned(2102945100,32),
    to_unsigned(2102986804,32),
    to_unsigned(2103028489,32),
    to_unsigned(2103070155,32),
    to_unsigned(2103111802,32),
    to_unsigned(2103153429,32),
    to_unsigned(2103195037,32),
    to_unsigned(2103236626,32),
    to_unsigned(2103278195,32),
    to_unsigned(2103319745,32),
    to_unsigned(2103361275,32),
    to_unsigned(2103402787,32),
    to_unsigned(2103444279,32),
    to_unsigned(2103485751,32),
    to_unsigned(2103527204,32),
    to_unsigned(2103568638,32),
    to_unsigned(2103610053,32),
    to_unsigned(2103651448,32),
    to_unsigned(2103692824,32),
    to_unsigned(2103734181,32),
    to_unsigned(2103775518,32),
    to_unsigned(2103816836,32),
    to_unsigned(2103858134,32),
    to_unsigned(2103899414,32),
    to_unsigned(2103940673,32),
    to_unsigned(2103981914,32),
    to_unsigned(2104023135,32),
    to_unsigned(2104064337,32),
    to_unsigned(2104105520,32),
    to_unsigned(2104146683,32),
    to_unsigned(2104187827,32),
    to_unsigned(2104228951,32),
    to_unsigned(2104270056,32),
    to_unsigned(2104311142,32),
    to_unsigned(2104352209,32),
    to_unsigned(2104393256,32),
    to_unsigned(2104434283,32),
    to_unsigned(2104475292,32),
    to_unsigned(2104516281,32),
    to_unsigned(2104557251,32),
    to_unsigned(2104598201,32),
    to_unsigned(2104639132,32),
    to_unsigned(2104680044,32),
    to_unsigned(2104720936,32),
    to_unsigned(2104761809,32),
    to_unsigned(2104802663,32),
    to_unsigned(2104843497,32),
    to_unsigned(2104884312,32),
    to_unsigned(2104925108,32),
    to_unsigned(2104965884,32),
    to_unsigned(2105006641,32),
    to_unsigned(2105047379,32),
    to_unsigned(2105088097,32),
    to_unsigned(2105128796,32),
    to_unsigned(2105169476,32),
    to_unsigned(2105210136,32),
    to_unsigned(2105250777,32),
    to_unsigned(2105291398,32),
    to_unsigned(2105332000,32),
    to_unsigned(2105372583,32),
    to_unsigned(2105413147,32),
    to_unsigned(2105453691,32),
    to_unsigned(2105494215,32),
    to_unsigned(2105534721,32),
    to_unsigned(2105575207,32),
    to_unsigned(2105615673,32),
    to_unsigned(2105656121,32),
    to_unsigned(2105696549,32),
    to_unsigned(2105736957,32),
    to_unsigned(2105777347,32),
    to_unsigned(2105817717,32),
    to_unsigned(2105858067,32),
    to_unsigned(2105898398,32),
    to_unsigned(2105938710,32),
    to_unsigned(2105979003,32),
    to_unsigned(2106019276,32),
    to_unsigned(2106059529,32),
    to_unsigned(2106099764,32),
    to_unsigned(2106139979,32),
    to_unsigned(2106180175,32),
    to_unsigned(2106220351,32),
    to_unsigned(2106260508,32),
    to_unsigned(2106300645,32),
    to_unsigned(2106340764,32),
    to_unsigned(2106380863,32),
    to_unsigned(2106420942,32),
    to_unsigned(2106461002,32),
    to_unsigned(2106501043,32),
    to_unsigned(2106541064,32),
    to_unsigned(2106581067,32),
    to_unsigned(2106621049,32),
    to_unsigned(2106661013,32),
    to_unsigned(2106700957,32),
    to_unsigned(2106740881,32),
    to_unsigned(2106780786,32),
    to_unsigned(2106820672,32),
    to_unsigned(2106860539,32),
    to_unsigned(2106900386,32),
    to_unsigned(2106940214,32),
    to_unsigned(2106980022,32),
    to_unsigned(2107019811,32),
    to_unsigned(2107059581,32),
    to_unsigned(2107099331,32),
    to_unsigned(2107139062,32),
    to_unsigned(2107178774,32),
    to_unsigned(2107218466,32),
    to_unsigned(2107258139,32),
    to_unsigned(2107297792,32),
    to_unsigned(2107337426,32),
    to_unsigned(2107377041,32),
    to_unsigned(2107416637,32),
    to_unsigned(2107456213,32),
    to_unsigned(2107495769,32),
    to_unsigned(2107535306,32),
    to_unsigned(2107574824,32),
    to_unsigned(2107614323,32),
    to_unsigned(2107653802,32),
    to_unsigned(2107693262,32),
    to_unsigned(2107732702,32),
    to_unsigned(2107772123,32),
    to_unsigned(2107811525,32),
    to_unsigned(2107850907,32),
    to_unsigned(2107890270,32),
    to_unsigned(2107929613,32),
    to_unsigned(2107968938,32),
    to_unsigned(2108008242,32),
    to_unsigned(2108047528,32),
    to_unsigned(2108086794,32),
    to_unsigned(2108126040,32),
    to_unsigned(2108165268,32),
    to_unsigned(2108204475,32),
    to_unsigned(2108243664,32),
    to_unsigned(2108282833,32),
    to_unsigned(2108321983,32),
    to_unsigned(2108361113,32),
    to_unsigned(2108400224,32),
    to_unsigned(2108439316,32),
    to_unsigned(2108478388,32),
    to_unsigned(2108517441,32),
    to_unsigned(2108556474,32),
    to_unsigned(2108595488,32),
    to_unsigned(2108634483,32),
    to_unsigned(2108673458,32),
    to_unsigned(2108712414,32),
    to_unsigned(2108751351,32),
    to_unsigned(2108790268,32),
    to_unsigned(2108829166,32),
    to_unsigned(2108868044,32),
    to_unsigned(2108906903,32),
    to_unsigned(2108945743,32),
    to_unsigned(2108984563,32),
    to_unsigned(2109023364,32),
    to_unsigned(2109062145,32),
    to_unsigned(2109100908,32),
    to_unsigned(2109139650,32),
    to_unsigned(2109178374,32),
    to_unsigned(2109217077,32),
    to_unsigned(2109255762,32),
    to_unsigned(2109294427,32),
    to_unsigned(2109333073,32),
    to_unsigned(2109371699,32),
    to_unsigned(2109410306,32),
    to_unsigned(2109448894,32),
    to_unsigned(2109487462,32),
    to_unsigned(2109526011,32),
    to_unsigned(2109564540,32),
    to_unsigned(2109603050,32),
    to_unsigned(2109641541,32),
    to_unsigned(2109680012,32),
    to_unsigned(2109718464,32),
    to_unsigned(2109756897,32),
    to_unsigned(2109795310,32),
    to_unsigned(2109833703,32),
    to_unsigned(2109872078,32),
    to_unsigned(2109910433,32),
    to_unsigned(2109948768,32),
    to_unsigned(2109987084,32),
    to_unsigned(2110025381,32),
    to_unsigned(2110063658,32),
    to_unsigned(2110101916,32),
    to_unsigned(2110140155,32),
    to_unsigned(2110178374,32),
    to_unsigned(2110216574,32),
    to_unsigned(2110254754,32),
    to_unsigned(2110292915,32),
    to_unsigned(2110331056,32),
    to_unsigned(2110369179,32),
    to_unsigned(2110407281,32),
    to_unsigned(2110445365,32),
    to_unsigned(2110483429,32),
    to_unsigned(2110521473,32),
    to_unsigned(2110559498,32),
    to_unsigned(2110597504,32),
    to_unsigned(2110635490,32),
    to_unsigned(2110673457,32),
    to_unsigned(2110711405,32),
    to_unsigned(2110749333,32),
    to_unsigned(2110787242,32),
    to_unsigned(2110825131,32),
    to_unsigned(2110863001,32),
    to_unsigned(2110900852,32),
    to_unsigned(2110938683,32),
    to_unsigned(2110976495,32),
    to_unsigned(2111014287,32),
    to_unsigned(2111052060,32),
    to_unsigned(2111089813,32),
    to_unsigned(2111127548,32),
    to_unsigned(2111165262,32),
    to_unsigned(2111202958,32),
    to_unsigned(2111240633,32),
    to_unsigned(2111278290,32),
    to_unsigned(2111315927,32),
    to_unsigned(2111353545,32),
    to_unsigned(2111391143,32),
    to_unsigned(2111428722,32),
    to_unsigned(2111466281,32),
    to_unsigned(2111503821,32),
    to_unsigned(2111541342,32),
    to_unsigned(2111578843,32),
    to_unsigned(2111616325,32),
    to_unsigned(2111653788,32),
    to_unsigned(2111691231,32),
    to_unsigned(2111728654,32),
    to_unsigned(2111766058,32),
    to_unsigned(2111803443,32),
    to_unsigned(2111840808,32),
    to_unsigned(2111878154,32),
    to_unsigned(2111915481,32),
    to_unsigned(2111952788,32),
    to_unsigned(2111990076,32),
    to_unsigned(2112027344,32),
    to_unsigned(2112064593,32),
    to_unsigned(2112101823,32),
    to_unsigned(2112139033,32),
    to_unsigned(2112176223,32),
    to_unsigned(2112213394,32),
    to_unsigned(2112250546,32),
    to_unsigned(2112287679,32),
    to_unsigned(2112324792,32),
    to_unsigned(2112361885,32),
    to_unsigned(2112398959,32),
    to_unsigned(2112436014,32),
    to_unsigned(2112473049,32),
    to_unsigned(2112510065,32),
    to_unsigned(2112547062,32),
    to_unsigned(2112584039,32),
    to_unsigned(2112620997,32),
    to_unsigned(2112657935,32),
    to_unsigned(2112694854,32),
    to_unsigned(2112731753,32),
    to_unsigned(2112768633,32),
    to_unsigned(2112805494,32),
    to_unsigned(2112842335,32),
    to_unsigned(2112879156,32),
    to_unsigned(2112915959,32),
    to_unsigned(2112952742,32),
    to_unsigned(2112989505,32),
    to_unsigned(2113026249,32),
    to_unsigned(2113062974,32),
    to_unsigned(2113099679,32),
    to_unsigned(2113136365,32),
    to_unsigned(2113173031,32),
    to_unsigned(2113209678,32),
    to_unsigned(2113246305,32),
    to_unsigned(2113282913,32),
    to_unsigned(2113319502,32),
    to_unsigned(2113356071,32),
    to_unsigned(2113392621,32),
    to_unsigned(2113429151,32),
    to_unsigned(2113465662,32),
    to_unsigned(2113502154,32),
    to_unsigned(2113538626,32),
    to_unsigned(2113575079,32),
    to_unsigned(2113611512,32),
    to_unsigned(2113647926,32),
    to_unsigned(2113684320,32),
    to_unsigned(2113720695,32),
    to_unsigned(2113757050,32),
    to_unsigned(2113793387,32),
    to_unsigned(2113829703,32),
    to_unsigned(2113866000,32),
    to_unsigned(2113902278,32),
    to_unsigned(2113938537,32),
    to_unsigned(2113974776,32),
    to_unsigned(2114010995,32),
    to_unsigned(2114047195,32),
    to_unsigned(2114083376,32),
    to_unsigned(2114119537,32),
    to_unsigned(2114155679,32),
    to_unsigned(2114191801,32),
    to_unsigned(2114227904,32),
    to_unsigned(2114263987,32),
    to_unsigned(2114300051,32),
    to_unsigned(2114336096,32),
    to_unsigned(2114372121,32),
    to_unsigned(2114408127,32),
    to_unsigned(2114444113,32),
    to_unsigned(2114480080,32),
    to_unsigned(2114516028,32),
    to_unsigned(2114551956,32),
    to_unsigned(2114587864,32),
    to_unsigned(2114623753,32),
    to_unsigned(2114659623,32),
    to_unsigned(2114695473,32),
    to_unsigned(2114731304,32),
    to_unsigned(2114767115,32),
    to_unsigned(2114802907,32),
    to_unsigned(2114838680,32),
    to_unsigned(2114874433,32),
    to_unsigned(2114910166,32),
    to_unsigned(2114945881,32),
    to_unsigned(2114981575,32),
    to_unsigned(2115017251,32),
    to_unsigned(2115052907,32),
    to_unsigned(2115088543,32),
    to_unsigned(2115124160,32),
    to_unsigned(2115159757,32),
    to_unsigned(2115195336,32),
    to_unsigned(2115230894,32),
    to_unsigned(2115266433,32),
    to_unsigned(2115301953,32),
    to_unsigned(2115337453,32),
    to_unsigned(2115372934,32),
    to_unsigned(2115408396,32),
    to_unsigned(2115443838,32),
    to_unsigned(2115479260,32),
    to_unsigned(2115514663,32),
    to_unsigned(2115550047,32),
    to_unsigned(2115585411,32),
    to_unsigned(2115620756,32),
    to_unsigned(2115656081,32),
    to_unsigned(2115691387,32),
    to_unsigned(2115726674,32),
    to_unsigned(2115761941,32),
    to_unsigned(2115797188,32),
    to_unsigned(2115832416,32),
    to_unsigned(2115867625,32),
    to_unsigned(2115902814,32),
    to_unsigned(2115937984,32),
    to_unsigned(2115973134,32),
    to_unsigned(2116008265,32),
    to_unsigned(2116043376,32),
    to_unsigned(2116078468,32),
    to_unsigned(2116113541,32),
    to_unsigned(2116148594,32),
    to_unsigned(2116183627,32),
    to_unsigned(2116218641,32),
    to_unsigned(2116253636,32),
    to_unsigned(2116288611,32),
    to_unsigned(2116323567,32),
    to_unsigned(2116358503,32),
    to_unsigned(2116393420,32),
    to_unsigned(2116428318,32),
    to_unsigned(2116463196,32),
    to_unsigned(2116498054,32),
    to_unsigned(2116532893,32),
    to_unsigned(2116567713,32),
    to_unsigned(2116602513,32),
    to_unsigned(2116637293,32),
    to_unsigned(2116672055,32),
    to_unsigned(2116706796,32),
    to_unsigned(2116741519,32),
    to_unsigned(2116776222,32),
    to_unsigned(2116810905,32),
    to_unsigned(2116845569,32),
    to_unsigned(2116880213,32),
    to_unsigned(2116914839,32),
    to_unsigned(2116949444,32),
    to_unsigned(2116984030,32),
    to_unsigned(2117018597,32),
    to_unsigned(2117053144,32),
    to_unsigned(2117087672,32),
    to_unsigned(2117122180,32),
    to_unsigned(2117156669,32),
    to_unsigned(2117191138,32),
    to_unsigned(2117225588,32),
    to_unsigned(2117260019,32),
    to_unsigned(2117294430,32),
    to_unsigned(2117328821,32),
    to_unsigned(2117363193,32),
    to_unsigned(2117397546,32),
    to_unsigned(2117431879,32),
    to_unsigned(2117466192,32),
    to_unsigned(2117500487,32),
    to_unsigned(2117534761,32),
    to_unsigned(2117569017,32),
    to_unsigned(2117603252,32),
    to_unsigned(2117637469,32),
    to_unsigned(2117671666,32),
    to_unsigned(2117705843,32),
    to_unsigned(2117740001,32),
    to_unsigned(2117774139,32),
    to_unsigned(2117808258,32),
    to_unsigned(2117842358,32),
    to_unsigned(2117876438,32),
    to_unsigned(2117910499,32),
    to_unsigned(2117944540,32),
    to_unsigned(2117978562,32),
    to_unsigned(2118012564,32),
    to_unsigned(2118046546,32),
    to_unsigned(2118080510,32),
    to_unsigned(2118114454,32),
    to_unsigned(2118148378,32),
    to_unsigned(2118182283,32),
    to_unsigned(2118216168,32),
    to_unsigned(2118250034,32),
    to_unsigned(2118283881,32),
    to_unsigned(2118317707,32),
    to_unsigned(2118351515,32),
    to_unsigned(2118385303,32),
    to_unsigned(2118419072,32),
    to_unsigned(2118452821,32),
    to_unsigned(2118486550,32),
    to_unsigned(2118520260,32),
    to_unsigned(2118553951,32),
    to_unsigned(2118587622,32),
    to_unsigned(2118621274,32),
    to_unsigned(2118654906,32),
    to_unsigned(2118688519,32),
    to_unsigned(2118722112,32),
    to_unsigned(2118755686,32),
    to_unsigned(2118789241,32),
    to_unsigned(2118822775,32),
    to_unsigned(2118856291,32),
    to_unsigned(2118889787,32),
    to_unsigned(2118923263,32),
    to_unsigned(2118956720,32),
    to_unsigned(2118990158,32),
    to_unsigned(2119023576,32),
    to_unsigned(2119056974,32),
    to_unsigned(2119090353,32),
    to_unsigned(2119123713,32),
    to_unsigned(2119157053,32),
    to_unsigned(2119190374,32),
    to_unsigned(2119223675,32),
    to_unsigned(2119256957,32),
    to_unsigned(2119290219,32),
    to_unsigned(2119323461,32),
    to_unsigned(2119356685,32),
    to_unsigned(2119389888,32),
    to_unsigned(2119423073,32),
    to_unsigned(2119456238,32),
    to_unsigned(2119489383,32),
    to_unsigned(2119522509,32),
    to_unsigned(2119555615,32),
    to_unsigned(2119588702,32),
    to_unsigned(2119621769,32),
    to_unsigned(2119654817,32),
    to_unsigned(2119687846,32),
    to_unsigned(2119720854,32),
    to_unsigned(2119753844,32),
    to_unsigned(2119786814,32),
    to_unsigned(2119819764,32),
    to_unsigned(2119852695,32),
    to_unsigned(2119885607,32),
    to_unsigned(2119918499,32),
    to_unsigned(2119951371,32),
    to_unsigned(2119984224,32),
    to_unsigned(2120017058,32),
    to_unsigned(2120049872,32),
    to_unsigned(2120082667,32),
    to_unsigned(2120115442,32),
    to_unsigned(2120148197,32),
    to_unsigned(2120180934,32),
    to_unsigned(2120213650,32),
    to_unsigned(2120246347,32),
    to_unsigned(2120279025,32),
    to_unsigned(2120311683,32),
    to_unsigned(2120344322,32),
    to_unsigned(2120376941,32),
    to_unsigned(2120409541,32),
    to_unsigned(2120442121,32),
    to_unsigned(2120474682,32),
    to_unsigned(2120507223,32),
    to_unsigned(2120539745,32),
    to_unsigned(2120572247,32),
    to_unsigned(2120604730,32),
    to_unsigned(2120637193,32),
    to_unsigned(2120669637,32),
    to_unsigned(2120702061,32),
    to_unsigned(2120734466,32),
    to_unsigned(2120766851,32),
    to_unsigned(2120799217,32),
    to_unsigned(2120831563,32),
    to_unsigned(2120863890,32),
    to_unsigned(2120896197,32),
    to_unsigned(2120928485,32),
    to_unsigned(2120960753,32),
    to_unsigned(2120993002,32),
    to_unsigned(2121025232,32),
    to_unsigned(2121057441,32),
    to_unsigned(2121089632,32),
    to_unsigned(2121121803,32),
    to_unsigned(2121153954,32),
    to_unsigned(2121186086,32),
    to_unsigned(2121218198,32),
    to_unsigned(2121250291,32),
    to_unsigned(2121282364,32),
    to_unsigned(2121314418,32),
    to_unsigned(2121346453,32),
    to_unsigned(2121378467,32),
    to_unsigned(2121410463,32),
    to_unsigned(2121442439,32),
    to_unsigned(2121474395,32),
    to_unsigned(2121506332,32),
    to_unsigned(2121538249,32),
    to_unsigned(2121570147,32),
    to_unsigned(2121602025,32),
    to_unsigned(2121633884,32),
    to_unsigned(2121665724,32),
    to_unsigned(2121697543,32),
    to_unsigned(2121729344,32),
    to_unsigned(2121761125,32),
    to_unsigned(2121792886,32),
    to_unsigned(2121824628,32),
    to_unsigned(2121856350,32),
    to_unsigned(2121888053,32),
    to_unsigned(2121919736,32),
    to_unsigned(2121951400,32),
    to_unsigned(2121983045,32),
    to_unsigned(2122014669,32),
    to_unsigned(2122046275,32),
    to_unsigned(2122077860,32),
    to_unsigned(2122109427,32),
    to_unsigned(2122140974,32),
    to_unsigned(2122172501,32),
    to_unsigned(2122204009,32),
    to_unsigned(2122235497,32),
    to_unsigned(2122266966,32),
    to_unsigned(2122298415,32),
    to_unsigned(2122329845,32),
    to_unsigned(2122361255,32),
    to_unsigned(2122392646,32),
    to_unsigned(2122424017,32),
    to_unsigned(2122455369,32),
    to_unsigned(2122486701,32),
    to_unsigned(2122518014,32),
    to_unsigned(2122549307,32),
    to_unsigned(2122580580,32),
    to_unsigned(2122611835,32),
    to_unsigned(2122643069,32),
    to_unsigned(2122674284,32),
    to_unsigned(2122705480,32),
    to_unsigned(2122736656,32),
    to_unsigned(2122767813,32),
    to_unsigned(2122798950,32),
    to_unsigned(2122830068,32),
    to_unsigned(2122861166,32),
    to_unsigned(2122892244,32),
    to_unsigned(2122923303,32),
    to_unsigned(2122954343,32),
    to_unsigned(2122985363,32),
    to_unsigned(2123016363,32),
    to_unsigned(2123047344,32),
    to_unsigned(2123078306,32),
    to_unsigned(2123109248,32),
    to_unsigned(2123140170,32),
    to_unsigned(2123171073,32),
    to_unsigned(2123201957,32),
    to_unsigned(2123232821,32),
    to_unsigned(2123263665,32),
    to_unsigned(2123294490,32),
    to_unsigned(2123325295,32),
    to_unsigned(2123356081,32),
    to_unsigned(2123386847,32),
    to_unsigned(2123417594,32),
    to_unsigned(2123448321,32),
    to_unsigned(2123479029,32),
    to_unsigned(2123509717,32),
    to_unsigned(2123540386,32),
    to_unsigned(2123571035,32),
    to_unsigned(2123601665,32),
    to_unsigned(2123632275,32),
    to_unsigned(2123662866,32),
    to_unsigned(2123693437,32),
    to_unsigned(2123723989,32),
    to_unsigned(2123754521,32),
    to_unsigned(2123785033,32),
    to_unsigned(2123815526,32),
    to_unsigned(2123846000,32),
    to_unsigned(2123876454,32),
    to_unsigned(2123906888,32),
    to_unsigned(2123937303,32),
    to_unsigned(2123967699,32),
    to_unsigned(2123998075,32),
    to_unsigned(2124028431,32),
    to_unsigned(2124058768,32),
    to_unsigned(2124089085,32),
    to_unsigned(2124119383,32),
    to_unsigned(2124149661,32),
    to_unsigned(2124179920,32),
    to_unsigned(2124210159,32),
    to_unsigned(2124240379,32),
    to_unsigned(2124270579,32),
    to_unsigned(2124300760,32),
    to_unsigned(2124330921,32),
    to_unsigned(2124361063,32),
    to_unsigned(2124391185,32),
    to_unsigned(2124421287,32),
    to_unsigned(2124451370,32),
    to_unsigned(2124481434,32),
    to_unsigned(2124511478,32),
    to_unsigned(2124541502,32),
    to_unsigned(2124571507,32),
    to_unsigned(2124601493,32),
    to_unsigned(2124631459,32),
    to_unsigned(2124661405,32),
    to_unsigned(2124691332,32),
    to_unsigned(2124721239,32),
    to_unsigned(2124751127,32),
    to_unsigned(2124780995,32),
    to_unsigned(2124810844,32),
    to_unsigned(2124840673,32),
    to_unsigned(2124870482,32),
    to_unsigned(2124900273,32),
    to_unsigned(2124930043,32),
    to_unsigned(2124959794,32),
    to_unsigned(2124989526,32),
    to_unsigned(2125019238,32),
    to_unsigned(2125048930,32),
    to_unsigned(2125078603,32),
    to_unsigned(2125108256,32),
    to_unsigned(2125137890,32),
    to_unsigned(2125167504,32),
    to_unsigned(2125197099,32),
    to_unsigned(2125226674,32),
    to_unsigned(2125256230,32),
    to_unsigned(2125285766,32),
    to_unsigned(2125315283,32),
    to_unsigned(2125344780,32),
    to_unsigned(2125374258,32),
    to_unsigned(2125403716,32),
    to_unsigned(2125433154,32),
    to_unsigned(2125462573,32),
    to_unsigned(2125491972,32),
    to_unsigned(2125521352,32),
    to_unsigned(2125550713,32),
    to_unsigned(2125580053,32),
    to_unsigned(2125609375,32),
    to_unsigned(2125638676,32),
    to_unsigned(2125667959,32),
    to_unsigned(2125697221,32),
    to_unsigned(2125726464,32),
    to_unsigned(2125755688,32),
    to_unsigned(2125784892,32),
    to_unsigned(2125814076,32),
    to_unsigned(2125843241,32),
    to_unsigned(2125872387,32),
    to_unsigned(2125901513,32),
    to_unsigned(2125930619,32),
    to_unsigned(2125959706,32),
    to_unsigned(2125988773,32),
    to_unsigned(2126017821,32),
    to_unsigned(2126046849,32),
    to_unsigned(2126075858,32),
    to_unsigned(2126104847,32),
    to_unsigned(2126133816,32),
    to_unsigned(2126162766,32),
    to_unsigned(2126191697,32),
    to_unsigned(2126220607,32),
    to_unsigned(2126249499,32),
    to_unsigned(2126278371,32),
    to_unsigned(2126307223,32),
    to_unsigned(2126336056,32),
    to_unsigned(2126364869,32),
    to_unsigned(2126393662,32),
    to_unsigned(2126422437,32),
    to_unsigned(2126451191,32),
    to_unsigned(2126479926,32),
    to_unsigned(2126508642,32),
    to_unsigned(2126537337,32),
    to_unsigned(2126566014,32),
    to_unsigned(2126594671,32),
    to_unsigned(2126623308,32),
    to_unsigned(2126651926,32),
    to_unsigned(2126680524,32),
    to_unsigned(2126709102,32),
    to_unsigned(2126737661,32),
    to_unsigned(2126766201,32),
    to_unsigned(2126794721,32),
    to_unsigned(2126823221,32),
    to_unsigned(2126851702,32),
    to_unsigned(2126880164,32),
    to_unsigned(2126908605,32),
    to_unsigned(2126937028,32),
    to_unsigned(2126965430,32),
    to_unsigned(2126993813,32),
    to_unsigned(2127022177,32),
    to_unsigned(2127050521,32),
    to_unsigned(2127078846,32),
    to_unsigned(2127107150,32),
    to_unsigned(2127135436,32),
    to_unsigned(2127163702,32),
    to_unsigned(2127191948,32),
    to_unsigned(2127220175,32),
    to_unsigned(2127248382,32),
    to_unsigned(2127276569,32),
    to_unsigned(2127304737,32),
    to_unsigned(2127332886,32),
    to_unsigned(2127361015,32),
    to_unsigned(2127389124,32),
    to_unsigned(2127417214,32),
    to_unsigned(2127445284,32),
    to_unsigned(2127473335,32),
    to_unsigned(2127501366,32),
    to_unsigned(2127529378,32),
    to_unsigned(2127557370,32),
    to_unsigned(2127585342,32),
    to_unsigned(2127613295,32),
    to_unsigned(2127641229,32),
    to_unsigned(2127669143,32),
    to_unsigned(2127697037,32),
    to_unsigned(2127724912,32),
    to_unsigned(2127752767,32),
    to_unsigned(2127780602,32),
    to_unsigned(2127808418,32),
    to_unsigned(2127836215,32),
    to_unsigned(2127863992,32),
    to_unsigned(2127891749,32),
    to_unsigned(2127919487,32),
    to_unsigned(2127947205,32),
    to_unsigned(2127974904,32),
    to_unsigned(2128002583,32),
    to_unsigned(2128030243,32),
    to_unsigned(2128057883,32),
    to_unsigned(2128085503,32),
    to_unsigned(2128113104,32),
    to_unsigned(2128140685,32),
    to_unsigned(2128168247,32),
    to_unsigned(2128195789,32),
    to_unsigned(2128223312,32),
    to_unsigned(2128250815,32),
    to_unsigned(2128278299,32),
    to_unsigned(2128305763,32),
    to_unsigned(2128333207,32),
    to_unsigned(2128360632,32),
    to_unsigned(2128388037,32),
    to_unsigned(2128415423,32),
    to_unsigned(2128442789,32),
    to_unsigned(2128470136,32),
    to_unsigned(2128497463,32),
    to_unsigned(2128524770,32),
    to_unsigned(2128552058,32),
    to_unsigned(2128579326,32),
    to_unsigned(2128606575,32),
    to_unsigned(2128633804,32),
    to_unsigned(2128661014,32),
    to_unsigned(2128688204,32),
    to_unsigned(2128715374,32),
    to_unsigned(2128742525,32),
    to_unsigned(2128769657,32),
    to_unsigned(2128796768,32),
    to_unsigned(2128823861,32),
    to_unsigned(2128850933,32),
    to_unsigned(2128877986,32),
    to_unsigned(2128905020,32),
    to_unsigned(2128932034,32),
    to_unsigned(2128959028,32),
    to_unsigned(2128986003,32),
    to_unsigned(2129012958,32),
    to_unsigned(2129039894,32),
    to_unsigned(2129066810,32),
    to_unsigned(2129093707,32),
    to_unsigned(2129120584,32),
    to_unsigned(2129147441,32),
    to_unsigned(2129174279,32),
    to_unsigned(2129201097,32),
    to_unsigned(2129227896,32),
    to_unsigned(2129254675,32),
    to_unsigned(2129281434,32),
    to_unsigned(2129308174,32),
    to_unsigned(2129334895,32),
    to_unsigned(2129361595,32),
    to_unsigned(2129388277,32),
    to_unsigned(2129414938,32),
    to_unsigned(2129441580,32),
    to_unsigned(2129468203,32),
    to_unsigned(2129494806,32),
    to_unsigned(2129521389,32),
    to_unsigned(2129547953,32),
    to_unsigned(2129574497,32),
    to_unsigned(2129601022,32),
    to_unsigned(2129627527,32),
    to_unsigned(2129654013,32),
    to_unsigned(2129680479,32),
    to_unsigned(2129706925,32),
    to_unsigned(2129733352,32),
    to_unsigned(2129759759,32),
    to_unsigned(2129786147,32),
    to_unsigned(2129812515,32),
    to_unsigned(2129838863,32),
    to_unsigned(2129865192,32),
    to_unsigned(2129891501,32),
    to_unsigned(2129917791,32),
    to_unsigned(2129944061,32),
    to_unsigned(2129970312,32),
    to_unsigned(2129996543,32),
    to_unsigned(2130022754,32),
    to_unsigned(2130048946,32),
    to_unsigned(2130075118,32),
    to_unsigned(2130101271,32),
    to_unsigned(2130127404,32),
    to_unsigned(2130153518,32),
    to_unsigned(2130179612,32),
    to_unsigned(2130205686,32),
    to_unsigned(2130231741,32),
    to_unsigned(2130257776,32),
    to_unsigned(2130283792,32),
    to_unsigned(2130309788,32),
    to_unsigned(2130335764,32),
    to_unsigned(2130361721,32),
    to_unsigned(2130387658,32),
    to_unsigned(2130413576,32),
    to_unsigned(2130439474,32),
    to_unsigned(2130465353,32),
    to_unsigned(2130491212,32),
    to_unsigned(2130517051,32),
    to_unsigned(2130542871,32),
    to_unsigned(2130568671,32),
    to_unsigned(2130594452,32),
    to_unsigned(2130620213,32),
    to_unsigned(2130645954,32),
    to_unsigned(2130671676,32),
    to_unsigned(2130697379,32),
    to_unsigned(2130723061,32),
    to_unsigned(2130748724,32),
    to_unsigned(2130774368,32),
    to_unsigned(2130799992,32),
    to_unsigned(2130825596,32),
    to_unsigned(2130851181,32),
    to_unsigned(2130876746,32),
    to_unsigned(2130902292,32),
    to_unsigned(2130927818,32),
    to_unsigned(2130953324,32),
    to_unsigned(2130978811,32),
    to_unsigned(2131004279,32),
    to_unsigned(2131029726,32),
    to_unsigned(2131055154,32),
    to_unsigned(2131080563,32),
    to_unsigned(2131105952,32),
    to_unsigned(2131131321,32),
    to_unsigned(2131156671,32),
    to_unsigned(2131182001,32),
    to_unsigned(2131207312,32),
    to_unsigned(2131232603,32),
    to_unsigned(2131257874,32),
    to_unsigned(2131283126,32),
    to_unsigned(2131308358,32),
    to_unsigned(2131333571,32),
    to_unsigned(2131358764,32),
    to_unsigned(2131383937,32),
    to_unsigned(2131409091,32),
    to_unsigned(2131434225,32),
    to_unsigned(2131459340,32),
    to_unsigned(2131484435,32),
    to_unsigned(2131509510,32),
    to_unsigned(2131534566,32),
    to_unsigned(2131559602,32),
    to_unsigned(2131584619,32),
    to_unsigned(2131609616,32),
    to_unsigned(2131634594,32),
    to_unsigned(2131659552,32),
    to_unsigned(2131684490,32),
    to_unsigned(2131709409,32),
    to_unsigned(2131734308,32),
    to_unsigned(2131759187,32),
    to_unsigned(2131784047,32),
    to_unsigned(2131808888,32),
    to_unsigned(2131833708,32),
    to_unsigned(2131858510,32),
    to_unsigned(2131883291,32),
    to_unsigned(2131908053,32),
    to_unsigned(2131932795,32),
    to_unsigned(2131957518,32),
    to_unsigned(2131982221,32),
    to_unsigned(2132006905,32),
    to_unsigned(2132031569,32),
    to_unsigned(2132056213,32),
    to_unsigned(2132080838,32),
    to_unsigned(2132105443,32),
    to_unsigned(2132130029,32),
    to_unsigned(2132154595,32),
    to_unsigned(2132179141,32),
    to_unsigned(2132203668,32),
    to_unsigned(2132228175,32),
    to_unsigned(2132252663,32),
    to_unsigned(2132277131,32),
    to_unsigned(2132301579,32),
    to_unsigned(2132326008,32),
    to_unsigned(2132350417,32),
    to_unsigned(2132374807,32),
    to_unsigned(2132399177,32),
    to_unsigned(2132423527,32),
    to_unsigned(2132447858,32),
    to_unsigned(2132472169,32),
    to_unsigned(2132496461,32),
    to_unsigned(2132520733,32),
    to_unsigned(2132544985,32),
    to_unsigned(2132569218,32),
    to_unsigned(2132593431,32),
    to_unsigned(2132617625,32),
    to_unsigned(2132641799,32),
    to_unsigned(2132665953,32),
    to_unsigned(2132690088,32),
    to_unsigned(2132714203,32),
    to_unsigned(2132738299,32),
    to_unsigned(2132762375,32),
    to_unsigned(2132786431,32),
    to_unsigned(2132810468,32),
    to_unsigned(2132834485,32),
    to_unsigned(2132858483,32),
    to_unsigned(2132882461,32),
    to_unsigned(2132906419,32),
    to_unsigned(2132930358,32),
    to_unsigned(2132954277,32),
    to_unsigned(2132978176,32),
    to_unsigned(2133002056,32),
    to_unsigned(2133025917,32),
    to_unsigned(2133049757,32),
    to_unsigned(2133073578,32),
    to_unsigned(2133097380,32),
    to_unsigned(2133121162,32),
    to_unsigned(2133144924,32),
    to_unsigned(2133168667,32),
    to_unsigned(2133192390,32),
    to_unsigned(2133216093,32),
    to_unsigned(2133239777,32),
    to_unsigned(2133263441,32),
    to_unsigned(2133287086,32),
    to_unsigned(2133310711,32),
    to_unsigned(2133334316,32),
    to_unsigned(2133357902,32),
    to_unsigned(2133381468,32),
    to_unsigned(2133405015,32),
    to_unsigned(2133428542,32),
    to_unsigned(2133452049,32),
    to_unsigned(2133475537,32),
    to_unsigned(2133499005,32),
    to_unsigned(2133522454,32),
    to_unsigned(2133545883,32),
    to_unsigned(2133569292,32),
    to_unsigned(2133592682,32),
    to_unsigned(2133616052,32),
    to_unsigned(2133639402,32),
    to_unsigned(2133662733,32),
    to_unsigned(2133686045,32),
    to_unsigned(2133709336,32),
    to_unsigned(2133732608,32),
    to_unsigned(2133755861,32),
    to_unsigned(2133779093,32),
    to_unsigned(2133802307,32),
    to_unsigned(2133825500,32),
    to_unsigned(2133848674,32),
    to_unsigned(2133871829,32),
    to_unsigned(2133894963,32),
    to_unsigned(2133918078,32),
    to_unsigned(2133941174,32),
    to_unsigned(2133964250,32),
    to_unsigned(2133987306,32),
    to_unsigned(2134010343,32),
    to_unsigned(2134033360,32),
    to_unsigned(2134056357,32),
    to_unsigned(2134079335,32),
    to_unsigned(2134102293,32),
    to_unsigned(2134125232,32),
    to_unsigned(2134148151,32),
    to_unsigned(2134171050,32),
    to_unsigned(2134193930,32),
    to_unsigned(2134216790,32),
    to_unsigned(2134239631,32),
    to_unsigned(2134262451,32),
    to_unsigned(2134285253,32),
    to_unsigned(2134308034,32),
    to_unsigned(2134330796,32),
    to_unsigned(2134353539,32),
    to_unsigned(2134376262,32),
    to_unsigned(2134398965,32),
    to_unsigned(2134421648,32),
    to_unsigned(2134444312,32),
    to_unsigned(2134466957,32),
    to_unsigned(2134489581,32),
    to_unsigned(2134512186,32),
    to_unsigned(2134534772,32),
    to_unsigned(2134557338,32),
    to_unsigned(2134579884,32),
    to_unsigned(2134602410,32),
    to_unsigned(2134624917,32),
    to_unsigned(2134647405,32),
    to_unsigned(2134669872,32),
    to_unsigned(2134692321,32),
    to_unsigned(2134714749,32),
    to_unsigned(2134737158,32),
    to_unsigned(2134759547,32),
    to_unsigned(2134781917,32),
    to_unsigned(2134804267,32),
    to_unsigned(2134826597,32),
    to_unsigned(2134848908,32),
    to_unsigned(2134871199,32),
    to_unsigned(2134893471,32),
    to_unsigned(2134915722,32),
    to_unsigned(2134937955,32),
    to_unsigned(2134960167,32),
    to_unsigned(2134982360,32),
    to_unsigned(2135004534,32),
    to_unsigned(2135026688,32),
    to_unsigned(2135048822,32),
    to_unsigned(2135070936,32),
    to_unsigned(2135093031,32),
    to_unsigned(2135115106,32),
    to_unsigned(2135137162,32),
    to_unsigned(2135159198,32),
    to_unsigned(2135181214,32),
    to_unsigned(2135203211,32),
    to_unsigned(2135225188,32),
    to_unsigned(2135247146,32),
    to_unsigned(2135269084,32),
    to_unsigned(2135291002,32),
    to_unsigned(2135312901,32),
    to_unsigned(2135334780,32),
    to_unsigned(2135356639,32),
    to_unsigned(2135378479,32),
    to_unsigned(2135400299,32),
    to_unsigned(2135422099,32),
    to_unsigned(2135443880,32),
    to_unsigned(2135465641,32),
    to_unsigned(2135487383,32),
    to_unsigned(2135509105,32),
    to_unsigned(2135530807,32),
    to_unsigned(2135552490,32),
    to_unsigned(2135574153,32),
    to_unsigned(2135595797,32),
    to_unsigned(2135617420,32),
    to_unsigned(2135639025,32),
    to_unsigned(2135660609,32),
    to_unsigned(2135682174,32),
    to_unsigned(2135703719,32),
    to_unsigned(2135725245,32),
    to_unsigned(2135746751,32),
    to_unsigned(2135768238,32),
    to_unsigned(2135789704,32),
    to_unsigned(2135811152,32),
    to_unsigned(2135832579,32),
    to_unsigned(2135853987,32),
    to_unsigned(2135875375,32),
    to_unsigned(2135896744,32),
    to_unsigned(2135918093,32),
    to_unsigned(2135939422,32),
    to_unsigned(2135960732,32),
    to_unsigned(2135982022,32),
    to_unsigned(2136003292,32),
    to_unsigned(2136024543,32),
    to_unsigned(2136045774,32),
    to_unsigned(2136066986,32),
    to_unsigned(2136088178,32),
    to_unsigned(2136109350,32),
    to_unsigned(2136130503,32),
    to_unsigned(2136151636,32),
    to_unsigned(2136172749,32),
    to_unsigned(2136193843,32),
    to_unsigned(2136214917,32),
    to_unsigned(2136235972,32),
    to_unsigned(2136257006,32),
    to_unsigned(2136278022,32),
    to_unsigned(2136299017,32),
    to_unsigned(2136319993,32),
    to_unsigned(2136340949,32),
    to_unsigned(2136361886,32),
    to_unsigned(2136382803,32),
    to_unsigned(2136403700,32),
    to_unsigned(2136424578,32),
    to_unsigned(2136445436,32),
    to_unsigned(2136466275,32),
    to_unsigned(2136487094,32),
    to_unsigned(2136507893,32),
    to_unsigned(2136528672,32),
    to_unsigned(2136549432,32),
    to_unsigned(2136570173,32),
    to_unsigned(2136590893,32),
    to_unsigned(2136611594,32),
    to_unsigned(2136632276,32),
    to_unsigned(2136652937,32),
    to_unsigned(2136673579,32),
    to_unsigned(2136694202,32),
    to_unsigned(2136714805,32),
    to_unsigned(2136735388,32),
    to_unsigned(2136755951,32),
    to_unsigned(2136776495,32),
    to_unsigned(2136797019,32),
    to_unsigned(2136817524,32),
    to_unsigned(2136838009,32),
    to_unsigned(2136858474,32),
    to_unsigned(2136878920,32),
    to_unsigned(2136899346,32),
    to_unsigned(2136919752,32),
    to_unsigned(2136940139,32),
    to_unsigned(2136960506,32),
    to_unsigned(2136980854,32),
    to_unsigned(2137001182,32),
    to_unsigned(2137021490,32),
    to_unsigned(2137041778,32),
    to_unsigned(2137062047,32),
    to_unsigned(2137082296,32),
    to_unsigned(2137102526,32),
    to_unsigned(2137122736,32),
    to_unsigned(2137142926,32),
    to_unsigned(2137163097,32),
    to_unsigned(2137183248,32),
    to_unsigned(2137203379,32),
    to_unsigned(2137223491,32),
    to_unsigned(2137243583,32),
    to_unsigned(2137263656,32),
    to_unsigned(2137283708,32),
    to_unsigned(2137303742,32),
    to_unsigned(2137323755,32),
    to_unsigned(2137343749,32),
    to_unsigned(2137363723,32),
    to_unsigned(2137383678,32),
    to_unsigned(2137403613,32),
    to_unsigned(2137423528,32),
    to_unsigned(2137443424,32),
    to_unsigned(2137463300,32),
    to_unsigned(2137483156,32),
    to_unsigned(2137502993,32),
    to_unsigned(2137522810,32),
    to_unsigned(2137542607,32),
    to_unsigned(2137562385,32),
    to_unsigned(2137582143,32),
    to_unsigned(2137601881,32),
    to_unsigned(2137621600,32),
    to_unsigned(2137641299,32),
    to_unsigned(2137660979,32),
    to_unsigned(2137680639,32),
    to_unsigned(2137700279,32),
    to_unsigned(2137719900,32),
    to_unsigned(2137739500,32),
    to_unsigned(2137759082,32),
    to_unsigned(2137778643,32),
    to_unsigned(2137798185,32),
    to_unsigned(2137817708,32),
    to_unsigned(2137837210,32),
    to_unsigned(2137856693,32),
    to_unsigned(2137876157,32),
    to_unsigned(2137895600,32),
    to_unsigned(2137915024,32),
    to_unsigned(2137934429,32),
    to_unsigned(2137953814,32),
    to_unsigned(2137973179,32),
    to_unsigned(2137992524,32),
    to_unsigned(2138011850,32),
    to_unsigned(2138031156,32),
    to_unsigned(2138050443,32),
    to_unsigned(2138069709,32),
    to_unsigned(2138088957,32),
    to_unsigned(2138108184,32),
    to_unsigned(2138127392,32),
    to_unsigned(2138146580,32),
    to_unsigned(2138165749,32),
    to_unsigned(2138184898,32),
    to_unsigned(2138204027,32),
    to_unsigned(2138223137,32),
    to_unsigned(2138242227,32),
    to_unsigned(2138261297,32),
    to_unsigned(2138280348,32),
    to_unsigned(2138299379,32),
    to_unsigned(2138318390,32),
    to_unsigned(2138337382,32),
    to_unsigned(2138356354,32),
    to_unsigned(2138375306,32),
    to_unsigned(2138394239,32),
    to_unsigned(2138413152,32),
    to_unsigned(2138432045,32),
    to_unsigned(2138450919,32),
    to_unsigned(2138469773,32),
    to_unsigned(2138488608,32),
    to_unsigned(2138507422,32),
    to_unsigned(2138526217,32),
    to_unsigned(2138544993,32),
    to_unsigned(2138563749,32),
    to_unsigned(2138582485,32),
    to_unsigned(2138601201,32),
    to_unsigned(2138619898,32),
    to_unsigned(2138638575,32),
    to_unsigned(2138657233,32),
    to_unsigned(2138675871,32),
    to_unsigned(2138694489,32),
    to_unsigned(2138713088,32),
    to_unsigned(2138731667,32),
    to_unsigned(2138750226,32),
    to_unsigned(2138768765,32),
    to_unsigned(2138787285,32),
    to_unsigned(2138805786,32),
    to_unsigned(2138824266,32),
    to_unsigned(2138842727,32),
    to_unsigned(2138861168,32),
    to_unsigned(2138879590,32),
    to_unsigned(2138897992,32),
    to_unsigned(2138916374,32),
    to_unsigned(2138934737,32),
    to_unsigned(2138953080,32),
    to_unsigned(2138971403,32),
    to_unsigned(2138989707,32),
    to_unsigned(2139007991,32),
    to_unsigned(2139026255,32),
    to_unsigned(2139044500,32),
    to_unsigned(2139062725,32),
    to_unsigned(2139080930,32),
    to_unsigned(2139099116,32),
    to_unsigned(2139117282,32),
    to_unsigned(2139135428,32),
    to_unsigned(2139153555,32),
    to_unsigned(2139171662,32),
    to_unsigned(2139189749,32),
    to_unsigned(2139207817,32),
    to_unsigned(2139225865,32),
    to_unsigned(2139243894,32),
    to_unsigned(2139261902,32),
    to_unsigned(2139279891,32),
    to_unsigned(2139297861,32),
    to_unsigned(2139315811,32),
    to_unsigned(2139333741,32),
    to_unsigned(2139351651,32),
    to_unsigned(2139369542,32),
    to_unsigned(2139387413,32),
    to_unsigned(2139405264,32),
    to_unsigned(2139423096,32),
    to_unsigned(2139440908,32),
    to_unsigned(2139458700,32),
    to_unsigned(2139476473,32),
    to_unsigned(2139494226,32),
    to_unsigned(2139511960,32),
    to_unsigned(2139529673,32),
    to_unsigned(2139547368,32),
    to_unsigned(2139565042,32),
    to_unsigned(2139582697,32),
    to_unsigned(2139600332,32),
    to_unsigned(2139617947,32),
    to_unsigned(2139635543,32),
    to_unsigned(2139653119,32),
    to_unsigned(2139670675,32),
    to_unsigned(2139688212,32),
    to_unsigned(2139705729,32),
    to_unsigned(2139723227,32),
    to_unsigned(2139740704,32),
    to_unsigned(2139758163,32),
    to_unsigned(2139775601,32),
    to_unsigned(2139793020,32),
    to_unsigned(2139810419,32),
    to_unsigned(2139827798,32),
    to_unsigned(2139845158,32),
    to_unsigned(2139862498,32),
    to_unsigned(2139879818,32),
    to_unsigned(2139897119,32),
    to_unsigned(2139914400,32),
    to_unsigned(2139931662,32),
    to_unsigned(2139948903,32),
    to_unsigned(2139966125,32),
    to_unsigned(2139983328,32),
    to_unsigned(2140000510,32),
    to_unsigned(2140017673,32),
    to_unsigned(2140034817,32),
    to_unsigned(2140051941,32),
    to_unsigned(2140069045,32),
    to_unsigned(2140086129,32),
    to_unsigned(2140103194,32),
    to_unsigned(2140120239,32),
    to_unsigned(2140137264,32),
    to_unsigned(2140154270,32),
    to_unsigned(2140171256,32),
    to_unsigned(2140188222,32),
    to_unsigned(2140205169,32),
    to_unsigned(2140222096,32),
    to_unsigned(2140239003,32),
    to_unsigned(2140255891,32),
    to_unsigned(2140272759,32),
    to_unsigned(2140289607,32),
    to_unsigned(2140306435,32),
    to_unsigned(2140323244,32),
    to_unsigned(2140340034,32),
    to_unsigned(2140356803,32),
    to_unsigned(2140373553,32),
    to_unsigned(2140390283,32),
    to_unsigned(2140406994,32),
    to_unsigned(2140423685,32),
    to_unsigned(2140440356,32),
    to_unsigned(2140457008,32),
    to_unsigned(2140473640,32),
    to_unsigned(2140490252,32),
    to_unsigned(2140506844,32),
    to_unsigned(2140523417,32),
    to_unsigned(2140539970,32),
    to_unsigned(2140556504,32),
    to_unsigned(2140573018,32),
    to_unsigned(2140589512,32),
    to_unsigned(2140605986,32),
    to_unsigned(2140622441,32),
    to_unsigned(2140638876,32),
    to_unsigned(2140655292,32),
    to_unsigned(2140671687,32),
    to_unsigned(2140688064,32),
    to_unsigned(2140704420,32),
    to_unsigned(2140720757,32),
    to_unsigned(2140737074,32),
    to_unsigned(2140753371,32),
    to_unsigned(2140769649,32),
    to_unsigned(2140785907,32),
    to_unsigned(2140802145,32),
    to_unsigned(2140818364,32),
    to_unsigned(2140834563,32),
    to_unsigned(2140850742,32),
    to_unsigned(2140866902,32),
    to_unsigned(2140883042,32),
    to_unsigned(2140899162,32),
    to_unsigned(2140915263,32),
    to_unsigned(2140931344,32),
    to_unsigned(2140947405,32),
    to_unsigned(2140963447,32),
    to_unsigned(2140979468,32),
    to_unsigned(2140995471,32),
    to_unsigned(2141011453,32),
    to_unsigned(2141027416,32),
    to_unsigned(2141043359,32),
    to_unsigned(2141059283,32),
    to_unsigned(2141075187,32),
    to_unsigned(2141091071,32),
    to_unsigned(2141106935,32),
    to_unsigned(2141122780,32),
    to_unsigned(2141138605,32),
    to_unsigned(2141154410,32),
    to_unsigned(2141170196,32),
    to_unsigned(2141185962,32),
    to_unsigned(2141201709,32),
    to_unsigned(2141217435,32),
    to_unsigned(2141233142,32),
    to_unsigned(2141248830,32),
    to_unsigned(2141264497,32),
    to_unsigned(2141280145,32),
    to_unsigned(2141295773,32),
    to_unsigned(2141311382,32),
    to_unsigned(2141326971,32),
    to_unsigned(2141342540,32),
    to_unsigned(2141358090,32),
    to_unsigned(2141373620,32),
    to_unsigned(2141389130,32),
    to_unsigned(2141404620,32),
    to_unsigned(2141420091,32),
    to_unsigned(2141435542,32),
    to_unsigned(2141450974,32),
    to_unsigned(2141466385,32),
    to_unsigned(2141481777,32),
    to_unsigned(2141497150,32),
    to_unsigned(2141512503,32),
    to_unsigned(2141527836,32),
    to_unsigned(2141543149,32),
    to_unsigned(2141558443,32),
    to_unsigned(2141573717,32),
    to_unsigned(2141588971,32),
    to_unsigned(2141604205,32),
    to_unsigned(2141619420,32),
    to_unsigned(2141634616,32),
    to_unsigned(2141649791,32),
    to_unsigned(2141664947,32),
    to_unsigned(2141680083,32),
    to_unsigned(2141695200,32),
    to_unsigned(2141710296,32),
    to_unsigned(2141725374,32),
    to_unsigned(2141740431,32),
    to_unsigned(2141755469,32),
    to_unsigned(2141770487,32),
    to_unsigned(2141785485,32),
    to_unsigned(2141800464,32),
    to_unsigned(2141815423,32),
    to_unsigned(2141830362,32),
    to_unsigned(2141845282,32),
    to_unsigned(2141860182,32),
    to_unsigned(2141875062,32),
    to_unsigned(2141889923,32),
    to_unsigned(2141904763,32),
    to_unsigned(2141919585,32),
    to_unsigned(2141934386,32),
    to_unsigned(2141949168,32),
    to_unsigned(2141963930,32),
    to_unsigned(2141978672,32),
    to_unsigned(2141993395,32),
    to_unsigned(2142008098,32),
    to_unsigned(2142022782,32),
    to_unsigned(2142037445,32),
    to_unsigned(2142052089,32),
    to_unsigned(2142066714,32),
    to_unsigned(2142081318,32),
    to_unsigned(2142095903,32),
    to_unsigned(2142110468,32),
    to_unsigned(2142125014,32),
    to_unsigned(2142139540,32),
    to_unsigned(2142154046,32),
    to_unsigned(2142168532,32),
    to_unsigned(2142182999,32),
    to_unsigned(2142197446,32),
    to_unsigned(2142211874,32),
    to_unsigned(2142226281,32),
    to_unsigned(2142240669,32),
    to_unsigned(2142255038,32),
    to_unsigned(2142269386,32),
    to_unsigned(2142283715,32),
    to_unsigned(2142298025,32),
    to_unsigned(2142312314,32),
    to_unsigned(2142326584,32),
    to_unsigned(2142340834,32),
    to_unsigned(2142355065,32),
    to_unsigned(2142369275,32),
    to_unsigned(2142383467,32),
    to_unsigned(2142397638,32),
    to_unsigned(2142411790,32),
    to_unsigned(2142425922,32),
    to_unsigned(2142440034,32),
    to_unsigned(2142454127,32),
    to_unsigned(2142468200,32),
    to_unsigned(2142482253,32),
    to_unsigned(2142496286,32),
    to_unsigned(2142510300,32),
    to_unsigned(2142524294,32),
    to_unsigned(2142538269,32),
    to_unsigned(2142552224,32),
    to_unsigned(2142566159,32),
    to_unsigned(2142580074,32),
    to_unsigned(2142593970,32),
    to_unsigned(2142607846,32),
    to_unsigned(2142621702,32),
    to_unsigned(2142635539,32),
    to_unsigned(2142649356,32),
    to_unsigned(2142663153,32),
    to_unsigned(2142676930,32),
    to_unsigned(2142690688,32),
    to_unsigned(2142704426,32),
    to_unsigned(2142718145,32),
    to_unsigned(2142731844,32),
    to_unsigned(2142745523,32),
    to_unsigned(2142759182,32),
    to_unsigned(2142772822,32),
    to_unsigned(2142786442,32),
    to_unsigned(2142800042,32),
    to_unsigned(2142813623,32),
    to_unsigned(2142827183,32),
    to_unsigned(2142840725,32),
    to_unsigned(2142854246,32),
    to_unsigned(2142867748,32),
    to_unsigned(2142881230,32),
    to_unsigned(2142894692,32),
    to_unsigned(2142908135,32),
    to_unsigned(2142921558,32),
    to_unsigned(2142934961,32),
    to_unsigned(2142948345,32),
    to_unsigned(2142961709,32),
    to_unsigned(2142975053,32),
    to_unsigned(2142988378,32),
    to_unsigned(2143001682,32),
    to_unsigned(2143014968,32),
    to_unsigned(2143028233,32),
    to_unsigned(2143041479,32),
    to_unsigned(2143054705,32),
    to_unsigned(2143067911,32),
    to_unsigned(2143081098,32),
    to_unsigned(2143094265,32),
    to_unsigned(2143107412,32),
    to_unsigned(2143120539,32),
    to_unsigned(2143133647,32),
    to_unsigned(2143146735,32),
    to_unsigned(2143159804,32),
    to_unsigned(2143172853,32),
    to_unsigned(2143185882,32),
    to_unsigned(2143198891,32),
    to_unsigned(2143211881,32),
    to_unsigned(2143224851,32),
    to_unsigned(2143237801,32),
    to_unsigned(2143250731,32),
    to_unsigned(2143263642,32),
    to_unsigned(2143276533,32),
    to_unsigned(2143289405,32),
    to_unsigned(2143302256,32),
    to_unsigned(2143315088,32),
    to_unsigned(2143327901,32),
    to_unsigned(2143340693,32),
    to_unsigned(2143353466,32),
    to_unsigned(2143366220,32),
    to_unsigned(2143378953,32),
    to_unsigned(2143391667,32),
    to_unsigned(2143404361,32),
    to_unsigned(2143417035,32),
    to_unsigned(2143429690,32),
    to_unsigned(2143442325,32),
    to_unsigned(2143454941,32),
    to_unsigned(2143467536,32),
    to_unsigned(2143480112,32),
    to_unsigned(2143492668,32),
    to_unsigned(2143505205,32),
    to_unsigned(2143517722,32),
    to_unsigned(2143530219,32),
    to_unsigned(2143542696,32),
    to_unsigned(2143555154,32),
    to_unsigned(2143567592,32),
    to_unsigned(2143580010,32),
    to_unsigned(2143592409,32),
    to_unsigned(2143604788,32),
    to_unsigned(2143617147,32),
    to_unsigned(2143629486,32),
    to_unsigned(2143641806,32),
    to_unsigned(2143654106,32),
    to_unsigned(2143666386,32),
    to_unsigned(2143678647,32),
    to_unsigned(2143690888,32),
    to_unsigned(2143703109,32),
    to_unsigned(2143715311,32),
    to_unsigned(2143727493,32),
    to_unsigned(2143739655,32),
    to_unsigned(2143751797,32),
    to_unsigned(2143763920,32),
    to_unsigned(2143776023,32),
    to_unsigned(2143788106,32),
    to_unsigned(2143800170,32),
    to_unsigned(2143812214,32),
    to_unsigned(2143824238,32),
    to_unsigned(2143836243,32),
    to_unsigned(2143848227,32),
    to_unsigned(2143860192,32),
    to_unsigned(2143872138,32),
    to_unsigned(2143884063,32),
    to_unsigned(2143895969,32),
    to_unsigned(2143907856,32),
    to_unsigned(2143919722,32),
    to_unsigned(2143931569,32),
    to_unsigned(2143943396,32),
    to_unsigned(2143955204,32),
    to_unsigned(2143966991,32),
    to_unsigned(2143978759,32),
    to_unsigned(2143990508,32),
    to_unsigned(2144002236,32),
    to_unsigned(2144013945,32),
    to_unsigned(2144025634,32),
    to_unsigned(2144037304,32),
    to_unsigned(2144048954,32),
    to_unsigned(2144060584,32),
    to_unsigned(2144072194,32),
    to_unsigned(2144083785,32),
    to_unsigned(2144095356,32),
    to_unsigned(2144106907,32),
    to_unsigned(2144118438,32),
    to_unsigned(2144129950,32),
    to_unsigned(2144141442,32),
    to_unsigned(2144152915,32),
    to_unsigned(2144164368,32),
    to_unsigned(2144175801,32),
    to_unsigned(2144187214,32),
    to_unsigned(2144198607,32),
    to_unsigned(2144209981,32),
    to_unsigned(2144221335,32),
    to_unsigned(2144232670,32),
    to_unsigned(2144243985,32),
    to_unsigned(2144255280,32),
    to_unsigned(2144266555,32),
    to_unsigned(2144277810,32),
    to_unsigned(2144289046,32),
    to_unsigned(2144300263,32),
    to_unsigned(2144311459,32),
    to_unsigned(2144322636,32),
    to_unsigned(2144333793,32),
    to_unsigned(2144344930,32),
    to_unsigned(2144356048,32),
    to_unsigned(2144367146,32),
    to_unsigned(2144378224,32),
    to_unsigned(2144389282,32),
    to_unsigned(2144400321,32),
    to_unsigned(2144411340,32),
    to_unsigned(2144422340,32),
    to_unsigned(2144433319,32),
    to_unsigned(2144444279,32),
    to_unsigned(2144455220,32),
    to_unsigned(2144466140,32),
    to_unsigned(2144477041,32),
    to_unsigned(2144487922,32),
    to_unsigned(2144498783,32),
    to_unsigned(2144509625,32),
    to_unsigned(2144520447,32),
    to_unsigned(2144531249,32),
    to_unsigned(2144542032,32),
    to_unsigned(2144552795,32),
    to_unsigned(2144563538,32),
    to_unsigned(2144574261,32),
    to_unsigned(2144584965,32),
    to_unsigned(2144595649,32),
    to_unsigned(2144606313,32),
    to_unsigned(2144616958,32),
    to_unsigned(2144627583,32),
    to_unsigned(2144638188,32),
    to_unsigned(2144648773,32),
    to_unsigned(2144659339,32),
    to_unsigned(2144669885,32),
    to_unsigned(2144680411,32),
    to_unsigned(2144690918,32),
    to_unsigned(2144701404,32),
    to_unsigned(2144711872,32),
    to_unsigned(2144722319,32),
    to_unsigned(2144732747,32),
    to_unsigned(2144743155,32),
    to_unsigned(2144753543,32),
    to_unsigned(2144763912,32),
    to_unsigned(2144774260,32),
    to_unsigned(2144784590,32),
    to_unsigned(2144794899,32),
    to_unsigned(2144805189,32),
    to_unsigned(2144815459,32),
    to_unsigned(2144825709,32),
    to_unsigned(2144835940,32),
    to_unsigned(2144846150,32),
    to_unsigned(2144856342,32),
    to_unsigned(2144866513,32),
    to_unsigned(2144876665,32),
    to_unsigned(2144886797,32),
    to_unsigned(2144896909,32),
    to_unsigned(2144907001,32),
    to_unsigned(2144917074,32),
    to_unsigned(2144927127,32),
    to_unsigned(2144937161,32),
    to_unsigned(2144947175,32),
    to_unsigned(2144957169,32),
    to_unsigned(2144967143,32),
    to_unsigned(2144977097,32),
    to_unsigned(2144987032,32),
    to_unsigned(2144996947,32),
    to_unsigned(2145006843,32),
    to_unsigned(2145016718,32),
    to_unsigned(2145026574,32),
    to_unsigned(2145036411,32),
    to_unsigned(2145046227,32),
    to_unsigned(2145056024,32),
    to_unsigned(2145065801,32),
    to_unsigned(2145075558,32),
    to_unsigned(2145085296,32),
    to_unsigned(2145095014,32),
    to_unsigned(2145104712,32),
    to_unsigned(2145114391,32),
    to_unsigned(2145124050,32),
    to_unsigned(2145133689,32),
    to_unsigned(2145143308,32),
    to_unsigned(2145152908,32),
    to_unsigned(2145162488,32),
    to_unsigned(2145172048,32),
    to_unsigned(2145181588,32),
    to_unsigned(2145191109,32),
    to_unsigned(2145200610,32),
    to_unsigned(2145210091,32),
    to_unsigned(2145219553,32),
    to_unsigned(2145228995,32),
    to_unsigned(2145238417,32),
    to_unsigned(2145247820,32),
    to_unsigned(2145257202,32),
    to_unsigned(2145266565,32),
    to_unsigned(2145275909,32),
    to_unsigned(2145285232,32),
    to_unsigned(2145294536,32),
    to_unsigned(2145303820,32),
    to_unsigned(2145313085,32),
    to_unsigned(2145322329,32),
    to_unsigned(2145331554,32),
    to_unsigned(2145340760,32),
    to_unsigned(2145349945,32),
    to_unsigned(2145359111,32),
    to_unsigned(2145368257,32),
    to_unsigned(2145377384,32),
    to_unsigned(2145386490,32),
    to_unsigned(2145395577,32),
    to_unsigned(2145404644,32),
    to_unsigned(2145413692,32),
    to_unsigned(2145422720,32),
    to_unsigned(2145431728,32),
    to_unsigned(2145440716,32),
    to_unsigned(2145449685,32),
    to_unsigned(2145458634,32),
    to_unsigned(2145467563,32),
    to_unsigned(2145476472,32),
    to_unsigned(2145485362,32),
    to_unsigned(2145494232,32),
    to_unsigned(2145503082,32),
    to_unsigned(2145511913,32),
    to_unsigned(2145520724,32),
    to_unsigned(2145529515,32),
    to_unsigned(2145538286,32),
    to_unsigned(2145547038,32),
    to_unsigned(2145555770,32),
    to_unsigned(2145564482,32),
    to_unsigned(2145573175,32),
    to_unsigned(2145581848,32),
    to_unsigned(2145590501,32),
    to_unsigned(2145599134,32),
    to_unsigned(2145607748,32),
    to_unsigned(2145616342,32),
    to_unsigned(2145624916,32),
    to_unsigned(2145633470,32),
    to_unsigned(2145642005,32),
    to_unsigned(2145650520,32),
    to_unsigned(2145659016,32),
    to_unsigned(2145667491,32),
    to_unsigned(2145675947,32),
    to_unsigned(2145684383,32),
    to_unsigned(2145692800,32),
    to_unsigned(2145701196,32),
    to_unsigned(2145709573,32),
    to_unsigned(2145717931,32),
    to_unsigned(2145726268,32),
    to_unsigned(2145734586,32),
    to_unsigned(2145742884,32),
    to_unsigned(2145751162,32),
    to_unsigned(2145759421,32),
    to_unsigned(2145767660,32),
    to_unsigned(2145775879,32),
    to_unsigned(2145784079,32),
    to_unsigned(2145792258,32),
    to_unsigned(2145800418,32),
    to_unsigned(2145808559,32),
    to_unsigned(2145816679,32),
    to_unsigned(2145824780,32),
    to_unsigned(2145832861,32),
    to_unsigned(2145840923,32),
    to_unsigned(2145848964,32),
    to_unsigned(2145856986,32),
    to_unsigned(2145864989,32),
    to_unsigned(2145872971,32),
    to_unsigned(2145880934,32),
    to_unsigned(2145888877,32),
    to_unsigned(2145896800,32),
    to_unsigned(2145904704,32),
    to_unsigned(2145912588,32),
    to_unsigned(2145920452,32),
    to_unsigned(2145928296,32),
    to_unsigned(2145936121,32),
    to_unsigned(2145943926,32),
    to_unsigned(2145951711,32),
    to_unsigned(2145959477,32),
    to_unsigned(2145967223,32),
    to_unsigned(2145974949,32),
    to_unsigned(2145982655,32),
    to_unsigned(2145990342,32),
    to_unsigned(2145998009,32),
    to_unsigned(2146005656,32),
    to_unsigned(2146013283,32),
    to_unsigned(2146020891,32),
    to_unsigned(2146028479,32),
    to_unsigned(2146036047,32),
    to_unsigned(2146043596,32),
    to_unsigned(2146051125,32),
    to_unsigned(2146058634,32),
    to_unsigned(2146066123,32),
    to_unsigned(2146073593,32),
    to_unsigned(2146081043,32),
    to_unsigned(2146088473,32),
    to_unsigned(2146095883,32),
    to_unsigned(2146103274,32),
    to_unsigned(2146110645,32),
    to_unsigned(2146117996,32),
    to_unsigned(2146125328,32),
    to_unsigned(2146132640,32),
    to_unsigned(2146139932,32),
    to_unsigned(2146147204,32),
    to_unsigned(2146154457,32),
    to_unsigned(2146161690,32),
    to_unsigned(2146168903,32),
    to_unsigned(2146176097,32),
    to_unsigned(2146183270,32),
    to_unsigned(2146190424,32),
    to_unsigned(2146197559,32),
    to_unsigned(2146204673,32),
    to_unsigned(2146211768,32),
    to_unsigned(2146218843,32),
    to_unsigned(2146225899,32),
    to_unsigned(2146232934,32),
    to_unsigned(2146239950,32),
    to_unsigned(2146246946,32),
    to_unsigned(2146253923,32),
    to_unsigned(2146260880,32),
    to_unsigned(2146267817,32),
    to_unsigned(2146274734,32),
    to_unsigned(2146281631,32),
    to_unsigned(2146288509,32),
    to_unsigned(2146295367,32),
    to_unsigned(2146302206,32),
    to_unsigned(2146309024,32),
    to_unsigned(2146315823,32),
    to_unsigned(2146322603,32),
    to_unsigned(2146329362,32),
    to_unsigned(2146336102,32),
    to_unsigned(2146342822,32),
    to_unsigned(2146349522,32),
    to_unsigned(2146356203,32),
    to_unsigned(2146362863,32),
    to_unsigned(2146369504,32),
    to_unsigned(2146376126,32),
    to_unsigned(2146382727,32),
    to_unsigned(2146389309,32),
    to_unsigned(2146395872,32),
    to_unsigned(2146402414,32),
    to_unsigned(2146408937,32),
    to_unsigned(2146415440,32),
    to_unsigned(2146421923,32),
    to_unsigned(2146428387,32),
    to_unsigned(2146434830,32),
    to_unsigned(2146441254,32),
    to_unsigned(2146447659,32),
    to_unsigned(2146454043,32),
    to_unsigned(2146460408,32),
    to_unsigned(2146466753,32),
    to_unsigned(2146473079,32),
    to_unsigned(2146479384,32),
    to_unsigned(2146485670,32),
    to_unsigned(2146491937,32),
    to_unsigned(2146498183,32),
    to_unsigned(2146504410,32),
    to_unsigned(2146510617,32),
    to_unsigned(2146516804,32),
    to_unsigned(2146522972,32),
    to_unsigned(2146529120,32),
    to_unsigned(2146535248,32),
    to_unsigned(2146541356,32),
    to_unsigned(2146547445,32),
    to_unsigned(2146553514,32),
    to_unsigned(2146559563,32),
    to_unsigned(2146565592,32),
    to_unsigned(2146571602,32),
    to_unsigned(2146577592,32),
    to_unsigned(2146583562,32),
    to_unsigned(2146589513,32),
    to_unsigned(2146595444,32),
    to_unsigned(2146601355,32),
    to_unsigned(2146607246,32),
    to_unsigned(2146613118,32),
    to_unsigned(2146618970,32),
    to_unsigned(2146624802,32),
    to_unsigned(2146630614,32),
    to_unsigned(2146636407,32),
    to_unsigned(2146642180,32),
    to_unsigned(2146647933,32),
    to_unsigned(2146653667,32),
    to_unsigned(2146659381,32),
    to_unsigned(2146665075,32),
    to_unsigned(2146670749,32),
    to_unsigned(2146676403,32),
    to_unsigned(2146682038,32),
    to_unsigned(2146687653,32),
    to_unsigned(2146693249,32),
    to_unsigned(2146698824,32),
    to_unsigned(2146704380,32),
    to_unsigned(2146709916,32),
    to_unsigned(2146715433,32),
    to_unsigned(2146720930,32),
    to_unsigned(2146726407,32),
    to_unsigned(2146731864,32),
    to_unsigned(2146737301,32),
    to_unsigned(2146742719,32),
    to_unsigned(2146748117,32),
    to_unsigned(2146753496,32),
    to_unsigned(2146758854,32),
    to_unsigned(2146764193,32),
    to_unsigned(2146769512,32),
    to_unsigned(2146774812,32),
    to_unsigned(2146780091,32),
    to_unsigned(2146785351,32),
    to_unsigned(2146790591,32),
    to_unsigned(2146795812,32),
    to_unsigned(2146801013,32),
    to_unsigned(2146806193,32),
    to_unsigned(2146811355,32),
    to_unsigned(2146816496,32),
    to_unsigned(2146821618,32),
    to_unsigned(2146826720,32),
    to_unsigned(2146831802,32),
    to_unsigned(2146836865,32),
    to_unsigned(2146841908,32),
    to_unsigned(2146846931,32),
    to_unsigned(2146851934,32),
    to_unsigned(2146856918,32),
    to_unsigned(2146861882,32),
    to_unsigned(2146866826,32),
    to_unsigned(2146871751,32),
    to_unsigned(2146876655,32),
    to_unsigned(2146881540,32),
    to_unsigned(2146886406,32),
    to_unsigned(2146891251,32),
    to_unsigned(2146896077,32),
    to_unsigned(2146900883,32),
    to_unsigned(2146905669,32),
    to_unsigned(2146910436,32),
    to_unsigned(2146915183,32),
    to_unsigned(2146919910,32),
    to_unsigned(2146924617,32),
    to_unsigned(2146929305,32),
    to_unsigned(2146933973,32),
    to_unsigned(2146938621,32),
    to_unsigned(2146943250,32),
    to_unsigned(2146947858,32),
    to_unsigned(2146952447,32),
    to_unsigned(2146957017,32),
    to_unsigned(2146961566,32),
    to_unsigned(2146966096,32),
    to_unsigned(2146970606,32),
    to_unsigned(2146975096,32),
    to_unsigned(2146979567,32),
    to_unsigned(2146984018,32),
    to_unsigned(2146988449,32),
    to_unsigned(2146992860,32),
    to_unsigned(2146997252,32),
    to_unsigned(2147001624,32),
    to_unsigned(2147005976,32),
    to_unsigned(2147010308,32),
    to_unsigned(2147014621,32),
    to_unsigned(2147018914,32),
    to_unsigned(2147023187,32),
    to_unsigned(2147027441,32),
    to_unsigned(2147031674,32),
    to_unsigned(2147035888,32),
    to_unsigned(2147040083,32),
    to_unsigned(2147044257,32),
    to_unsigned(2147048412,32),
    to_unsigned(2147052547,32),
    to_unsigned(2147056663,32),
    to_unsigned(2147060758,32),
    to_unsigned(2147064834,32),
    to_unsigned(2147068890,32),
    to_unsigned(2147072927,32),
    to_unsigned(2147076943,32),
    to_unsigned(2147080940,32),
    to_unsigned(2147084917,32),
    to_unsigned(2147088875,32),
    to_unsigned(2147092813,32),
    to_unsigned(2147096731,32),
    to_unsigned(2147100629,32),
    to_unsigned(2147104507,32),
    to_unsigned(2147108366,32),
    to_unsigned(2147112205,32),
    to_unsigned(2147116025,32),
    to_unsigned(2147119824,32),
    to_unsigned(2147123604,32),
    to_unsigned(2147127364,32),
    to_unsigned(2147131105,32),
    to_unsigned(2147134825,32),
    to_unsigned(2147138526,32),
    to_unsigned(2147142207,32),
    to_unsigned(2147145869,32),
    to_unsigned(2147149510,32),
    to_unsigned(2147153132,32),
    to_unsigned(2147156735,32),
    to_unsigned(2147160317,32),
    to_unsigned(2147163880,32),
    to_unsigned(2147167423,32),
    to_unsigned(2147170946,32),
    to_unsigned(2147174450,32),
    to_unsigned(2147177933,32),
    to_unsigned(2147181397,32),
    to_unsigned(2147184842,32),
    to_unsigned(2147188266,32),
    to_unsigned(2147191671,32),
    to_unsigned(2147195056,32),
    to_unsigned(2147198422,32),
    to_unsigned(2147201767,32),
    to_unsigned(2147205093,32),
    to_unsigned(2147208399,32),
    to_unsigned(2147211686,32),
    to_unsigned(2147214953,32),
    to_unsigned(2147218200,32),
    to_unsigned(2147221427,32),
    to_unsigned(2147224634,32),
    to_unsigned(2147227822,32),
    to_unsigned(2147230990,32),
    to_unsigned(2147234138,32),
    to_unsigned(2147237267,32),
    to_unsigned(2147240376,32),
    to_unsigned(2147243465,32),
    to_unsigned(2147246534,32),
    to_unsigned(2147249584,32),
    to_unsigned(2147252614,32),
    to_unsigned(2147255624,32),
    to_unsigned(2147258614,32),
    to_unsigned(2147261585,32),
    to_unsigned(2147264536,32),
    to_unsigned(2147267467,32),
    to_unsigned(2147270378,32),
    to_unsigned(2147273270,32),
    to_unsigned(2147276142,32),
    to_unsigned(2147278994,32),
    to_unsigned(2147281827,32),
    to_unsigned(2147284639,32),
    to_unsigned(2147287432,32),
    to_unsigned(2147290206,32),
    to_unsigned(2147292959,32),
    to_unsigned(2147295693,32),
    to_unsigned(2147298407,32),
    to_unsigned(2147301101,32),
    to_unsigned(2147303776,32),
    to_unsigned(2147306431,32),
    to_unsigned(2147309066,32),
    to_unsigned(2147311681,32),
    to_unsigned(2147314277,32),
    to_unsigned(2147316853,32),
    to_unsigned(2147319409,32),
    to_unsigned(2147321945,32),
    to_unsigned(2147324462,32),
    to_unsigned(2147326959,32),
    to_unsigned(2147329436,32),
    to_unsigned(2147331894,32),
    to_unsigned(2147334331,32),
    to_unsigned(2147336749,32),
    to_unsigned(2147339148,32),
    to_unsigned(2147341526,32),
    to_unsigned(2147343885,32),
    to_unsigned(2147346224,32),
    to_unsigned(2147348543,32),
    to_unsigned(2147350843,32),
    to_unsigned(2147353123,32),
    to_unsigned(2147355383,32),
    to_unsigned(2147357623,32),
    to_unsigned(2147359844,32),
    to_unsigned(2147362045,32),
    to_unsigned(2147364226,32),
    to_unsigned(2147366387,32),
    to_unsigned(2147368529,32),
    to_unsigned(2147370651,32),
    to_unsigned(2147372753,32),
    to_unsigned(2147374836,32),
    to_unsigned(2147376898,32),
    to_unsigned(2147378941,32),
    to_unsigned(2147380964,32),
    to_unsigned(2147382968,32),
    to_unsigned(2147384952,32),
    to_unsigned(2147386916,32),
    to_unsigned(2147388860,32),
    to_unsigned(2147390785,32),
    to_unsigned(2147392689,32),
    to_unsigned(2147394574,32),
    to_unsigned(2147396440,32),
    to_unsigned(2147398285,32),
    to_unsigned(2147400111,32),
    to_unsigned(2147401917,32),
    to_unsigned(2147403704,32),
    to_unsigned(2147405470,32),
    to_unsigned(2147407217,32),
    to_unsigned(2147408944,32),
    to_unsigned(2147410652,32),
    to_unsigned(2147412340,32),
    to_unsigned(2147414007,32),
    to_unsigned(2147415656,32),
    to_unsigned(2147417284,32),
    to_unsigned(2147418893,32),
    to_unsigned(2147420482,32),
    to_unsigned(2147422051,32),
    to_unsigned(2147423601,32),
    to_unsigned(2147425130,32),
    to_unsigned(2147426640,32),
    to_unsigned(2147428131,32),
    to_unsigned(2147429601,32),
    to_unsigned(2147431052,32),
    to_unsigned(2147432483,32),
    to_unsigned(2147433895,32),
    to_unsigned(2147435286,32),
    to_unsigned(2147436658,32),
    to_unsigned(2147438010,32),
    to_unsigned(2147439342,32),
    to_unsigned(2147440655,32),
    to_unsigned(2147441948,32),
    to_unsigned(2147443221,32),
    to_unsigned(2147444475,32),
    to_unsigned(2147445708,32),
    to_unsigned(2147446922,32),
    to_unsigned(2147448117,32),
    to_unsigned(2147449291,32),
    to_unsigned(2147450446,32),
    to_unsigned(2147451581,32),
    to_unsigned(2147452696,32),
    to_unsigned(2147453792,32),
    to_unsigned(2147454867,32),
    to_unsigned(2147455923,32),
    to_unsigned(2147456960,32),
    to_unsigned(2147457976,32),
    to_unsigned(2147458973,32),
    to_unsigned(2147459950,32),
    to_unsigned(2147460907,32),
    to_unsigned(2147461845,32),
    to_unsigned(2147462763,32),
    to_unsigned(2147463661,32),
    to_unsigned(2147464539,32),
    to_unsigned(2147465398,32),
    to_unsigned(2147466237,32),
    to_unsigned(2147467056,32),
    to_unsigned(2147467856,32),
    to_unsigned(2147468635,32),
    to_unsigned(2147469395,32),
    to_unsigned(2147470136,32),
    to_unsigned(2147470856,32),
    to_unsigned(2147471557,32),
    to_unsigned(2147472238,32),
    to_unsigned(2147472899,32),
    to_unsigned(2147473541,32),
    to_unsigned(2147474162,32),
    to_unsigned(2147474764,32),
    to_unsigned(2147475347,32),
    to_unsigned(2147475909,32),
    to_unsigned(2147476452,32),
    to_unsigned(2147476975,32),
    to_unsigned(2147477479,32),
    to_unsigned(2147477962,32),
    to_unsigned(2147478426,32),
    to_unsigned(2147478870,32),
    to_unsigned(2147479295,32),
    to_unsigned(2147479699,32),
    to_unsigned(2147480084,32),
    to_unsigned(2147480449,32),
    to_unsigned(2147480795,32),
    to_unsigned(2147481120,32),
    to_unsigned(2147481426,32),
    to_unsigned(2147481713,32),
    to_unsigned(2147481979,32),
    to_unsigned(2147482226,32),
    to_unsigned(2147482453,32),
    to_unsigned(2147482660,32),
    to_unsigned(2147482848,32),
    to_unsigned(2147483015,32),
    to_unsigned(2147483163,32),
    to_unsigned(2147483292,32),
    to_unsigned(2147483400,32),
    to_unsigned(2147483489,32),
    to_unsigned(2147483558,32),
    to_unsigned(2147483608,32),
    to_unsigned(2147483608,32)
	);

end dds_sine_pack;

package body dds_sine_pack is
end dds_sine_pack;


-------------------------------------------------------------------------------
-- Digital Quadrature (2-phase) sine/cosine oscillator
-------------------------------------------------------------------------------
--
-- Author: John Clayton
-- Update: Jan.  3, 2014 Wrote code and description.  Tested in simulation,
--                       saw that there is amplitude creep, either growth
--                       or shrinkage over time.  Applied rounding to
--                       mitigate this, with no satisfaction.  Ended up
--                       using an "amplitude reset" technique mentioned in
--                       the book "Digital Signal Processing in VLSI."
--                       The inspiration for this module came from that
--                       book.
--
-- Description
-------------------------------------------------------------------------------
-- This is a discrete time, discrete amplitude binary recursion oscillator.
--
-- The sine and cosine outputs represent the projections of a rotating vector,
-- or complex phasor if you like, along the real and imaginary axes of a
-- 2-dimensional Cartesian coordinate space.  The vector is rotated a fixed
-- amount with each new sample.  Is this just as clear as mud?
--
-- Well, it does take some multipliers to implement the rotation matrix, but
-- otherwise, it's a fairly quick implementation...
--
-- The number of samples per cycle is given as a generic quantity, and the
-- initial values for the vector are zero for sin_o, and +1 for cos_o.
--
-- The numerical quantities are represented as signed 2's complement numbers,
-- in Q1.(AMPL_BITS-1) notation.
--
-- The frequency of the oscillator has been fixed at the lowest possible value.
-- The intention is that by varying the sample rate, sine and cosine waves of
-- different frequencies can be produced.
--
-- For example, if the system clock is at 50 MHz, and SAMPLES_PER_CYCLE=1000,
-- then it should be possible to create output at 50 kHz by setting the
-- clk_en_i input to '1'.  For lower frequencies, just provide a stream of
-- clock enable pulses at the appropriate rate.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library work;
use work.convert_pack.all;

entity quadrature_oscillator is
  generic(
    AMPL_BITS         : natural := 16;
    AMPL_VALUE        : natural := 31768; -- Set to some value below full scale.  There is no saturation!

    SAMPLES_PER_CYCLE : natural := 5000
  );
  port(
    clk_i     : in  std_logic; -- System clock
    rst_n_i   : in  std_logic; -- Low asserted reset
    clk_en_i  : in  std_logic; -- clock enable, determines sample rate

    -- Sine and Cosine outputs
    sin_o     : out signed(AMPL_BITS-1 downto 0);
    cos_o     : out signed(AMPL_BITS-1 downto 0)
  );
end quadrature_oscillator;

architecture beh of quadrature_oscillator is

-- Constants
constant alpha     : real := MATH_2_PI/real(SAMPLES_PER_CYCLE);
constant CA        : real := COS(alpha);
constant SA        : real := SIN(alpha);
constant FULLSCALE : real := 2.0**real(AMPL_BITS-1);
constant ROUNDVAL  : integer := integer(FULLSCALE);
constant C_INT     : integer := integer(CA * FULLSCALE);
constant S_INT     : integer := integer(SA * FULLSCALE);
constant C_VECT : signed(AMPL_BITS-1 downto 0) := to_signed(C_INT,AMPL_BITS);
constant S_VECT : signed(AMPL_BITS-1 downto 0) := to_signed(S_INT,AMPL_BITS);

-- Signals
signal sine     : signed(AMPL_BITS-1 downto 0);
signal cosine   : signed(AMPL_BITS-1 downto 0);
signal s_sop    : signed(2*AMPL_BITS-1 downto 0);
signal c_sop    : signed(2*AMPL_BITS-1 downto 0);
signal s_rnd    : signed(2*AMPL_BITS-1 downto 0);
signal c_rnd    : signed(2*AMPL_BITS-1 downto 0);
signal last_sine_sign : std_logic;

begin

  -- Calculate the sum of products, which is a vector twice as long, with two adjacent sign bits
  s_sop <= S_VECT*cosine + C_VECT*sine;
  c_sop <= C_VECT*cosine - S_VECT*sine;
  -- Get rid of the duplicated sign bit
  -- These signals were named "_rnd" because rounding was tried here...
  -- Alas, although the rounding itself seemed to work, the amplitude decayed anyway.
  -- So, I pulled out the rounding, but kept the names.
  -- To implement rounding, add ROUNDVAL to these.
  s_rnd <= (s_sop(2*AMPL_BITS-2 downto 0) & '0');
  c_rnd <= (c_sop(2*AMPL_BITS-2 downto 0) & '0');

  process (clk_i, rst_n_i)
  begin
    if (rst_n_i = '0') then
      sine   <= (others=>'0');
      last_sine_sign <= '0';
      cosine <= to_signed(AMPL_VALUE,cosine'length);
    elsif (clk_i'event and clk_i = '1') then
      if (clk_en_i = '1') then
        sine   <= s_rnd(2*AMPL_BITS-1 downto AMPL_BITS); -- select the upper half
        cosine <= c_rnd(2*AMPL_BITS-1 downto AMPL_BITS); -- select the upper half
      end if;
      -- Prevent amplitude creep by resetting the cosine component at the
      -- positive zero crossing of the sine signal.
      if s_rnd(2*AMPL_BITS-1)='0' and sine(sine'length-1)='1' then
        cosine <= to_signed(AMPL_VALUE,cosine'length);
      end if;

    end if;
  end process;

sin_o <= sine;
cos_o <= cosine;

end beh;

-------------------------------------------------------------------------------
-- Sinewave Generator Direct Digital Synthesizer (DDS) method
-------------------------------------------------------------------------------
--
-- Author: John Clayton
-- Update: Oct. 15, 2013 Copied code from dds_sine to make this module.
--
-- Description
-------------------------------------------------------------------------------
-- This is a direct digital synthesizer module, which uses a 1/4 wave lookup
-- to produce sinewave samples.  This module is the same as "dds_sine" except
-- that this module uses an internal lookup table instead of an external one.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.convert_pack.all;
use work.dds_sine_pack.all;

entity sine_generator_dds is
  generic(
    PHI_BITS     : natural := 24; -- Bits in phase accumulator, must be >= PHASE_BITS
    AMPL_BITS    : natural := 16;
    PHASE_BITS   : natural := 10
  );
  port(
    clk_i     : in  std_logic;
    rst_n_i   : in  std_logic;
    clk_en_i  : in  std_logic;

    -- Frequency Tuning Word input
    ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

    -- Outputs
    accum_o   : out unsigned(PHI_BITS-1 downto 0);
    sine_o    : out signed(AMPL_BITS-1 downto 0)
    );
end sine_generator_dds;

architecture beh of sine_generator_dds is

  -- Constants
  constant Q_PHASE_BITS     : integer := PHASE_BITS-2;  -- Quarter phase takes two bits less to represent
  constant Q_PHASE_LUT_BITS : integer := PHASE_BITS-2;  -- Quarter phase takes two bits less to represent

  -- Signals
  signal accum        : unsigned(PHI_BITS-1 downto 0);
  signal lut_val      : unsigned(AMPL_BITS-1 downto 0);
  signal lut_val_neg  : unsigned(AMPL_BITS-1 downto 0);
  signal q_phase      : unsigned(Q_PHASE_BITS-1 downto 0);
  signal q_phase_neg  : unsigned(Q_PHASE_BITS-1 downto 0);
  signal phase_value  : unsigned(Q_PHASE_BITS-1 downto 0);
  signal lut_adr      : unsigned(Q_PHASE_LUT_BITS-1 downto 0);

begin

  q_phase      <= u_resize(u_resize_l(accum,PHASE_BITS),q_phase'length); -- Discard the fractional portion
  q_phase_neg  <= (not q_phase)+1;

  process (clk_i, rst_n_i)
  begin
    if (rst_n_i = '0') then
      accum <= (others=>'0');
    elsif (clk_i'event and clk_i = '1') then
      if (clk_en_i = '1') then
        accum  <= accum + ftw_i;
      end if;
    end if;
  end process;

  phase_value  <= q_phase when accum(accum'length-2)='0' else q_phase_neg;
  lut_adr      <= u_resize_l(phase_value,lut_adr'length);
  lut_val      <= u_resize_l(sine_lut_65536_x_32(to_integer(lut_adr)),lut_val'length);
  lut_val_neg  <= (not lut_val) + 1;
  sine_o       <= signed(lut_val) when accum(accum'length-1)='0' else signed(lut_val_neg);
  accum_o      <= accum;

end beh;


-------------------------------------------------------------------------------
-- Direct Digital Synthesizer Power of 2 Length Sinewave Look Up Table module
-------------------------------------------------------------------------------
--
-- Author: John Clayton
-- Update: Sep.  5, 2013 Copied code from dds_sine_non_power_of_two to make
--                       this module.
--
-- Description
-------------------------------------------------------------------------------
-- This is a direct digital synthesizer module, which uses a 1/4 wave lookup
-- to produce sinewave samples.  An external look up table provides the
-- sinewave samples to be used.  The lookup table must be 2**(PHASE_BITS-2)
-- entries long.
--
-- An address bus is provided for indexing into the look up table, and the
-- response data is input via the lut_dat_i bus.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.convert_pack.all;

entity dds_sine is
  generic(
    PHI_BITS     : natural := 24; -- Bits in phase accumulator, must be >= PHASE_BITS
    AMPL_BITS    : natural := 16;
    PHASE_BITS   : natural := 10
  );
  port(
    clk_i     : in  std_logic;
    rst_n_i   : in  std_logic;
    clk_en_i  : in  std_logic;

    -- Look Up Table interface
    lut_adr_o : out unsigned(PHASE_BITS-3 downto 0); -- Quarter wave LUT
    lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

    -- Frequency Tuning Word input
    ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

    -- Outputs
    accum_o   : out unsigned(PHI_BITS-1 downto 0);
    sine_o    : out signed(AMPL_BITS-1 downto 0)
    );
end dds_sine;

architecture beh of dds_sine is

  -- Constants
  constant Q_PHASE_BITS : integer := PHASE_BITS-2;  -- Quarter phase takes two bits less to represent

  -- Signals
  signal accum        : unsigned(PHI_BITS-1 downto 0);
  signal lut_out      : unsigned(AMPL_BITS-1 downto 0);
  signal lut_out_neg  : unsigned(AMPL_BITS-1 downto 0);
  signal q_phase      : unsigned(Q_PHASE_BITS-1 downto 0);
  signal q_phase_neg  : unsigned(Q_PHASE_BITS-1 downto 0);

begin

  q_phase      <= u_resize(u_resize_l(accum,PHASE_BITS),q_phase'length); -- Discard the fractional portion
  q_phase_neg  <= (not q_phase)+1;

  process (clk_i, rst_n_i)
  begin
    if (rst_n_i = '0') then
      accum <= (others=>'0');
    elsif (clk_i'event and clk_i = '1') then
      if (clk_en_i = '1') then
        accum  <= accum + ftw_i;
      end if;
    end if;
  end process;

  lut_adr_o    <= q_phase when accum(accum'length-2)='0' else q_phase_neg;
  lut_out      <= lut_dat_i;
  lut_out_neg  <= (not lut_out) + 1;
  sine_o       <= signed(lut_out) when accum(accum'length-1)='0' else signed(lut_out_neg);
  accum_o      <= accum;

end beh;


-------------------------------------------------------------------------------
-- Direct Digital Synthesizer Arbitrary Length Sinewave Look Up Table module
-------------------------------------------------------------------------------
--
-- Author: John Clayton
-- Update: Jan. 24, 2013 Modified Matlab script "sine_arbitrary_length_lut_gen"
--                       to produce VHDL output which uses the "unsigned" type
--                       from ieee.numeric_std library.
--         Jan. 26, 2013 Rewrote accumulator folding logic.  Added saturation
--                       check to avoid indices beyond the end of the lookup
--                       table.
--         Sep.  5, 2013 Restructured the module to use external look up
--                       tables.  Created generics for AMPL_BITS, PHASE_LENGTH
--                       and PHASE_BITS.
--
-- Description
-------------------------------------------------------------------------------
-- This is a direct digital synthesizer module, which uses a 1/4 wave lookup
-- to produce waveform samples.  An external look up table provides the
-- sinewave samples to be used.  The lookup table can be any length, being
-- one quarter of PHASE_LENGTH entries long.
--
-- An address bus is provided for indexing into the look up table, and the
-- response data is input via the lut_dat_i bus.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.convert_pack.all;

entity dds_sine_non_power_of_two is
  generic(
    PHI_BITS     : natural := 24; -- Bits in phase accumulator, must be >= PHASE_BITS
    AMPL_BITS    : natural := 16;
    PHASE_LENGTH : natural := 1024;
    PHASE_BITS   : natural := 10
  );
  port(
    clk_i     : in  std_logic;
    rst_n_i   : in  std_logic;
    clk_en_i  : in  std_logic;

    -- Look Up Table interface
    lut_adr_o : out unsigned(PHASE_BITS-3 downto 0); -- Quarter wave LUT
    lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

    -- Frequency Tuning Word input
    ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

    -- Outputs
    accum_o   : out unsigned(PHI_BITS-1 downto 0);
    sine_o    : out signed(AMPL_BITS-1 downto 0)
    );
end dds_sine_non_power_of_two;

architecture beh of dds_sine_non_power_of_two is

  constant FRAC_BITS    : natural := PHI_BITS - PHASE_BITS;
  constant Q_PHASE_BITS : integer := PHASE_BITS-2;  -- Quarter phase takes two bits less to represent
  constant Q_LENGTH     : unsigned(Q_PHASE_BITS-1 downto 0) := to_unsigned(PHASE_LENGTH/4,Q_PHASE_BITS); -- Quadrant Length
  constant Q_THRESH     : unsigned(PHI_BITS-1 downto 0) := to_unsigned(2**FRAC_BITS*PHASE_LENGTH/4,PHI_BITS); -- Quadrant Length

  signal accum        : unsigned(PHI_BITS-1 downto 0);
  signal q_accum      : unsigned(PHI_BITS-1 downto 0);
  signal q_accum_next : unsigned(PHI_BITS-1 downto 0);
  signal accum_incr   : unsigned(PHI_BITS-1 downto 0);
  signal accum_folded : unsigned(PHI_BITS-1 downto 0);
  signal lut_out      : unsigned(AMPL_BITS-1 downto 0);
  signal lut_out_neg  : unsigned(AMPL_BITS-1 downto 0);

  signal q_phase      : unsigned(Q_PHASE_BITS-1 downto 0);
  signal q_phase_sat  : unsigned(Q_PHASE_BITS-1 downto 0);
  signal q_count      : unsigned(1 downto 0);
  signal q_count_r1   : unsigned(1 downto 0);

begin

  accum_incr   <= unsigned(ftw_i);
  q_accum_next   <= q_accum + accum_incr;
  accum_folded <=            q_accum when q_count(0)='0' else
                  Q_THRESH - q_accum;
  q_phase      <= u_resize(u_resize_l(accum_folded,PHASE_BITS),q_phase'length); -- Discard the fractional portion

  process (clk_i, rst_n_i)
  begin
    if (rst_n_i = '0') then
      accum       <= (others=>'0');
      q_accum     <= (others=>'0');
      q_count     <= (others=>'0');
      q_count_r1  <= (others=>'0');
      q_phase_sat <= (others=>'0');
    elsif (clk_i'event and clk_i = '1') then
      if (clk_en_i = '1') then
        if (q_accum_next > Q_THRESH) then
          q_accum <= q_accum_next - Q_THRESH;
          q_count <= q_count+1;
          if (q_count="11") then
            accum <= (others=>'0');
          else
            accum   <= accum + Q_THRESH;
          end if;
        else
          q_accum <= q_accum_next;
        end if;

        -- Delayed q_count, to match delayed q_phase
        q_count_r1 <= q_count;
        -- Saturate the quarter phase signal, to avoid overflows when looking up sine values
        if (q_phase>=(PHASE_LENGTH/4)) then
          q_phase_sat <= to_unsigned(PHASE_LENGTH/4-1,q_phase_sat'length);
        else
          q_phase_sat <= q_phase;
        end if;
      end if;
    end if;
  end process;

  lut_adr_o    <= q_phase_sat;
  lut_out      <= lut_dat_i;
  lut_out_neg  <= (not lut_out) + 1;
  sine_o       <= signed(lut_out_neg) when q_count_r1(1) = '1' else signed(lut_out);
  accum_o      <= accum+q_accum;

end beh;

-------------------------------------------------------------------------------
-- Direct Digital Synthesizer Arbitrary Waveform Look Up Table module
-------------------------------------------------------------------------------
--
-- Author: John Clayton
-- Update: Sep.  5, 2013 Copied code from dds_sine to make this module.
--
-- Description
-------------------------------------------------------------------------------
-- This is a direct digital synthesizer module, which uses a full wave lookup
-- to produce waveform samples.  The lookup table is external.
-- The lookup table must be 2**PHASE_BITS entries long.
--
-- An address bus is provided for indexing into the look up table, and the
-- response data is input via the lut_dat_i bus.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.convert_pack.all;

entity dds_arb is
  generic(
    PHI_BITS     : natural := 24; -- Bits in phase accumulator, must be >= PHASE_BITS
    AMPL_BITS    : natural := 16;
    PHASE_BITS   : natural := 10
  );
  port(
    clk_i     : in  std_logic;
    rst_n_i   : in  std_logic;
    clk_en_i  : in  std_logic;

    -- Look Up Table interface
    lut_adr_o : out unsigned(PHASE_BITS-1 downto 0); -- Full wave LUT
    lut_dat_i : in  unsigned(AMPL_BITS-1 downto 0);

    -- Frequency Tuning Word input
    ftw_i     : in  unsigned(PHI_BITS-1 downto 0);

    -- Outputs
    accum_o   : out unsigned(PHI_BITS-1 downto 0);
    arb_o     : out signed(AMPL_BITS-1 downto 0)
    );
end dds_arb;

architecture beh of dds_arb is

  -- Constants
  constant Q_PHASE_BITS : integer := PHASE_BITS-2;  -- Quarter phase takes two bits less to represent

  -- Signals
  signal accum        : unsigned(PHI_BITS-1 downto 0);

begin

  process (clk_i, rst_n_i)
  begin
    if (rst_n_i = '0') then
      accum <= (others=>'0');
    elsif (clk_i'event and clk_i = '1') then
      if (clk_en_i = '1') then
        accum   <= accum + ftw_i;
      end if;
    end if;
  end process;

  lut_adr_o <= u_resize_l(accum,PHASE_BITS); -- Discard the fractional portion
  accum_o   <= accum;
  arb_o     <= signed(lut_dat_i);

end beh;

