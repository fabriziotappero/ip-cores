-- DAC_AHB enable 
  constant CFG_DAC_AHB  : integer := CONFIG_DAC_AHB_ENABLE;

