----------------------------------------------------------------------------------
-- Company		: OCST Co.,Ltd.
-- Engineer		: RyuShinHyung
-- 
-- Create Date	: 02/23/2005
-- Design Name	: 
-- Module Name	: ENC8B10B - RTL
-- Project Name	: Fiber Optic Application
--
-- Revision
-- Revision 0.01 - File Created.
--          1.00 - publishing on the opencores.org.
--          1.01 - eliminate needing the VECTLIB.vhd in the original revision.(20110424)
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ENC8B10B is
	port
	(
		CLK_IN : in STD_LOGIC;
		RUNDP_RESET_IN : in STD_LOGIC;
		CTRL_IN : in STD_LOGIC;
		DATA_IN : in STD_LOGIC_VECTOR(7 downto 0);
		RUNDP_OUT : out STD_LOGIC;
		ENCODE_OUT : out STD_LOGIC_VECTOR(9 downto 0)
	);
end ENC8B10B;

architecture RTL of ENC8B10B is

type TYPE_ENC8b10b is array (0 to 1023) of std_logic_vector (10 downto 0); -- RD & Dx.y
signal TBL_ENC8b10b : TYPE_ENC8b10b:=
	(
	--	"Rjhgfiedcba"	-- RD(Pre) + Dx.y => RD(Post)
		"00010111001",	-- "00000000" -D00.0- [0]
		"00010101110",	-- "00000001" -D01.0- [1]
		"00010101101",	-- "00000010" -D02.0- [2]
		"11101100011",	-- "00000011" -D03.0+ [3]
		"00010101011",	-- "00000100" -D04.0- [4]
		"11101100101",	-- "00000101" -D05.0+ [5]
		"11101100110",	-- "00000110" -D06.0+ [6]
		"11101000111",	-- "00000111" -D07.0+ [7]
		"00010100111",	-- "00001000" -D08.0- [8]
		"11101101001",	-- "00001001" -D09.0+ [9]
		"11101101010",	-- "00001010" -D10.0+ [10]
		"11101001011",	-- "00001011" -D11.0+ [11]
		"11101101100",	-- "00001100" -D12.0+ [12]
		"11101001101",	-- "00001101" -D13.0+ [13]
		"11101001110",	-- "00001110" -D14.0+ [14]
		"00010111010",	-- "00001111" -D15.0- [15]
		"00010110110",	-- "00010000" -D16.0- [16]
		"11101110001",	-- "00010001" -D17.0+ [17]
		"11101110010",	-- "00010010" -D18.0+ [18]
		"11101010011",	-- "00010011" -D19.0+ [19]
		"11101110100",	-- "00010100" -D20.0+ [20]
		"11101010101",	-- "00010101" -D21.0+ [21]
		"11101010110",	-- "00010110" -D22.0+ [22]
		"00010010111",	-- "00010111" -D23.0- [23]
		"00010110011",	-- "00011000" -D24.0- [24]
		"11101011001",	-- "00011001" -D25.0+ [25]
		"11101011010",	-- "00011010" -D26.0+ [26]
		"00010011011",	-- "00011011" -D27.0- [27]
		"11101011100",	-- "00011100" -D28.0+ [28]
		"00010011101",	-- "00011101" -D29.0- [29]
		"00010011110",	-- "00011110" -D30.0- [30]
		"00010110101",	-- "00011111" -D31.0- [31]
		"11001111001",	-- "00100000" -D00.1+ [32]
		"11001101110",	-- "00100001" -D01.1+ [33]
		"11001101101",	-- "00100010" -D02.1+ [34]
		"01001100011",	-- "00100011" -D03.1- [35]
		"11001101011",	-- "00100100" -D04.1+ [36]
		"01001100101",	-- "00100101" -D05.1- [37]
		"01001100110",	-- "00100110" -D06.1- [38]
		"01001000111",	-- "00100111" -D07.1- [39]
		"11001100111",	-- "00101000" -D08.1+ [40]
		"01001101001",	-- "00101001" -D09.1- [41]
		"01001101010",	-- "00101010" -D10.1- [42]
		"01001001011",	-- "00101011" -D11.1- [43]
		"01001101100",	-- "00101100" -D12.1- [44]
		"01001001101",	-- "00101101" -D13.1- [45]
		"01001001110",	-- "00101110" -D14.1- [46]
		"11001111010",	-- "00101111" -D15.1+ [47]
		"11001110110",	-- "00110000" -D16.1+ [48]
		"01001110001",	-- "00110001" -D17.1- [49]
		"01001110010",	-- "00110010" -D18.1- [50]
		"01001010011",	-- "00110011" -D19.1- [51]
		"01001110100",	-- "00110100" -D20.1- [52]
		"01001010101",	-- "00110101" -D21.1- [53]
		"01001010110",	-- "00110110" -D22.1- [54]
		"11001010111",	-- "00110111" -D23.1+ [55]
		"11001110011",	-- "00111000" -D24.1+ [56]
		"01001011001",	-- "00111001" -D25.1- [57]
		"01001011010",	-- "00111010" -D26.1- [58]
		"11001011011",	-- "00111011" -D27.1+ [59]
		"01001011100",	-- "00111100" -D28.1- [60]
		"11001011101",	-- "00111101" -D29.1+ [61]
		"11001011110",	-- "00111110" -D30.1+ [62]
		"11001110101",	-- "00111111" -D31.1+ [63]
		"11010111001",	-- "01000000" -D00.2+ [64]
		"11010101110",	-- "01000001" -D01.2+ [65]
		"11010101101",	-- "01000010" -D02.2+ [66]
		"01010100011",	-- "01000011" -D03.2- [67]
		"11010101011",	-- "01000100" -D04.2+ [68]
		"01010100101",	-- "01000101" -D05.2- [69]
		"01010100110",	-- "01000110" -D06.2- [70]
		"01010000111",	-- "01000111" -D07.2- [71]
		"11010100111",	-- "01001000" -D08.2+ [72]
		"01010101001",	-- "01001001" -D09.2- [73]
		"01010101010",	-- "01001010" -D10.2- [74]
		"01010001011",	-- "01001011" -D11.2- [75]
		"01010101100",	-- "01001100" -D12.2- [76]
		"01010001101",	-- "01001101" -D13.2- [77]
		"01010001110",	-- "01001110" -D14.2- [78]
		"11010111010",	-- "01001111" -D15.2+ [79]
		"11010110110",	-- "01010000" -D16.2+ [80]
		"01010110001",	-- "01010001" -D17.2- [81]
		"01010110010",	-- "01010010" -D18.2- [82]
		"01010010011",	-- "01010011" -D19.2- [83]
		"01010110100",	-- "01010100" -D20.2- [84]
		"01010010101",	-- "01010101" -D21.2- [85]
		"01010010110",	-- "01010110" -D22.2- [86]
		"11010010111",	-- "01010111" -D23.2+ [87]
		"11010110011",	-- "01011000" -D24.2+ [88]
		"01010011001",	-- "01011001" -D25.2- [89]
		"01010011010",	-- "01011010" -D26.2- [90]
		"11010011011",	-- "01011011" -D27.2+ [91]
		"01010011100",	-- "01011100" -D28.2- [92]
		"11010011101",	-- "01011101" -D29.2+ [93]
		"11010011110",	-- "01011110" -D30.2+ [94]
		"11010110101",	-- "01011111" -D31.2+ [95]
		"11100111001",	-- "01100000" -D00.3+ [96]
		"11100101110",	-- "01100001" -D01.3+ [97]
		"11100101101",	-- "01100010" -D02.3+ [98]
		"00011100011",	-- "01100011" -D03.3- [99]
		"11100101011",	-- "01100100" -D04.3+ [100]
		"00011100101",	-- "01100101" -D05.3- [101]
		"00011100110",	-- "01100110" -D06.3- [102]
		"00011000111",	-- "01100111" -D07.3- [103]
		"11100100111",	-- "01101000" -D08.3+ [104]
		"00011101001",	-- "01101001" -D09.3- [105]
		"00011101010",	-- "01101010" -D10.3- [106]
		"00011001011",	-- "01101011" -D11.3- [107]
		"00011101100",	-- "01101100" -D12.3- [108]
		"00011001101",	-- "01101101" -D13.3- [109]
		"00011001110",	-- "01101110" -D14.3- [110]
		"11100111010",	-- "01101111" -D15.3+ [111]
		"11100110110",	-- "01110000" -D16.3+ [112]
		"00011110001",	-- "01110001" -D17.3- [113]
		"00011110010",	-- "01110010" -D18.3- [114]
		"00011010011",	-- "01110011" -D19.3- [115]
		"00011110100",	-- "01110100" -D20.3- [116]
		"00011010101",	-- "01110101" -D21.3- [117]
		"00011010110",	-- "01110110" -D22.3- [118]
		"11100010111",	-- "01110111" -D23.3+ [119]
		"11100110011",	-- "01111000" -D24.3+ [120]
		"00011011001",	-- "01111001" -D25.3- [121]
		"00011011010",	-- "01111010" -D26.3- [122]
		"11100011011",	-- "01111011" -D27.3+ [123]
		"00011011100",	-- "01111100" -D28.3- [124]
		"11100011101",	-- "01111101" -D29.3+ [125]
		"11100011110",	-- "01111110" -D30.3+ [126]
		"11100110101",	-- "01111111" -D31.3+ [127]
		"00100111001",	-- "10000000" -D00.4- [128]
		"00100101110",	-- "10000001" -D01.4- [129]
		"00100101101",	-- "10000010" -D02.4- [130]
		"11011100011",	-- "10000011" -D03.4+ [131]
		"00100101011",	-- "10000100" -D04.4- [132]
		"11011100101",	-- "10000101" -D05.4+ [133]
		"11011100110",	-- "10000110" -D06.4+ [134]
		"11011000111",	-- "10000111" -D07.4+ [135]
		"00100100111",	-- "10001000" -D08.4- [136]
		"11011101001",	-- "10001001" -D09.4+ [137]
		"11011101010",	-- "10001010" -D10.4+ [138]
		"11011001011",	-- "10001011" -D11.4+ [139]
		"11011101100",	-- "10001100" -D12.4+ [140]
		"11011001101",	-- "10001101" -D13.4+ [141]
		"11011001110",	-- "10001110" -D14.4+ [142]
		"00100111010",	-- "10001111" -D15.4- [143]
		"00100110110",	-- "10010000" -D16.4- [144]
		"11011110001",	-- "10010001" -D17.4+ [145]
		"11011110010",	-- "10010010" -D18.4+ [146]
		"11011010011",	-- "10010011" -D19.4+ [147]
		"11011110100",	-- "10010100" -D20.4+ [148]
		"11011010101",	-- "10010101" -D21.4+ [149]
		"11011010110",	-- "10010110" -D22.4+ [150]
		"00100010111",	-- "10010111" -D23.4- [151]
		"00100110011",	-- "10011000" -D24.4- [152]
		"11011011001",	-- "10011001" -D25.4+ [153]
		"11011011010",	-- "10011010" -D26.4+ [154]
		"00100011011",	-- "10011011" -D27.4- [155]
		"11011011100",	-- "10011100" -D28.4+ [156]
		"00100011101",	-- "10011101" -D29.4- [157]
		"00100011110",	-- "10011110" -D30.4- [158]
		"00100110101",	-- "10011111" -D31.4- [159]
		"10101111001",	-- "10100000" -D00.5+ [160]
		"10101101110",	-- "10100001" -D01.5+ [161]
		"10101101101",	-- "10100010" -D02.5+ [162]
		"00101100011",	-- "10100011" -D03.5- [163]
		"10101101011",	-- "10100100" -D04.5+ [164]
		"00101100101",	-- "10100101" -D05.5- [165]
		"00101100110",	-- "10100110" -D06.5- [166]
		"00101000111",	-- "10100111" -D07.5- [167]
		"10101100111",	-- "10101000" -D08.5+ [168]
		"00101101001",	-- "10101001" -D09.5- [169]
		"00101101010",	-- "10101010" -D10.5- [170]
		"00101001011",	-- "10101011" -D11.5- [171]
		"00101101100",	-- "10101100" -D12.5- [172]
		"00101001101",	-- "10101101" -D13.5- [173]
		"00101001110",	-- "10101110" -D14.5- [174]
		"10101111010",	-- "10101111" -D15.5+ [175]
		"10101110110",	-- "10110000" -D16.5+ [176]
		"00101110001",	-- "10110001" -D17.5- [177]
		"00101110010",	-- "10110010" -D18.5- [178]
		"00101010011",	-- "10110011" -D19.5- [179]
		"00101110100",	-- "10110100" -D20.5- [180]
		"00101010101",	-- "10110101" -D21.5- [181]
		"00101010110",	-- "10110110" -D22.5- [182]
		"10101010111",	-- "10110111" -D23.5+ [183]
		"10101110011",	-- "10111000" -D24.5+ [184]
		"00101011001",	-- "10111001" -D25.5- [185]
		"00101011010",	-- "10111010" -D26.5- [186]
		"10101011011",	-- "10111011" -D27.5+ [187]
		"00101011100",	-- "10111100" -D28.5- [188]
		"10101011101",	-- "10111101" -D29.5+ [189]
		"10101011110",	-- "10111110" -D30.5+ [190]
		"10101110101",	-- "10111111" -D31.5+ [191]
		"10110111001",	-- "11000000" -D00.6+ [192]
		"10110101110",	-- "11000001" -D01.6+ [193]
		"10110101101",	-- "11000010" -D02.6+ [194]
		"00110100011",	-- "11000011" -D03.6- [195]
		"10110101011",	-- "11000100" -D04.6+ [196]
		"00110100101",	-- "11000101" -D05.6- [197]
		"00110100110",	-- "11000110" -D06.6- [198]
		"00110000111",	-- "11000111" -D07.6- [199]
		"10110100111",	-- "11001000" -D08.6+ [200]
		"00110101001",	-- "11001001" -D09.6- [201]
		"00110101010",	-- "11001010" -D10.6- [202]
		"00110001011",	-- "11001011" -D11.6- [203]
		"00110101100",	-- "11001100" -D12.6- [204]
		"00110001101",	-- "11001101" -D13.6- [205]
		"00110001110",	-- "11001110" -D14.6- [206]
		"10110111010",	-- "11001111" -D15.6+ [207]
		"10110110110",	-- "11010000" -D16.6+ [208]
		"00110110001",	-- "11010001" -D17.6- [209]
		"00110110010",	-- "11010010" -D18.6- [210]
		"00110010011",	-- "11010011" -D19.6- [211]
		"00110110100",	-- "11010100" -D20.6- [212]
		"00110010101",	-- "11010101" -D21.6- [213]
		"00110010110",	-- "11010110" -D22.6- [214]
		"10110010111",	-- "11010111" -D23.6+ [215]
		"10110110011",	-- "11011000" -D24.6+ [216]
		"00110011001",	-- "11011001" -D25.6- [217]
		"00110011010",	-- "11011010" -D26.6- [218]
		"10110011011",	-- "11011011" -D27.6+ [219]
		"00110011100",	-- "11011100" -D28.6- [220]
		"10110011101",	-- "11011101" -D29.6+ [221]
		"10110011110",	-- "11011110" -D30.6+ [222]
		"10110110101",	-- "11011111" -D31.6+ [223]
		"01000111001",	-- "11100000" -D00.7- [224]
		"01000101110",	-- "11100001" -D01.7- [225]
		"01000101101",	-- "11100010" -D02.7- [226]
		"10111100011",	-- "11100011" -D03.7+ [227]
		"01000101011",	-- "11100100" -D04.7- [228]
		"10111100101",	-- "11100101" -D05.7+ [229]
		"10111100110",	-- "11100110" -D06.7+ [230]
		"10111000111",	-- "11100111" -D07.7+ [231]
		"01000100111",	-- "11101000" -D08.7- [232]
		"10111101001",	-- "11101001" -D09.7+ [233]
		"10111101010",	-- "11101010" -D10.7+ [234]
		"10111001011",	-- "11101011" -D11.7+ [235]
		"10111101100",	-- "11101100" -D12.7+ [236]
		"10111001101",	-- "11101101" -D13.7+ [237]
		"10111001110",	-- "11101110" -D14.7+ [238]
		"01000111010",	-- "11101111" -D15.7- [239]
		"01000110110",	-- "11110000" -D16.7- [240]
		"11110110001",	-- "11110001" -D17.7+ [241]
		"11110110010",	-- "11110010" -D18.7+ [242]
		"10111010011",	-- "11110011" -D19.7+ [243]
		"11110110100",	-- "11110100" -D20.7+ [244]
		"10111010101",	-- "11110101" -D21.7+ [245]
		"10111010110",	-- "11110110" -D22.7+ [246]
		"01000010111",	-- "11110111" -D23.7- [247]
		"01000110011",	-- "11111000" -D24.7- [248]
		"10111011001",	-- "11111001" -D25.7+ [249]
		"10111011010",	-- "11111010" -D26.7+ [250]
		"01000011011",	-- "11111011" -D27.7- [251]
		"10111011100",	-- "11111100" -D28.7+ [252]
		"01000011101",	-- "11111101" -D29.7- [253]
		"01000011110",	-- "11111110" -D30.7- [254]
		"01000110101",	-- "11111111" -D31.7- [255]
		"11101000110",	-- "00000000" +D00.0+ [256]
		"11101010001",	-- "00000001" +D01.0+ [257]
		"11101010010",	-- "00000010" +D02.0+ [258]
		"00010100011",	-- "00000011" +D03.0- [259]
		"11101010100",	-- "00000100" +D04.0+ [260]
		"00010100101",	-- "00000101" +D05.0- [261]
		"00010100110",	-- "00000110" +D06.0- [262]
		"00010111000",	-- "00000111" +D07.0- [263]
		"11101011000",	-- "00001000" +D08.0+ [264]
		"00010101001",	-- "00001001" +D09.0- [265]
		"00010101010",	-- "00001010" +D10.0- [266]
		"00010001011",	-- "00001011" +D11.0- [267]
		"00010101100",	-- "00001100" +D12.0- [268]
		"00010001101",	-- "00001101" +D13.0- [269]
		"00010001110",	-- "00001110" +D14.0- [270]
		"11101000101",	-- "00001111" +D15.0+ [271]
		"11101001001",	-- "00010000" +D16.0+ [272]
		"00010110001",	-- "00010001" +D17.0- [273]
		"00010110010",	-- "00010010" +D18.0- [274]
		"00010010011",	-- "00010011" +D19.0- [275]
		"00010110100",	-- "00010100" +D20.0- [276]
		"00010010101",	-- "00010101" +D21.0- [277]
		"00010010110",	-- "00010110" +D22.0- [278]
		"11101101000",	-- "00010111" +D23.0+ [279]
		"11101001100",	-- "00011000" +D24.0+ [280]
		"00010011001",	-- "00011001" +D25.0- [281]
		"00010011010",	-- "00011010" +D26.0- [282]
		"11101100100",	-- "00011011" +D27.0+ [283]
		"00010011100",	-- "00011100" +D28.0- [284]
		"11101100010",	-- "00011101" +D29.0+ [285]
		"11101100001",	-- "00011110" +D30.0+ [286]
		"11101001010",	-- "00011111" +D31.0+ [287]
		"01001000110",	-- "00100000" +D00.1- [288]
		"01001010001",	-- "00100001" +D01.1- [289]
		"01001010010",	-- "00100010" +D02.1- [290]
		"11001100011",	-- "00100011" +D03.1+ [291]
		"01001010100",	-- "00100100" +D04.1- [292]
		"11001100101",	-- "00100101" +D05.1+ [293]
		"11001100110",	-- "00100110" +D06.1+ [294]
		"11001111000",	-- "00100111" +D07.1+ [295]
		"01001011000",	-- "00101000" +D08.1- [296]
		"11001101001",	-- "00101001" +D09.1+ [297]
		"11001101010",	-- "00101010" +D10.1+ [298]
		"11001001011",	-- "00101011" +D11.1+ [299]
		"11001101100",	-- "00101100" +D12.1+ [300]
		"11001001101",	-- "00101101" +D13.1+ [301]
		"11001001110",	-- "00101110" +D14.1+ [302]
		"01001000101",	-- "00101111" +D15.1- [303]
		"01001001001",	-- "00110000" +D16.1- [304]
		"11001110001",	-- "00110001" +D17.1+ [305]
		"11001110010",	-- "00110010" +D18.1+ [306]
		"11001010011",	-- "00110011" +D19.1+ [307]
		"11001110100",	-- "00110100" +D20.1+ [308]
		"11001010101",	-- "00110101" +D21.1+ [309]
		"11001010110",	-- "00110110" +D22.1+ [310]
		"01001101000",	-- "00110111" +D23.1- [311]
		"01001001100",	-- "00111000" +D24.1- [312]
		"11001011001",	-- "00111001" +D25.1+ [313]
		"11001011010",	-- "00111010" +D26.1+ [314]
		"01001100100",	-- "00111011" +D27.1- [315]
		"11001011100",	-- "00111100" +D28.1+ [316]
		"01001100010",	-- "00111101" +D29.1- [317]
		"01001100001",	-- "00111110" +D30.1- [318]
		"01001001010",	-- "00111111" +D31.1- [319]
		"01010000110",	-- "01000000" +D00.2- [320]
		"01010010001",	-- "01000001" +D01.2- [321]
		"01010010010",	-- "01000010" +D02.2- [322]
		"11010100011",	-- "01000011" +D03.2+ [323]
		"01010010100",	-- "01000100" +D04.2- [324]
		"11010100101",	-- "01000101" +D05.2+ [325]
		"11010100110",	-- "01000110" +D06.2+ [326]
		"11010111000",	-- "01000111" +D07.2+ [327]
		"01010011000",	-- "01001000" +D08.2- [328]
		"11010101001",	-- "01001001" +D09.2+ [329]
		"11010101010",	-- "01001010" +D10.2+ [330]
		"11010001011",	-- "01001011" +D11.2+ [331]
		"11010101100",	-- "01001100" +D12.2+ [332]
		"11010001101",	-- "01001101" +D13.2+ [333]
		"11010001110",	-- "01001110" +D14.2+ [334]
		"01010000101",	-- "01001111" +D15.2- [335]
		"01010001001",	-- "01010000" +D16.2- [336]
		"11010110001",	-- "01010001" +D17.2+ [337]
		"11010110010",	-- "01010010" +D18.2+ [338]
		"11010010011",	-- "01010011" +D19.2+ [339]
		"11010110100",	-- "01010100" +D20.2+ [340]
		"11010010101",	-- "01010101" +D21.2+ [341]
		"11010010110",	-- "01010110" +D22.2+ [342]
		"01010101000",	-- "01010111" +D23.2- [343]
		"01010001100",	-- "01011000" +D24.2- [344]
		"11010011001",	-- "01011001" +D25.2+ [345]
		"11010011010",	-- "01011010" +D26.2+ [346]
		"01010100100",	-- "01011011" +D27.2- [347]
		"11010011100",	-- "01011100" +D28.2+ [348]
		"01010100010",	-- "01011101" +D29.2- [349]
		"01010100001",	-- "01011110" +D30.2- [350]
		"01010001010",	-- "01011111" +D31.2- [351]
		"00011000110",	-- "01100000" +D00.3- [352]
		"00011010001",	-- "01100001" +D01.3- [353]
		"00011010010",	-- "01100010" +D02.3- [354]
		"11100100011",	-- "01100011" +D03.3+ [355]
		"00011010100",	-- "01100100" +D04.3- [356]
		"11100100101",	-- "01100101" +D05.3+ [357]
		"11100100110",	-- "01100110" +D06.3+ [358]
		"11100111000",	-- "01100111" +D07.3+ [359]
		"00011011000",	-- "01101000" +D08.3- [360]
		"11100101001",	-- "01101001" +D09.3+ [361]
		"11100101010",	-- "01101010" +D10.3+ [362]
		"11100001011",	-- "01101011" +D11.3+ [363]
		"11100101100",	-- "01101100" +D12.3+ [364]
		"11100001101",	-- "01101101" +D13.3+ [365]
		"11100001110",	-- "01101110" +D14.3+ [366]
		"00011000101",	-- "01101111" +D15.3- [367]
		"00011001001",	-- "01110000" +D16.3- [368]
		"11100110001",	-- "01110001" +D17.3+ [369]
		"11100110010",	-- "01110010" +D18.3+ [370]
		"11100010011",	-- "01110011" +D19.3+ [371]
		"11100110100",	-- "01110100" +D20.3+ [372]
		"11100010101",	-- "01110101" +D21.3+ [373]
		"11100010110",	-- "01110110" +D22.3+ [374]
		"00011101000",	-- "01110111" +D23.3- [375]
		"00011001100",	-- "01111000" +D24.3- [376]
		"11100011001",	-- "01111001" +D25.3+ [377]
		"11100011010",	-- "01111010" +D26.3+ [378]
		"00011100100",	-- "01111011" +D27.3- [379]
		"11100011100",	-- "01111100" +D28.3+ [380]
		"00011100010",	-- "01111101" +D29.3- [381]
		"00011100001",	-- "01111110" +D30.3- [382]
		"00011001010",	-- "01111111" +D31.3- [383]
		"11011000110",	-- "10000000" +D00.4+ [384]
		"11011010001",	-- "10000001" +D01.4+ [385]
		"11011010010",	-- "10000010" +D02.4+ [386]
		"00100100011",	-- "10000011" +D03.4- [387]
		"11011010100",	-- "10000100" +D04.4+ [388]
		"00100100101",	-- "10000101" +D05.4- [389]
		"00100100110",	-- "10000110" +D06.4- [390]
		"00100111000",	-- "10000111" +D07.4- [391]
		"11011011000",	-- "10001000" +D08.4+ [392]
		"00100101001",	-- "10001001" +D09.4- [393]
		"00100101010",	-- "10001010" +D10.4- [394]
		"00100001011",	-- "10001011" +D11.4- [395]
		"00100101100",	-- "10001100" +D12.4- [396]
		"00100001101",	-- "10001101" +D13.4- [397]
		"00100001110",	-- "10001110" +D14.4- [398]
		"11011000101",	-- "10001111" +D15.4+ [399]
		"11011001001",	-- "10010000" +D16.4+ [400]
		"00100110001",	-- "10010001" +D17.4- [401]
		"00100110010",	-- "10010010" +D18.4- [402]
		"00100010011",	-- "10010011" +D19.4- [403]
		"00100110100",	-- "10010100" +D20.4- [404]
		"00100010101",	-- "10010101" +D21.4- [405]
		"00100010110",	-- "10010110" +D22.4- [406]
		"11011101000",	-- "10010111" +D23.4+ [407]
		"11011001100",	-- "10011000" +D24.4+ [408]
		"00100011001",	-- "10011001" +D25.4- [409]
		"00100011010",	-- "10011010" +D26.4- [410]
		"11011100100",	-- "10011011" +D27.4+ [411]
		"00100011100",	-- "10011100" +D28.4- [412]
		"11011100010",	-- "10011101" +D29.4+ [413]
		"11011100001",	-- "10011110" +D30.4+ [414]
		"11011001010",	-- "10011111" +D31.4+ [415]
		"00101000110",	-- "10100000" +D00.5- [416]
		"00101010001",	-- "10100001" +D01.5- [417]
		"00101010010",	-- "10100010" +D02.5- [418]
		"10101100011",	-- "10100011" +D03.5+ [419]
		"00101010100",	-- "10100100" +D04.5- [420]
		"10101100101",	-- "10100101" +D05.5+ [421]
		"10101100110",	-- "10100110" +D06.5+ [422]
		"10101111000",	-- "10100111" +D07.5+ [423]
		"00101011000",	-- "10101000" +D08.5- [424]
		"10101101001",	-- "10101001" +D09.5+ [425]
		"10101101010",	-- "10101010" +D10.5+ [426]
		"10101001011",	-- "10101011" +D11.5+ [427]
		"10101101100",	-- "10101100" +D12.5+ [428]
		"10101001101",	-- "10101101" +D13.5+ [429]
		"10101001110",	-- "10101110" +D14.5+ [430]
		"00101000101",	-- "10101111" +D15.5- [431]
		"00101001001",	-- "10110000" +D16.5- [432]
		"10101110001",	-- "10110001" +D17.5+ [433]
		"10101110010",	-- "10110010" +D18.5+ [434]
		"10101010011",	-- "10110011" +D19.5+ [435]
		"10101110100",	-- "10110100" +D20.5+ [436]
		"10101010101",	-- "10110101" +D21.5+ [437]
		"10101010110",	-- "10110110" +D22.5+ [438]
		"00101101000",	-- "10110111" +D23.5- [439]
		"00101001100",	-- "10111000" +D24.5- [440]
		"10101011001",	-- "10111001" +D25.5+ [441]
		"10101011010",	-- "10111010" +D26.5+ [442]
		"00101100100",	-- "10111011" +D27.5- [443]
		"10101011100",	-- "10111100" +D28.5+ [444]
		"00101100010",	-- "10111101" +D29.5- [445]
		"00101100001",	-- "10111110" +D30.5- [446]
		"00101001010",	-- "10111111" +D31.5- [447]
		"00110000110",	-- "11000000" +D00.6- [448]
		"00110010001",	-- "11000001" +D01.6- [449]
		"00110010010",	-- "11000010" +D02.6- [450]
		"10110100011",	-- "11000011" +D03.6+ [451]
		"00110010100",	-- "11000100" +D04.6- [452]
		"10110100101",	-- "11000101" +D05.6+ [453]
		"10110100110",	-- "11000110" +D06.6+ [454]
		"10110111000",	-- "11000111" +D07.6+ [455]
		"00110011000",	-- "11001000" +D08.6- [456]
		"10110101001",	-- "11001001" +D09.6+ [457]
		"10110101010",	-- "11001010" +D10.6+ [458]
		"10110001011",	-- "11001011" +D11.6+ [459]
		"10110101100",	-- "11001100" +D12.6+ [460]
		"10110001101",	-- "11001101" +D13.6+ [461]
		"10110001110",	-- "11001110" +D14.6+ [462]
		"00110000101",	-- "11001111" +D15.6- [463]
		"00110001001",	-- "11010000" +D16.6- [464]
		"10110110001",	-- "11010001" +D17.6+ [465]
		"10110110010",	-- "11010010" +D18.6+ [466]
		"10110010011",	-- "11010011" +D19.6+ [467]
		"10110110100",	-- "11010100" +D20.6+ [468]
		"10110010101",	-- "11010101" +D21.6+ [469]
		"10110010110",	-- "11010110" +D22.6+ [470]
		"00110101000",	-- "11010111" +D23.6- [471]
		"00110001100",	-- "11011000" +D24.6- [472]
		"10110011001",	-- "11011001" +D25.6+ [473]
		"10110011010",	-- "11011010" +D26.6+ [474]
		"00110100100",	-- "11011011" +D27.6- [475]
		"10110011100",	-- "11011100" +D28.6+ [476]
		"00110100010",	-- "11011101" +D29.6- [477]
		"00110100001",	-- "11011110" +D30.6- [478]
		"00110001010",	-- "11011111" +D31.6- [479]
		"10111000110",	-- "11100000" +D00.7+ [480]
		"10111010001",	-- "11100001" +D01.7+ [481]
		"10111010010",	-- "11100010" +D02.7+ [482]
		"01000100011",	-- "11100011" +D03.7- [483]
		"10111010100",	-- "11100100" +D04.7+ [484]
		"01000100101",	-- "11100101" +D05.7- [485]
		"01000100110",	-- "11100110" +D06.7- [486]
		"01000111000",	-- "11100111" +D07.7- [487]
		"10111011000",	-- "11101000" +D08.7+ [488]
		"01000101001",	-- "11101001" +D09.7- [489]
		"01000101010",	-- "11101010" +D10.7- [490]
		"00001001011",	-- "11101011" +D11.7- [491]
		"01000101100",	-- "11101100" +D12.7- [492]
		"00001001101",	-- "11101101" +D13.7- [493]
		"00001001110",	-- "11101110" +D14.7- [494]
		"10111000101",	-- "11101111" +D15.7+ [495]
		"10111001001",	-- "11110000" +D16.7+ [496]
		"01000110001",	-- "11110001" +D17.7- [497]
		"01000110010",	-- "11110010" +D18.7- [498]
		"01000010011",	-- "11110011" +D19.7- [499]
		"01000110100",	-- "11110100" +D20.7- [500]
		"01000010101",	-- "11110101" +D21.7- [501]
		"01000010110",	-- "11110110" +D22.7- [502]
		"10111101000",	-- "11110111" +D23.7+ [503]
		"10111001100",	-- "11111000" +D24.7+ [504]
		"01000011001",	-- "11111001" +D25.7- [505]
		"01000011010",	-- "11111010" +D26.7- [506]
		"10111100100",	-- "11111011" +D27.7+ [507]
		"01000011100",	-- "11111100" +D28.7- [508]
		"10111100010",	-- "11111101" +D29.7+ [509]
		"10111100001",	-- "11111110" +D30.7+ [510]
		"10111001010",	-- "11111111" +D31.7+ [511]
		"00010111001",	-- "00000000" -K00.0- [512]
		"00010101110",	-- "00000001" -K01.0- [513]
		"00010101101",	-- "00000010" -K02.0- [514]
		"11101100011",	-- "00000011" -K03.0+ [515]
		"00010101011",	-- "00000100" -K04.0- [516]
		"11101100101",	-- "00000101" -K05.0+ [517]
		"11101100110",	-- "00000110" -K06.0+ [518]
		"11101000111",	-- "00000111" -K07.0+ [519]
		"00010100111",	-- "00001000" -K08.0- [520]
		"11101101001",	-- "00001001" -K09.0+ [521]
		"11101101010",	-- "00001010" -K10.0+ [522]
		"11101001011",	-- "00001011" -K11.0+ [523]
		"11101101100",	-- "00001100" -K12.0+ [524]
		"11101001101",	-- "00001101" -K13.0+ [525]
		"11101001110",	-- "00001110" -K14.0+ [526]
		"00010111010",	-- "00001111" -K15.0- [527]
		"00010110110",	-- "00010000" -K16.0- [528]
		"11101110001",	-- "00010001" -K17.0+ [529]
		"11101110010",	-- "00010010" -K18.0+ [530]
		"11101010011",	-- "00010011" -K19.0+ [531]
		"11101110100",	-- "00010100" -K20.0+ [532]
		"11101010101",	-- "00010101" -K21.0+ [533]
		"11101010110",	-- "00010110" -K22.0+ [534]
		"00010010111",	-- "00010111" -K23.0- [535]
		"00010110011",	-- "00011000" -K24.0- [536]
		"11101011001",	-- "00011001" -K25.0+ [537]
		"11101011010",	-- "00011010" -K26.0+ [538]
		"00010011011",	-- "00011011" -K27.0- [539]
		"00010111100",	-- "00011100" -K28.0- [540]
		"00010011101",	-- "00011101" -K29.0- [541]
		"00010011110",	-- "00011110" -K30.0- [542]
		"00010110101",	-- "00011111" -K31.0- [543]
		"11001111001",	-- "00100000" -K00.1+ [544]
		"11001101110",	-- "00100001" -K01.1+ [545]
		"11001101101",	-- "00100010" -K02.1+ [546]
		"00110100011",	-- "00100011" -K03.1- [547]
		"11001101011",	-- "00100100" -K04.1+ [548]
		"00110100101",	-- "00100101" -K05.1- [549]
		"00110100110",	-- "00100110" -K06.1- [550]
		"00110000111",	-- "00100111" -K07.1- [551]
		"11001100111",	-- "00101000" -K08.1+ [552]
		"00110101001",	-- "00101001" -K09.1- [553]
		"00110101010",	-- "00101010" -K10.1- [554]
		"00110001011",	-- "00101011" -K11.1- [555]
		"00110101100",	-- "00101100" -K12.1- [556]
		"00110001101",	-- "00101101" -K13.1- [557]
		"00110001110",	-- "00101110" -K14.1- [558]
		"11001111010",	-- "00101111" -K15.1+ [559]
		"11001110110",	-- "00110000" -K16.1+ [560]
		"00110110001",	-- "00110001" -K17.1- [561]
		"00110110010",	-- "00110010" -K18.1- [562]
		"00110010011",	-- "00110011" -K19.1- [563]
		"00110110100",	-- "00110100" -K20.1- [564]
		"00110010101",	-- "00110101" -K21.1- [565]
		"00110010110",	-- "00110110" -K22.1- [566]
		"11001010111",	-- "00110111" -K23.1+ [567]
		"11001110011",	-- "00111000" -K24.1+ [568]
		"00110011001",	-- "00111001" -K25.1- [569]
		"00110011010",	-- "00111010" -K26.1- [570]
		"11001011011",	-- "00111011" -K27.1+ [571]
		"11001111100",	-- "00111100" -K28.1+ [572]
		"11001011101",	-- "00111101" -K29.1+ [573]
		"11001011110",	-- "00111110" -K30.1+ [574]
		"11001110101",	-- "00111111" -K31.1+ [575]
		"11010111001",	-- "01000000" -K00.2+ [576]
		"11010101110",	-- "01000001" -K01.2+ [577]
		"11010101101",	-- "01000010" -K02.2+ [578]
		"00101100011",	-- "01000011" -K03.2- [579]
		"11010101011",	-- "01000100" -K04.2+ [580]
		"00101100101",	-- "01000101" -K05.2- [581]
		"00101100110",	-- "01000110" -K06.2- [582]
		"00101000111",	-- "01000111" -K07.2- [583]
		"11010100111",	-- "01001000" -K08.2+ [584]
		"00101101001",	-- "01001001" -K09.2- [585]
		"00101101010",	-- "01001010" -K10.2- [586]
		"00101001011",	-- "01001011" -K11.2- [587]
		"00101101100",	-- "01001100" -K12.2- [588]
		"00101001101",	-- "01001101" -K13.2- [589]
		"00101001110",	-- "01001110" -K14.2- [590]
		"11010111010",	-- "01001111" -K15.2+ [591]
		"11010110110",	-- "01010000" -K16.2+ [592]
		"00101110001",	-- "01010001" -K17.2- [593]
		"00101110010",	-- "01010010" -K18.2- [594]
		"00101010011",	-- "01010011" -K19.2- [595]
		"00101110100",	-- "01010100" -K20.2- [596]
		"00101010101",	-- "01010101" -K21.2- [597]
		"00101010110",	-- "01010110" -K22.2- [598]
		"11010010111",	-- "01010111" -K23.2+ [599]
		"11010110011",	-- "01011000" -K24.2+ [600]
		"00101011001",	-- "01011001" -K25.2- [601]
		"00101011010",	-- "01011010" -K26.2- [602]
		"11010011011",	-- "01011011" -K27.2+ [603]
		"11010111100",	-- "01011100" -K28.2+ [604]
		"11010011101",	-- "01011101" -K29.2+ [605]
		"11010011110",	-- "01011110" -K30.2+ [606]
		"11010110101",	-- "01011111" -K31.2+ [607]
		"11100111001",	-- "01100000" -K00.3+ [608]
		"11100101110",	-- "01100001" -K01.3+ [609]
		"11100101101",	-- "01100010" -K02.3+ [610]
		"00011100011",	-- "01100011" -K03.3- [611]
		"11100101011",	-- "01100100" -K04.3+ [612]
		"00011100101",	-- "01100101" -K05.3- [613]
		"00011100110",	-- "01100110" -K06.3- [614]
		"00011000111",	-- "01100111" -K07.3- [615]
		"11100100111",	-- "01101000" -K08.3+ [616]
		"00011101001",	-- "01101001" -K09.3- [617]
		"00011101010",	-- "01101010" -K10.3- [618]
		"00011001011",	-- "01101011" -K11.3- [619]
		"00011101100",	-- "01101100" -K12.3- [620]
		"00011001101",	-- "01101101" -K13.3- [621]
		"00011001110",	-- "01101110" -K14.3- [622]
		"11100111010",	-- "01101111" -K15.3+ [623]
		"11100110110",	-- "01110000" -K16.3+ [624]
		"00011110001",	-- "01110001" -K17.3- [625]
		"00011110010",	-- "01110010" -K18.3- [626]
		"00011010011",	-- "01110011" -K19.3- [627]
		"00011110100",	-- "01110100" -K20.3- [628]
		"00011010101",	-- "01110101" -K21.3- [629]
		"00011010110",	-- "01110110" -K22.3- [630]
		"11100010111",	-- "01110111" -K23.3+ [631]
		"11100110011",	-- "01111000" -K24.3+ [632]
		"00011011001",	-- "01111001" -K25.3- [633]
		"00011011010",	-- "01111010" -K26.3- [634]
		"11100011011",	-- "01111011" -K27.3+ [635]
		"11100111100",	-- "01111100" -K28.3+ [636]
		"11100011101",	-- "01111101" -K29.3+ [637]
		"11100011110",	-- "01111110" -K30.3+ [638]
		"11100110101",	-- "01111111" -K31.3+ [639]
		"00100111001",	-- "10000000" -K00.4- [640]
		"00100101110",	-- "10000001" -K01.4- [641]
		"00100101101",	-- "10000010" -K02.4- [642]
		"11011100011",	-- "10000011" -K03.4+ [643]
		"00100101011",	-- "10000100" -K04.4- [644]
		"11011100101",	-- "10000101" -K05.4+ [645]
		"11011100110",	-- "10000110" -K06.4+ [646]
		"11011000111",	-- "10000111" -K07.4+ [647]
		"00100100111",	-- "10001000" -K08.4- [648]
		"11011101001",	-- "10001001" -K09.4+ [649]
		"11011101010",	-- "10001010" -K10.4+ [650]
		"11011001011",	-- "10001011" -K11.4+ [651]
		"11011101100",	-- "10001100" -K12.4+ [652]
		"11011001101",	-- "10001101" -K13.4+ [653]
		"11011001110",	-- "10001110" -K14.4+ [654]
		"00100111010",	-- "10001111" -K15.4- [655]
		"00100110110",	-- "10010000" -K16.4- [656]
		"11011110001",	-- "10010001" -K17.4+ [657]
		"11011110010",	-- "10010010" -K18.4+ [658]
		"11011010011",	-- "10010011" -K19.4+ [659]
		"11011110100",	-- "10010100" -K20.4+ [660]
		"11011010101",	-- "10010101" -K21.4+ [661]
		"11011010110",	-- "10010110" -K22.4+ [662]
		"00100010111",	-- "10010111" -K23.4- [663]
		"00100110011",	-- "10011000" -K24.4- [664]
		"11011011001",	-- "10011001" -K25.4+ [665]
		"11011011010",	-- "10011010" -K26.4+ [666]
		"00100011011",	-- "10011011" -K27.4- [667]
		"00100111100",	-- "10011100" -K28.4- [668]
		"00100011101",	-- "10011101" -K29.4- [669]
		"00100011110",	-- "10011110" -K30.4- [670]
		"00100110101",	-- "10011111" -K31.4- [671]
		"10101111001",	-- "10100000" -K00.5+ [672]
		"10101101110",	-- "10100001" -K01.5+ [673]
		"10101101101",	-- "10100010" -K02.5+ [674]
		"01010100011",	-- "10100011" -K03.5- [675]
		"10101101011",	-- "10100100" -K04.5+ [676]
		"01010100101",	-- "10100101" -K05.5- [677]
		"01010100110",	-- "10100110" -K06.5- [678]
		"01010000111",	-- "10100111" -K07.5- [679]
		"10101100111",	-- "10101000" -K08.5+ [680]
		"01010101001",	-- "10101001" -K09.5- [681]
		"01010101010",	-- "10101010" -K10.5- [682]
		"01010001011",	-- "10101011" -K11.5- [683]
		"01010101100",	-- "10101100" -K12.5- [684]
		"01010001101",	-- "10101101" -K13.5- [685]
		"01010001110",	-- "10101110" -K14.5- [686]
		"10101111010",	-- "10101111" -K15.5+ [687]
		"10101110110",	-- "10110000" -K16.5+ [688]
		"01010110001",	-- "10110001" -K17.5- [689]
		"01010110010",	-- "10110010" -K18.5- [690]
		"01010010011",	-- "10110011" -K19.5- [691]
		"01010110100",	-- "10110100" -K20.5- [692]
		"01010010101",	-- "10110101" -K21.5- [693]
		"01010010110",	-- "10110110" -K22.5- [694]
		"10101010111",	-- "10110111" -K23.5+ [695]
		"10101110011",	-- "10111000" -K24.5+ [696]
		"01010011001",	-- "10111001" -K25.5- [697]
		"01010011010",	-- "10111010" -K26.5- [698]
		"10101011011",	-- "10111011" -K27.5+ [699]
		"10101111100",	-- "10111100" -K28.5+ [700]
		"10101011101",	-- "10111101" -K29.5+ [701]
		"10101011110",	-- "10111110" -K30.5+ [702]
		"10101110101",	-- "10111111" -K31.5+ [703]
		"10110111001",	-- "11000000" -K00.6+ [704]
		"10110101110",	-- "11000001" -K01.6+ [705]
		"10110101101",	-- "11000010" -K02.6+ [706]
		"01001100011",	-- "11000011" -K03.6- [707]
		"10110101011",	-- "11000100" -K04.6+ [708]
		"01001100101",	-- "11000101" -K05.6- [709]
		"01001100110",	-- "11000110" -K06.6- [710]
		"01001000111",	-- "11000111" -K07.6- [711]
		"10110100111",	-- "11001000" -K08.6+ [712]
		"01001101001",	-- "11001001" -K09.6- [713]
		"01001101010",	-- "11001010" -K10.6- [714]
		"01001001011",	-- "11001011" -K11.6- [715]
		"01001101100",	-- "11001100" -K12.6- [716]
		"01001001101",	-- "11001101" -K13.6- [717]
		"01001001110",	-- "11001110" -K14.6- [718]
		"10110111010",	-- "11001111" -K15.6+ [719]
		"10110110110",	-- "11010000" -K16.6+ [720]
		"01001110001",	-- "11010001" -K17.6- [721]
		"01001110010",	-- "11010010" -K18.6- [722]
		"01001010011",	-- "11010011" -K19.6- [723]
		"01001110100",	-- "11010100" -K20.6- [724]
		"01001010101",	-- "11010101" -K21.6- [725]
		"01001010110",	-- "11010110" -K22.6- [726]
		"10110010111",	-- "11010111" -K23.6+ [727]
		"10110110011",	-- "11011000" -K24.6+ [728]
		"01001011001",	-- "11011001" -K25.6- [729]
		"01001011010",	-- "11011010" -K26.6- [730]
		"10110011011",	-- "11011011" -K27.6+ [731]
		"10110111100",	-- "11011100" -K28.6+ [732]
		"10110011101",	-- "11011101" -K29.6+ [733]
		"10110011110",	-- "11011110" -K30.6+ [734]
		"10110110101",	-- "11011111" -K31.6+ [735]
		"00001111001",	-- "11100000" -K00.7- [736]
		"00001101110",	-- "11100001" -K01.7- [737]
		"00001101101",	-- "11100010" -K02.7- [738]
		"11110100011",	-- "11100011" -K03.7+ [739]
		"00001101011",	-- "11100100" -K04.7- [740]
		"11110100101",	-- "11100101" -K05.7+ [741]
		"11110100110",	-- "11100110" -K06.7+ [742]
		"11110000111",	-- "11100111" -K07.7+ [743]
		"00001100111",	-- "11101000" -K08.7- [744]
		"11110101001",	-- "11101001" -K09.7+ [745]
		"11110101010",	-- "11101010" -K10.7+ [746]
		"11110001011",	-- "11101011" -K11.7+ [747]
		"11110101100",	-- "11101100" -K12.7+ [748]
		"11110001101",	-- "11101101" -K13.7+ [749]
		"11110001110",	-- "11101110" -K14.7+ [750]
		"00001111010",	-- "11101111" -K15.7- [751]
		"00001110110",	-- "11110000" -K16.7- [752]
		"11110110001",	-- "11110001" -K17.7+ [753]
		"11110110010",	-- "11110010" -K18.7+ [754]
		"11110010011",	-- "11110011" -K19.7+ [755]
		"11110110100",	-- "11110100" -K20.7+ [756]
		"11110010101",	-- "11110101" -K21.7+ [757]
		"11110010110",	-- "11110110" -K22.7+ [758]
		"00001010111",	-- "11110111" -K23.7- [759]
		"00001110011",	-- "11111000" -K24.7- [760]
		"11110011001",	-- "11111001" -K25.7+ [761]
		"11110011010",	-- "11111010" -K26.7+ [762]
		"00001011011",	-- "11111011" -K27.7- [763]
		"00001111100",	-- "11111100" -K28.7- [764]
		"00001011101",	-- "11111101" -K29.7- [765]
		"00001011110",	-- "11111110" -K30.7- [766]
		"00001110101",	-- "11111111" -K31.7- [767]
		"11101000110",	-- "00000000" +K00.0+ [768]
		"11101010001",	-- "00000001" +K01.0+ [769]
		"11101010010",	-- "00000010" +K02.0+ [770]
		"00010100011",	-- "00000011" +K03.0- [771]
		"11101010100",	-- "00000100" +K04.0+ [772]
		"00010100101",	-- "00000101" +K05.0- [773]
		"00010100110",	-- "00000110" +K06.0- [774]
		"00010111000",	-- "00000111" +K07.0- [775]
		"11101011000",	-- "00001000" +K08.0+ [776]
		"00010101001",	-- "00001001" +K09.0- [777]
		"00010101010",	-- "00001010" +K10.0- [778]
		"00010001011",	-- "00001011" +K11.0- [779]
		"00010101100",	-- "00001100" +K12.0- [780]
		"00010001101",	-- "00001101" +K13.0- [781]
		"00010001110",	-- "00001110" +K14.0- [782]
		"11101000101",	-- "00001111" +K15.0+ [783]
		"11101001001",	-- "00010000" +K16.0+ [784]
		"00010110001",	-- "00010001" +K17.0- [785]
		"00010110010",	-- "00010010" +K18.0- [786]
		"00010010011",	-- "00010011" +K19.0- [787]
		"00010110100",	-- "00010100" +K20.0- [788]
		"00010010101",	-- "00010101" +K21.0- [789]
		"00010010110",	-- "00010110" +K22.0- [790]
		"11101101000",	-- "00010111" +K23.0+ [791]
		"11101001100",	-- "00011000" +K24.0+ [792]
		"00010011001",	-- "00011001" +K25.0- [793]
		"00010011010",	-- "00011010" +K26.0- [794]
		"11101100100",	-- "00011011" +K27.0+ [795]
		"11101000011",	-- "00011100" +K28.0+ [796]
		"11101100010",	-- "00011101" +K29.0+ [797]
		"11101100001",	-- "00011110" +K30.0+ [798]
		"11101001010",	-- "00011111" +K31.0+ [799]
		"00110000110",	-- "00100000" +K00.1- [800]
		"00110010001",	-- "00100001" +K01.1- [801]
		"00110010010",	-- "00100010" +K02.1- [802]
		"11001100011",	-- "00100011" +K03.1+ [803]
		"00110010100",	-- "00100100" +K04.1- [804]
		"11001100101",	-- "00100101" +K05.1+ [805]
		"11001100110",	-- "00100110" +K06.1+ [806]
		"11001111000",	-- "00100111" +K07.1+ [807]
		"00110011000",	-- "00101000" +K08.1- [808]
		"11001101001",	-- "00101001" +K09.1+ [809]
		"11001101010",	-- "00101010" +K10.1+ [810]
		"11001001011",	-- "00101011" +K11.1+ [811]
		"11001101100",	-- "00101100" +K12.1+ [812]
		"11001001101",	-- "00101101" +K13.1+ [813]
		"11001001110",	-- "00101110" +K14.1+ [814]
		"00110000101",	-- "00101111" +K15.1- [815]
		"00110001001",	-- "00110000" +K16.1- [816]
		"11001110001",	-- "00110001" +K17.1+ [817]
		"11001110010",	-- "00110010" +K18.1+ [818]
		"11001010011",	-- "00110011" +K19.1+ [819]
		"11001110100",	-- "00110100" +K20.1+ [820]
		"11001010101",	-- "00110101" +K21.1+ [821]
		"11001010110",	-- "00110110" +K22.1+ [822]
		"00110101000",	-- "00110111" +K23.1- [823]
		"00110001100",	-- "00111000" +K24.1- [824]
		"11001011001",	-- "00111001" +K25.1+ [825]
		"11001011010",	-- "00111010" +K26.1+ [826]
		"00110100100",	-- "00111011" +K27.1- [827]
		"00110000011",	-- "00111100" +K28.1- [828]
		"00110100010",	-- "00111101" +K29.1- [829]
		"00110100001",	-- "00111110" +K30.1- [830]
		"00110001010",	-- "00111111" +K31.1- [831]
		"00101000110",	-- "01000000" +K00.2- [832]
		"00101010001",	-- "01000001" +K01.2- [833]
		"00101010010",	-- "01000010" +K02.2- [834]
		"11010100011",	-- "01000011" +K03.2+ [835]
		"00101010100",	-- "01000100" +K04.2- [836]
		"11010100101",	-- "01000101" +K05.2+ [837]
		"11010100110",	-- "01000110" +K06.2+ [838]
		"11010111000",	-- "01000111" +K07.2+ [839]
		"00101011000",	-- "01001000" +K08.2- [840]
		"11010101001",	-- "01001001" +K09.2+ [841]
		"11010101010",	-- "01001010" +K10.2+ [842]
		"11010001011",	-- "01001011" +K11.2+ [843]
		"11010101100",	-- "01001100" +K12.2+ [844]
		"11010001101",	-- "01001101" +K13.2+ [845]
		"11010001110",	-- "01001110" +K14.2+ [846]
		"00101000101",	-- "01001111" +K15.2- [847]
		"00101001001",	-- "01010000" +K16.2- [848]
		"11010110001",	-- "01010001" +K17.2+ [849]
		"11010110010",	-- "01010010" +K18.2+ [850]
		"11010010011",	-- "01010011" +K19.2+ [851]
		"11010110100",	-- "01010100" +K20.2+ [852]
		"11010010101",	-- "01010101" +K21.2+ [853]
		"11010010110",	-- "01010110" +K22.2+ [854]
		"00101101000",	-- "01010111" +K23.2- [855]
		"00101001100",	-- "01011000" +K24.2- [856]
		"11010011001",	-- "01011001" +K25.2+ [857]
		"11010011010",	-- "01011010" +K26.2+ [858]
		"00101100100",	-- "01011011" +K27.2- [859]
		"00101000011",	-- "01011100" +K28.2- [860]
		"00101100010",	-- "01011101" +K29.2- [861]
		"00101100001",	-- "01011110" +K30.2- [862]
		"00101001010",	-- "01011111" +K31.2- [863]
		"00011000110",	-- "01100000" +K00.3- [864]
		"00011010001",	-- "01100001" +K01.3- [865]
		"00011010010",	-- "01100010" +K02.3- [866]
		"11100100011",	-- "01100011" +K03.3+ [867]
		"00011010100",	-- "01100100" +K04.3- [868]
		"11100100101",	-- "01100101" +K05.3+ [869]
		"11100100110",	-- "01100110" +K06.3+ [870]
		"11100111000",	-- "01100111" +K07.3+ [871]
		"00011011000",	-- "01101000" +K08.3- [872]
		"11100101001",	-- "01101001" +K09.3+ [873]
		"11100101010",	-- "01101010" +K10.3+ [874]
		"11100001011",	-- "01101011" +K11.3+ [875]
		"11100101100",	-- "01101100" +K12.3+ [876]
		"11100001101",	-- "01101101" +K13.3+ [877]
		"11100001110",	-- "01101110" +K14.3+ [878]
		"00011000101",	-- "01101111" +K15.3- [879]
		"00011001001",	-- "01110000" +K16.3- [880]
		"11100110001",	-- "01110001" +K17.3+ [881]
		"11100110010",	-- "01110010" +K18.3+ [882]
		"11100010011",	-- "01110011" +K19.3+ [883]
		"11100110100",	-- "01110100" +K20.3+ [884]
		"11100010101",	-- "01110101" +K21.3+ [885]
		"11100010110",	-- "01110110" +K22.3+ [886]
		"00011101000",	-- "01110111" +K23.3- [887]
		"00011001100",	-- "01111000" +K24.3- [888]
		"11100011001",	-- "01111001" +K25.3+ [889]
		"11100011010",	-- "01111010" +K26.3+ [890]
		"00011100100",	-- "01111011" +K27.3- [891]
		"00011000011",	-- "01111100" +K28.3- [892]
		"00011100010",	-- "01111101" +K29.3- [893]
		"00011100001",	-- "01111110" +K30.3- [894]
		"00011001010",	-- "01111111" +K31.3- [895]
		"11011000110",	-- "10000000" +K00.4+ [896]
		"11011010001",	-- "10000001" +K01.4+ [897]
		"11011010010",	-- "10000010" +K02.4+ [898]
		"00100100011",	-- "10000011" +K03.4- [899]
		"11011010100",	-- "10000100" +K04.4+ [900]
		"00100100101",	-- "10000101" +K05.4- [901]
		"00100100110",	-- "10000110" +K06.4- [902]
		"00100111000",	-- "10000111" +K07.4- [903]
		"11011011000",	-- "10001000" +K08.4+ [904]
		"00100101001",	-- "10001001" +K09.4- [905]
		"00100101010",	-- "10001010" +K10.4- [906]
		"00100001011",	-- "10001011" +K11.4- [907]
		"00100101100",	-- "10001100" +K12.4- [908]
		"00100001101",	-- "10001101" +K13.4- [909]
		"00100001110",	-- "10001110" +K14.4- [910]
		"11011000101",	-- "10001111" +K15.4+ [911]
		"11011001001",	-- "10010000" +K16.4+ [912]
		"00100110001",	-- "10010001" +K17.4- [913]
		"00100110010",	-- "10010010" +K18.4- [914]
		"00100010011",	-- "10010011" +K19.4- [915]
		"00100110100",	-- "10010100" +K20.4- [916]
		"00100010101",	-- "10010101" +K21.4- [917]
		"00100010110",	-- "10010110" +K22.4- [918]
		"11011101000",	-- "10010111" +K23.4+ [919]
		"11011001100",	-- "10011000" +K24.4+ [920]
		"00100011001",	-- "10011001" +K25.4- [921]
		"00100011010",	-- "10011010" +K26.4- [922]
		"11011100100",	-- "10011011" +K27.4+ [923]
		"11011000011",	-- "10011100" +K28.4+ [924]
		"11011100010",	-- "10011101" +K29.4+ [925]
		"11011100001",	-- "10011110" +K30.4+ [926]
		"11011001010",	-- "10011111" +K31.4+ [927]
		"01010000110",	-- "10100000" +K00.5- [928]
		"01010010001",	-- "10100001" +K01.5- [929]
		"01010010010",	-- "10100010" +K02.5- [930]
		"10101100011",	-- "10100011" +K03.5+ [931]
		"01010010100",	-- "10100100" +K04.5- [932]
		"10101100101",	-- "10100101" +K05.5+ [933]
		"10101100110",	-- "10100110" +K06.5+ [934]
		"10101111000",	-- "10100111" +K07.5+ [935]
		"01010011000",	-- "10101000" +K08.5- [936]
		"10101101001",	-- "10101001" +K09.5+ [937]
		"10101101010",	-- "10101010" +K10.5+ [938]
		"10101001011",	-- "10101011" +K11.5+ [939]
		"10101101100",	-- "10101100" +K12.5+ [940]
		"10101001101",	-- "10101101" +K13.5+ [941]
		"10101001110",	-- "10101110" +K14.5+ [942]
		"01010000101",	-- "10101111" +K15.5- [943]
		"01010001001",	-- "10110000" +K16.5- [944]
		"10101110001",	-- "10110001" +K17.5+ [945]
		"10101110010",	-- "10110010" +K18.5+ [946]
		"10101010011",	-- "10110011" +K19.5+ [947]
		"10101110100",	-- "10110100" +K20.5+ [948]
		"10101010101",	-- "10110101" +K21.5+ [949]
		"10101010110",	-- "10110110" +K22.5+ [950]
		"01010101000",	-- "10110111" +K23.5- [951]
		"01010001100",	-- "10111000" +K24.5- [952]
		"10101011001",	-- "10111001" +K25.5+ [953]
		"10101011010",	-- "10111010" +K26.5+ [954]
		"01010100100",	-- "10111011" +K27.5- [955]
		"01010000011",	-- "10111100" +K28.5- [956]
		"01010100010",	-- "10111101" +K29.5- [957]
		"01010100001",	-- "10111110" +K30.5- [958]
		"01010001010",	-- "10111111" +K31.5- [959]
		"01001000110",	-- "11000000" +K00.6- [960]
		"01001010001",	-- "11000001" +K01.6- [961]
		"01001010010",	-- "11000010" +K02.6- [962]
		"10110100011",	-- "11000011" +K03.6+ [963]
		"01001010100",	-- "11000100" +K04.6- [964]
		"10110100101",	-- "11000101" +K05.6+ [965]
		"10110100110",	-- "11000110" +K06.6+ [966]
		"10110111000",	-- "11000111" +K07.6+ [967]
		"01001011000",	-- "11001000" +K08.6- [968]
		"10110101001",	-- "11001001" +K09.6+ [969]
		"10110101010",	-- "11001010" +K10.6+ [970]
		"10110001011",	-- "11001011" +K11.6+ [971]
		"10110101100",	-- "11001100" +K12.6+ [972]
		"10110001101",	-- "11001101" +K13.6+ [973]
		"10110001110",	-- "11001110" +K14.6+ [974]
		"01001000101",	-- "11001111" +K15.6- [975]
		"01001001001",	-- "11010000" +K16.6- [976]
		"10110110001",	-- "11010001" +K17.6+ [977]
		"10110110010",	-- "11010010" +K18.6+ [978]
		"10110010011",	-- "11010011" +K19.6+ [979]
		"10110110100",	-- "11010100" +K20.6+ [980]
		"10110010101",	-- "11010101" +K21.6+ [981]
		"10110010110",	-- "11010110" +K22.6+ [982]
		"01001101000",	-- "11010111" +K23.6- [983]
		"01001001100",	-- "11011000" +K24.6- [984]
		"10110011001",	-- "11011001" +K25.6+ [985]
		"10110011010",	-- "11011010" +K26.6+ [986]
		"01001100100",	-- "11011011" +K27.6- [987]
		"01001000011",	-- "11011100" +K28.6- [988]
		"01001100010",	-- "11011101" +K29.6- [989]
		"01001100001",	-- "11011110" +K30.6- [990]
		"01001001010",	-- "11011111" +K31.6- [991]
		"11110000110",	-- "11100000" +K00.7+ [992]
		"11110010001",	-- "11100001" +K01.7+ [993]
		"11110010010",	-- "11100010" +K02.7+ [994]
		"00001100011",	-- "11100011" +K03.7- [995]
		"11110010100",	-- "11100100" +K04.7+ [996]
		"00001100101",	-- "11100101" +K05.7- [997]
		"00001100110",	-- "11100110" +K06.7- [998]
		"00001111000",	-- "11100111" +K07.7- [999]
		"11110011000",	-- "11101000" +K08.7+ [1000]
		"00001101001",	-- "11101001" +K09.7- [1001]
		"00001101010",	-- "11101010" +K10.7- [1002]
		"00001001011",	-- "11101011" +K11.7- [1003]
		"00001101100",	-- "11101100" +K12.7- [1004]
		"00001001101",	-- "11101101" +K13.7- [1005]
		"00001001110",	-- "11101110" +K14.7- [1006]
		"11110000101",	-- "11101111" +K15.7+ [1007]
		"11110001001",	-- "11110000" +K16.7+ [1008]
		"00001110001",	-- "11110001" +K17.7- [1009]
		"00001110010",	-- "11110010" +K18.7- [1010]
		"00001010011",	-- "11110011" +K19.7- [1011]
		"00001110100",	-- "11110100" +K20.7- [1012]
		"00001010101",	-- "11110101" +K21.7- [1013]
		"00001010110",	-- "11110110" +K22.7- [1014]
		"11110101000",	-- "11110111" +K23.7+ [1015]
		"11110001100",	-- "11111000" +K24.7+ [1016]
		"00001011001",	-- "11111001" +K25.7- [1017]
		"00001011010",	-- "11111010" +K26.7- [1018]
		"11110100100",	-- "11111011" +K27.7+ [1019]
		"11110000011",	-- "11111100" +K28.7+ [1020]
		"11110100010",	-- "11111101" +K29.7+ [1021]
		"11110100001",	-- "11111110" +K30.7+ [1022]
		"11110001010"	-- "11111111" +K31.7+ [1023]
	);

constant ENC_K28D0R0 : std_logic_vector := "00010111100";	-- -1 + K28.0 => -1
constant ENC_K28D1R0 : std_logic_vector := "11001111100";	-- -1 + K28.1 => 1
constant ENC_K28D2R0 : std_logic_vector := "11010111100";	-- -1 + K28.2 => 1
constant ENC_K28D3R0 : std_logic_vector := "11100111100";	-- -1 + K28.3 => 1
constant ENC_K28D4R0 : std_logic_vector := "00100111100";	-- -1 + K28.4 => -1
constant ENC_K28D5R0 : std_logic_vector := "10101111100";	-- -1 + K28.5 => 1

constant ENC_K28D6R0 : std_logic_vector := "10110111100";	-- -1 + K28.6 => 1
constant ENC_K28D7R0 : std_logic_vector := "00001111100";	-- -1 + K28.7 => -1
constant ENC_K23D7R0 : std_logic_vector := "00001010111";	-- -1 + K23.7 => -1
constant ENC_K27D7R0 : std_logic_vector := "00001011011";	-- -1 + K27.7 => -1
constant ENC_K29D7R0 : std_logic_vector := "00001011101";	-- -1 + K29.7 => -1
constant ENC_K30D7R0 : std_logic_vector := "00001011110";	-- -1 + K30.7 => -1
constant ENC_K28D0R1 : std_logic_vector := "11101000011";	-- 1 + K28.0 => 1
constant ENC_K28D1R1 : std_logic_vector := "00110000011";	-- 1 + K28.1 => -1
constant ENC_K28D2R1 : std_logic_vector := "00101000011";	-- 1 + K28.2 => -1
constant ENC_K28D3R1 : std_logic_vector := "00011000011";	-- 1 + K28.3 => -1
constant ENC_K28D4R1 : std_logic_vector := "11011000011";	-- 1 + K28.4 => 1
constant ENC_K28D5R1 : std_logic_vector := "01010000011";	-- 1 + K28.5 => -1
constant ENC_K28D6R1 : std_logic_vector := "01001000011";	-- 1 + K28.6 => -1
constant ENC_K28D7R1 : std_logic_vector := "11110000011";	-- 1 + K28.7 => 1
constant ENC_K23D7R1 : std_logic_vector := "11110101000";	-- 1 + K23.7 => 1
constant ENC_K27D7R1 : std_logic_vector := "11110100100";	-- 1 + K27.7 => 1
constant ENC_K29D7R1 : std_logic_vector := "11110100010";	-- 1 + K29.7 => 1
constant ENC_K30D7R1 : std_logic_vector := "11110100001";	-- 1 + K30.7 => 1
constant DEC_K28D0 : std_logic_vector := "00011100";	-- K28.0
constant DEC_K28D1 : std_logic_vector := "00111100";	-- K28.1
constant DEC_K28D2 : std_logic_vector := "01011100";	-- K28.2
constant DEC_K28D3 : std_logic_vector := "01111100";	-- K28.3
constant DEC_K28D4 : std_logic_vector := "10011100";	-- K28.4
constant DEC_K28D5 : std_logic_vector := "10111100";	-- K28.5
constant DEC_K28D6 : std_logic_vector := "11011100";	-- K28.6
constant DEC_K28D7 : std_logic_vector := "11111100";	-- K28.7
constant DEC_K23D7 : std_logic_vector := "11110111";	-- K23.7
constant DEC_K27D7 : std_logic_vector := "11111011";	-- K27.7
constant DEC_K29D7 : std_logic_vector := "11111101";	-- K29.7
constant DEC_K30D7 : std_logic_vector := "11111110";	-- K30.7

signal ENCODE : std_logic_vector (10 downto 0);
begin

	RUNDP_OUT <= ENCODE(10);
	ENCODE_OUT <= ENCODE(9 downto 0);
	
	process (CLK_IN)
	begin
		if (CLK_IN='1' and CLK_IN'event)
		then
			ENCODE <= TBL_ENC8b10b(conv_integer(CTRL_IN & ((not RUNDP_RESET_IN) and ENCODE(10)) & DATA_IN));
		end if;
	end process;

end RTL;

