//-------------------------------------------------------------------------
//
// File name    :  ldpc_edgetable.v
// Title        :
//              :
// Purpose      : ROM, holds DVB-S2 edge table
//              : Format:
//              : Code pointer: points to the beginning of a code group
//              :   address[12:0]
//              :
//              : Line descriptor : describes the group of parity
//              :                   descriptors that follow
//              :   bits 13:9: # of parity descriptors in this group
//              :   bit 8: indicate that this is the last group of
//              :          parity descriptors for this code group
//              :   bits 7:0: q value for this group
//              : 
//              : Parity descriptor
//              :   bits 15:9: parity location/q, indicates the distance
//              :              to shift VN input to align with CN
//              :   bits 8:0: parity location MOD q, indicates the CN
//              :             address for this check node
//
// ----------------------------------------------------------------------
// Revision History :
// ----------------------------------------------------------------------
//   Ver  :| Author   :| Mod. Date   :| Changes Made:
//   v1.0  | JTC      :| 2008/07/02  :|
// ----------------------------------------------------------------------
`timescale 1ns/10ps

module ldpc_edgetable(
  input        clk,
  input        rst,
  input[12:0]  romaddr,
  output[16:0] romdata
);

reg[16:0] romdata_int;

assign romdata = romdata_int;

always @( posedge rst, posedge clk )
  if( rst )
    romdata_int <= 0;
  else
  case( romaddr )
    0: romdata_int  <= 'h15;   // Code pointer for 1_4
    1: romdata_int  <= 'h150;  // Code pointer for 1_3
    2: romdata_int  <= 'h2f4;  // Code pointer for 2_5
    3: romdata_int  <= 'h4ec;  // Code pointer for 1_2
    4: romdata_int  <= 'h708;  // Code pointer for 3_5
    5: romdata_int  <= 'h9fc;  // Code pointer for 2_3
    6: romdata_int  <= 'hc54;  // Code pointer for 3_4
    7: romdata_int  <= 'hef7;  // Code pointer for 4_5
    8: romdata_int  <= 'h11c7; // Code pointer for 5_6
    9: romdata_int  <= 'h14b5; // Code pointer for 8_9
    10: romdata_int <= 'h1749; // Code pointer for 9_10
    11: romdata_int <= 'h19e3; // Code pointer for 1_5s
    12: romdata_int <= 'h1a2b; // Code pointer for 1_3s
    13: romdata_int <= 'h1a94; // Code pointer for 2_5s
    14: romdata_int <= 'h1b12; // Code pointer for 4_9s
    15: romdata_int <= 'h1b7b; // Code pointer for 3_5s
    16: romdata_int <= 'h1c38; // Code pointer for 2_3s
    17: romdata_int <= 'h1cce; // Code pointer for 11_15s
    18: romdata_int <= 'h1d5b; // Code pointer for 7_9s
    19: romdata_int <= 'h1de7; // Code pointer for 37_45s
    20: romdata_int <= 'h1e85; // Code pointer for 8_9s
    21: romdata_int <= 'h1687; // Line Descriptor
    22: romdata_int <= 'he8ae;
    23: romdata_int <= 'h6b0b;
    24: romdata_int <= 'h7808;
    25: romdata_int <= 'hd0d5;
    26: romdata_int <= 'h7486;
    27: romdata_int <= 'h1e89;
    28: romdata_int <= 'h202e;
    29: romdata_int <= 'h4;
    30: romdata_int <= 'h3b37;
    31: romdata_int <= 'hb29a;
    32: romdata_int <= 'h54b0;
    33: romdata_int <= 'hd95c;
    34: romdata_int <= 'h1687; // Line Descriptor
    35: romdata_int <= 'ha879;
    36: romdata_int <= 'hb0b8;
    37: romdata_int <= 'h87b;
    38: romdata_int <= 'hce7f;
    39: romdata_int <= 'h10a38;
    40: romdata_int <= 'h2cb9;
    41: romdata_int <= 'h7d3b;
    42: romdata_int <= 'hec7c;
    43: romdata_int <= 'hb702;
    44: romdata_int <= 'hea9b;
    45: romdata_int <= 'h4512;
    46: romdata_int <= 'h4a99;
    47: romdata_int <= 'h1687; // Line Descriptor
    48: romdata_int <= 'hee0d;
    49: romdata_int <= 'h10d28;
    50: romdata_int <= 'h948a;
    51: romdata_int <= 'h3a6b;
    52: romdata_int <= 'hc667;
    53: romdata_int <= 'h5855;
    54: romdata_int <= 'h1661;
    55: romdata_int <= 'h8ed5;
    56: romdata_int <= 'h771e;
    57: romdata_int <= 'hb0a5;
    58: romdata_int <= 'h1ee0;
    59: romdata_int <= 'h6ee6;
    60: romdata_int <= 'h1687; // Line Descriptor
    61: romdata_int <= 'he4a4;
    62: romdata_int <= 'h812c;
    63: romdata_int <= 'hc8a7;
    64: romdata_int <= 'hf4a6;
    65: romdata_int <= 'h762d;
    66: romdata_int <= 'h10643;
    67: romdata_int <= 'h4d28;
    68: romdata_int <= 'h108b0;
    69: romdata_int <= 'h3642;
    70: romdata_int <= 'ha673;
    71: romdata_int <= 'he47c;
    72: romdata_int <= 'hbce5;
    73: romdata_int <= 'h1687; // Line Descriptor
    74: romdata_int <= 'h903b;
    75: romdata_int <= 'h492b;
    76: romdata_int <= 'h6464;
    77: romdata_int <= 'hac90;
    78: romdata_int <= 'h6936;
    79: romdata_int <= 'h36d5;
    80: romdata_int <= 'h9462;
    81: romdata_int <= 'hfcf2;
    82: romdata_int <= 'hdab6;
    83: romdata_int <= 'hac9;
    84: romdata_int <= 'ha154;
    85: romdata_int <= 'h3e4a;
    86: romdata_int <= 'h1687; // Line Descriptor
    87: romdata_int <= 'h512c;
    88: romdata_int <= 'ha749;
    89: romdata_int <= 'hc67;
    90: romdata_int <= 'h32a6;
    91: romdata_int <= 'h3ef2;
    92: romdata_int <= 'h5a88;
    93: romdata_int <= 'hd127;
    94: romdata_int <= 'hcbd;
    95: romdata_int <= 'h9a5c;
    96: romdata_int <= 'h10648;
    97: romdata_int <= 'h9322;
    98: romdata_int <= 'h10101;
    99: romdata_int <= 'h1687; // Line Descriptor
    100: romdata_int <= 'he270;
    101: romdata_int <= 'hd94f;
    102: romdata_int <= 'h5c25;
    103: romdata_int <= 'h314d;
    104: romdata_int <= 'ha152;
    105: romdata_int <= 'h3d38;
    106: romdata_int <= 'hde8f;
    107: romdata_int <= 'h40e;
    108: romdata_int <= 'h48ab;
    109: romdata_int <= 'h8275;
    110: romdata_int <= 'h7241;
    111: romdata_int <= 'h604c;
    112: romdata_int <= 'h1687; // Line Descriptor
    113: romdata_int <= 'h924d;
    114: romdata_int <= 'h2148;
    115: romdata_int <= 'hca1a;
    116: romdata_int <= 'h1040a;
    117: romdata_int <= 'h6716;
    118: romdata_int <= 'hf8ee;
    119: romdata_int <= 'h5e66;
    120: romdata_int <= 'h10a32;
    121: romdata_int <= 'haef3;
    122: romdata_int <= 'h392a;
    123: romdata_int <= 'hc558;
    124: romdata_int <= 'h7858;
    125: romdata_int <= 'h1687; // Line Descriptor
    126: romdata_int <= 'hb431;
    127: romdata_int <= 'h44a0;
    128: romdata_int <= 'h8cd0;
    129: romdata_int <= 'h2344;
    130: romdata_int <= 'haa06;
    131: romdata_int <= 'h8630;
    132: romdata_int <= 'h5a9b;
    133: romdata_int <= 'h30d6;
    134: romdata_int <= 'h18df;
    135: romdata_int <= 'hacbe;
    136: romdata_int <= 'h2735;
    137: romdata_int <= 'h6854;
    138: romdata_int <= 'h1687; // Line Descriptor
    139: romdata_int <= 'h108a2;
    140: romdata_int <= 'h8a2a;
    141: romdata_int <= 'h96c9;
    142: romdata_int <= 'h24ce;
    143: romdata_int <= 'h4afd;
    144: romdata_int <= 'h7319;
    145: romdata_int <= 'he650;
    146: romdata_int <= 'he233;
    147: romdata_int <= 'h581c;
    148: romdata_int <= 'h1538;
    149: romdata_int <= 'h4e21;
    150: romdata_int <= 'hc708;
    151: romdata_int <= 'h1687; // Line Descriptor
    152: romdata_int <= 'h143f;
    153: romdata_int <= 'hde08;
    154: romdata_int <= 'he65;
    155: romdata_int <= 'h46e5;
    156: romdata_int <= 'h2ec0;
    157: romdata_int <= 'hec5d;
    158: romdata_int <= 'hf27b;
    159: romdata_int <= 'hd4fd;
    160: romdata_int <= 'hceeb;
    161: romdata_int <= 'hc818;
    162: romdata_int <= 'hd640;
    163: romdata_int <= 'h9722;
    164: romdata_int <= 'h1687; // Line Descriptor
    165: romdata_int <= 'h9e8c;
    166: romdata_int <= 'h607e;
    167: romdata_int <= 'h833f;
    168: romdata_int <= 'h7a1f;
    169: romdata_int <= 'h8823;
    170: romdata_int <= 'h2946;
    171: romdata_int <= 'h1c90;
    172: romdata_int <= 'ha2da;
    173: romdata_int <= 'h963;
    174: romdata_int <= 'h6c70;
    175: romdata_int <= 'h42b4;
    176: romdata_int <= 'h628f;
    177: romdata_int <= 'h1687; // Line Descriptor
    178: romdata_int <= 'hb27b;
    179: romdata_int <= 'h163e;
    180: romdata_int <= 'h9adb;
    181: romdata_int <= 'h9958;
    182: romdata_int <= 'hbcee;
    183: romdata_int <= 'h26c3;
    184: romdata_int <= 'hb445;
    185: romdata_int <= 'h8687;
    186: romdata_int <= 'h225c;
    187: romdata_int <= 'h5cca;
    188: romdata_int <= 'hc106;
    189: romdata_int <= 'hf37;
    190: romdata_int <= 'h1687; // Line Descriptor
    191: romdata_int <= 'hea73;
    192: romdata_int <= 'h842b;
    193: romdata_int <= 'h6358;
    194: romdata_int <= 'h100c5;
    195: romdata_int <= 'h52ad;
    196: romdata_int <= 'hcc35;
    197: romdata_int <= 'h8042;
    198: romdata_int <= 'h6617;
    199: romdata_int <= 'h3315;
    200: romdata_int <= 'h74c;
    201: romdata_int <= 'h6b06;
    202: romdata_int <= 'h5264;
    203: romdata_int <= 'h1687; // Line Descriptor
    204: romdata_int <= 'h7f3d;
    205: romdata_int <= 'h1aed;
    206: romdata_int <= 'hd731;
    207: romdata_int <= 'h391f;
    208: romdata_int <= 'hdcc4;
    209: romdata_int <= 'h414;
    210: romdata_int <= 'hfac9;
    211: romdata_int <= 'h1035b;
    212: romdata_int <= 'hee0a;
    213: romdata_int <= 'hc29a;
    214: romdata_int <= 'h2acb;
    215: romdata_int <= 'h9d1d;
    216: romdata_int <= 'h487; // Line Descriptor
    217: romdata_int <= 'h18a4;
    218: romdata_int <= 'hc0b3;
    219: romdata_int <= 'h7c3d;
    220: romdata_int <= 'h487; // Line Descriptor
    221: romdata_int <= 'h548f;
    222: romdata_int <= 'hf649;
    223: romdata_int <= 'hfecd;
    224: romdata_int <= 'h487; // Line Descriptor
    225: romdata_int <= 'h3503;
    226: romdata_int <= 'h122f;
    227: romdata_int <= 'ha2f8;
    228: romdata_int <= 'h487; // Line Descriptor
    229: romdata_int <= 'ha4dc;
    230: romdata_int <= 'hbee4;
    231: romdata_int <= 'hbada;
    232: romdata_int <= 'h487; // Line Descriptor
    233: romdata_int <= 'hc444;
    234: romdata_int <= 'h5f67;
    235: romdata_int <= 'h4e6a;
    236: romdata_int <= 'h487; // Line Descriptor
    237: romdata_int <= 'hfd19;
    238: romdata_int <= 'he61e;
    239: romdata_int <= 'h745;
    240: romdata_int <= 'h487; // Line Descriptor
    241: romdata_int <= 'h563f;
    242: romdata_int <= 'hc2f5;
    243: romdata_int <= 'hf0fe;
    244: romdata_int <= 'h487; // Line Descriptor
    245: romdata_int <= 'hfaa6;
    246: romdata_int <= 'h70d5;
    247: romdata_int <= 'h6eb1;
    248: romdata_int <= 'h487; // Line Descriptor
    249: romdata_int <= 'h6c97;
    250: romdata_int <= 'he01d;
    251: romdata_int <= 'h2ab3;
    252: romdata_int <= 'h487; // Line Descriptor
    253: romdata_int <= 'h111e;
    254: romdata_int <= 'hae3c;
    255: romdata_int <= 'h40e5;
    256: romdata_int <= 'h487; // Line Descriptor
    257: romdata_int <= 'h4307;
    258: romdata_int <= 'hb45;
    259: romdata_int <= 'h1029e;
    260: romdata_int <= 'h487; // Line Descriptor
    261: romdata_int <= 'h8e34;
    262: romdata_int <= 'hf351;
    263: romdata_int <= 'h9c6f;
    264: romdata_int <= 'h487; // Line Descriptor
    265: romdata_int <= 'hd228;
    266: romdata_int <= 'h45;
    267: romdata_int <= 'h4ca2;
    268: romdata_int <= 'h487; // Line Descriptor
    269: romdata_int <= 'h30b;
    270: romdata_int <= 'hdaf3;
    271: romdata_int <= 'hb657;
    272: romdata_int <= 'h487; // Line Descriptor
    273: romdata_int <= 'h1c36;
    274: romdata_int <= 'hb926;
    275: romdata_int <= 'hd4f9;
    276: romdata_int <= 'h487; // Line Descriptor
    277: romdata_int <= 'h3c7d;
    278: romdata_int <= 'hfedd;
    279: romdata_int <= 'h2860;
    280: romdata_int <= 'h487; // Line Descriptor
    281: romdata_int <= 'hca52;
    282: romdata_int <= 'ha8af;
    283: romdata_int <= 'h64a6;
    284: romdata_int <= 'h487; // Line Descriptor
    285: romdata_int <= 'he8ff;
    286: romdata_int <= 'ha449;
    287: romdata_int <= 'hab49;
    288: romdata_int <= 'h487; // Line Descriptor
    289: romdata_int <= 'h10467;
    290: romdata_int <= 'h855e;
    291: romdata_int <= 'h5041;
    292: romdata_int <= 'h487; // Line Descriptor
    293: romdata_int <= 'h906f;
    294: romdata_int <= 'hf550;
    295: romdata_int <= 'h34b5;
    296: romdata_int <= 'h487; // Line Descriptor
    297: romdata_int <= 'h10e2;
    298: romdata_int <= 'h2d11;
    299: romdata_int <= 'h8a06;
    300: romdata_int <= 'h487; // Line Descriptor
    301: romdata_int <= 'h2e38;
    302: romdata_int <= 'h10c62;
    303: romdata_int <= 'h40b4;
    304: romdata_int <= 'h487; // Line Descriptor
    305: romdata_int <= 'h5603;
    306: romdata_int <= 'h70c8;
    307: romdata_int <= 'hb822;
    308: romdata_int <= 'h487; // Line Descriptor
    309: romdata_int <= 'h8859;
    310: romdata_int <= 'h74e8;
    311: romdata_int <= 'h8ca0;
    312: romdata_int <= 'h487; // Line Descriptor
    313: romdata_int <= 'h9e08;
    314: romdata_int <= 'h9885;
    315: romdata_int <= 'h7a10;
    316: romdata_int <= 'h487; // Line Descriptor
    317: romdata_int <= 'h247e;
    318: romdata_int <= 'hd31e;
    319: romdata_int <= 'h4645;
    320: romdata_int <= 'h487; // Line Descriptor
    321: romdata_int <= 'h7e80;
    322: romdata_int <= 'hbeb5;
    323: romdata_int <= 'h12db;
    324: romdata_int <= 'h487; // Line Descriptor
    325: romdata_int <= 'hbb55;
    326: romdata_int <= 'hf8e5;
    327: romdata_int <= 'h1af3;
    328: romdata_int <= 'h487; // Line Descriptor
    329: romdata_int <= 'hf696;
    330: romdata_int <= 'he111;
    331: romdata_int <= 'hf087;
    332: romdata_int <= 'h587; // Line Descriptor
    333: romdata_int <= 'hdd59;
    334: romdata_int <= 'hcc98;
    335: romdata_int <= 'h2f3;
    336: romdata_int <= 'h1678; // Line Descriptor
    337: romdata_int <= 'hcf22;
    338: romdata_int <= 'h5eae;
    339: romdata_int <= 'h6b0b;
    340: romdata_int <= 'hb808;
    341: romdata_int <= 'h66d5;
    342: romdata_int <= 'h1a86;
    343: romdata_int <= 'h1c89;
    344: romdata_int <= 'h2e;
    345: romdata_int <= 'h3404;
    346: romdata_int <= 'h9f37;
    347: romdata_int <= 'h4c9a;
    348: romdata_int <= 'hb0;
    349: romdata_int <= 'h1678; // Line Descriptor
    350: romdata_int <= 'he860;
    351: romdata_int <= 'h9479;
    352: romdata_int <= 'h9cb8;
    353: romdata_int <= 'h67b;
    354: romdata_int <= 'hba7f;
    355: romdata_int <= 'hec38;
    356: romdata_int <= 'h2cb9;
    357: romdata_int <= 'h713b;
    358: romdata_int <= 'hd27c;
    359: romdata_int <= 'ha302;
    360: romdata_int <= 'hd09b;
    361: romdata_int <= 'h3d12;
    362: romdata_int <= 'h1678; // Line Descriptor
    363: romdata_int <= 'h6291;
    364: romdata_int <= 'hd20d;
    365: romdata_int <= 'hef28;
    366: romdata_int <= 'h808a;
    367: romdata_int <= 'h366b;
    368: romdata_int <= 'hb267;
    369: romdata_int <= 'h5255;
    370: romdata_int <= 'h1461;
    371: romdata_int <= 'h7cd5;
    372: romdata_int <= 'h691e;
    373: romdata_int <= 'h9ca5;
    374: romdata_int <= 'h1ce0;
    375: romdata_int <= 'h1678; // Line Descriptor
    376: romdata_int <= 'h96f3;
    377: romdata_int <= 'hc8a4;
    378: romdata_int <= 'h712c;
    379: romdata_int <= 'hb2a7;
    380: romdata_int <= 'hdaa6;
    381: romdata_int <= 'h722d;
    382: romdata_int <= 'hea43;
    383: romdata_int <= 'h4528;
    384: romdata_int <= 'heab0;
    385: romdata_int <= 'h2e42;
    386: romdata_int <= 'h9273;
    387: romdata_int <= 'hc87c;
    388: romdata_int <= 'h1678; // Line Descriptor
    389: romdata_int <= 'h9052;
    390: romdata_int <= 'h7e3b;
    391: romdata_int <= 'h3f2b;
    392: romdata_int <= 'h5664;
    393: romdata_int <= 'ha090;
    394: romdata_int <= 'h6b36;
    395: romdata_int <= 'h38d5;
    396: romdata_int <= 'h8662;
    397: romdata_int <= 'he0f2;
    398: romdata_int <= 'hc0b6;
    399: romdata_int <= 'hac9;
    400: romdata_int <= 'h8d54;
    401: romdata_int <= 'h1678; // Line Descriptor
    402: romdata_int <= 'h2b53;
    403: romdata_int <= 'h472c;
    404: romdata_int <= 'h9949;
    405: romdata_int <= 'hc67;
    406: romdata_int <= 'h34a6;
    407: romdata_int <= 'h40f2;
    408: romdata_int <= 'h5a88;
    409: romdata_int <= 'hbf27;
    410: romdata_int <= 'hcbd;
    411: romdata_int <= 'h845c;
    412: romdata_int <= 'he848;
    413: romdata_int <= 'h7f22;
    414: romdata_int <= 'h1678; // Line Descriptor
    415: romdata_int <= 'haa9f;
    416: romdata_int <= 'hcc82;
    417: romdata_int <= 'hc070;
    418: romdata_int <= 'h4d4f;
    419: romdata_int <= 'h3225;
    420: romdata_int <= 'h954d;
    421: romdata_int <= 'h3d52;
    422: romdata_int <= 'hc938;
    423: romdata_int <= 'h48f;
    424: romdata_int <= 'h400e;
    425: romdata_int <= 'h72ab;
    426: romdata_int <= 'hc475;
    427: romdata_int <= 'h1678; // Line Descriptor
    428: romdata_int <= 'h2505;
    429: romdata_int <= 'h2ca1;
    430: romdata_int <= 'h7a4d;
    431: romdata_int <= 'h1f48;
    432: romdata_int <= 'hb61a;
    433: romdata_int <= 'he80a;
    434: romdata_int <= 'h6316;
    435: romdata_int <= 'hdcee;
    436: romdata_int <= 'h5466;
    437: romdata_int <= 'hec32;
    438: romdata_int <= 'h98f3;
    439: romdata_int <= 'h372a;
    440: romdata_int <= 'h1678; // Line Descriptor
    441: romdata_int <= 'hd05f;
    442: romdata_int <= 'h34fe;
    443: romdata_int <= 'heca2;
    444: romdata_int <= 'h782a;
    445: romdata_int <= 'h88c9;
    446: romdata_int <= 'h24ce;
    447: romdata_int <= 'h4afd;
    448: romdata_int <= 'h6f19;
    449: romdata_int <= 'hc650;
    450: romdata_int <= 'hbe33;
    451: romdata_int <= 'h4a1c;
    452: romdata_int <= 'h1738;
    453: romdata_int <= 'h1678; // Line Descriptor
    454: romdata_int <= 'h1321;
    455: romdata_int <= 'hacc0;
    456: romdata_int <= 'h163f;
    457: romdata_int <= 'hc408;
    458: romdata_int <= 'he65;
    459: romdata_int <= 'h4ce5;
    460: romdata_int <= 'h30c0;
    461: romdata_int <= 'hd25d;
    462: romdata_int <= 'hd67b;
    463: romdata_int <= 'hb6fd;
    464: romdata_int <= 'hb2eb;
    465: romdata_int <= 'hac18;
    466: romdata_int <= 'h1678; // Line Descriptor
    467: romdata_int <= 'h2861;
    468: romdata_int <= 'hbc7f;
    469: romdata_int <= 'h868c;
    470: romdata_int <= 'h507e;
    471: romdata_int <= 'h7f3f;
    472: romdata_int <= 'h741f;
    473: romdata_int <= 'h8223;
    474: romdata_int <= 'h2746;
    475: romdata_int <= 'h1a90;
    476: romdata_int <= 'h8ada;
    477: romdata_int <= 'h963;
    478: romdata_int <= 'h5c70;
    479: romdata_int <= 'h1678; // Line Descriptor
    480: romdata_int <= 'h7306;
    481: romdata_int <= 'h5a0b;
    482: romdata_int <= 'h887b;
    483: romdata_int <= 'h1a3e;
    484: romdata_int <= 'h8cdb;
    485: romdata_int <= 'h8558;
    486: romdata_int <= 'ha6ee;
    487: romdata_int <= 'h2ac3;
    488: romdata_int <= 'h9445;
    489: romdata_int <= 'h6e87;
    490: romdata_int <= 'h1e5c;
    491: romdata_int <= 'h4eca;
    492: romdata_int <= 'h1678; // Line Descriptor
    493: romdata_int <= 'hae82;
    494: romdata_int <= 'hd667;
    495: romdata_int <= 'hd473;
    496: romdata_int <= 'h6e2b;
    497: romdata_int <= 'h6158;
    498: romdata_int <= 'he6c5;
    499: romdata_int <= 'h50ad;
    500: romdata_int <= 'hae35;
    501: romdata_int <= 'h6442;
    502: romdata_int <= 'h5617;
    503: romdata_int <= 'h2d15;
    504: romdata_int <= 'h74c;
    505: romdata_int <= 'h1678; // Line Descriptor
    506: romdata_int <= 'ha62c;
    507: romdata_int <= 'h3abb;
    508: romdata_int <= 'h673d;
    509: romdata_int <= 'h22ed;
    510: romdata_int <= 'hc131;
    511: romdata_int <= 'h3f1f;
    512: romdata_int <= 'hc6c4;
    513: romdata_int <= 'h814;
    514: romdata_int <= 'hdac9;
    515: romdata_int <= 'he55b;
    516: romdata_int <= 'hc20a;
    517: romdata_int <= 'ha69a;
    518: romdata_int <= 'h1678; // Line Descriptor
    519: romdata_int <= 'h921e;
    520: romdata_int <= 'h8d45;
    521: romdata_int <= 'ha078;
    522: romdata_int <= 'h4efc;
    523: romdata_int <= 'h5738;
    524: romdata_int <= 'h283f;
    525: romdata_int <= 'heef5;
    526: romdata_int <= 'h4efe;
    527: romdata_int <= 'hdf4b;
    528: romdata_int <= 'hb8a8;
    529: romdata_int <= 'h1897;
    530: romdata_int <= 'hb4a6;
    531: romdata_int <= 'h1678; // Line Descriptor
    532: romdata_int <= 'h851e;
    533: romdata_int <= 'h683c;
    534: romdata_int <= 'h5ce5;
    535: romdata_int <= 'hdc6b;
    536: romdata_int <= 'h4639;
    537: romdata_int <= 'h7966;
    538: romdata_int <= 'hd07;
    539: romdata_int <= 'h8b45;
    540: romdata_int <= 'h329e;
    541: romdata_int <= 'h7a81;
    542: romdata_int <= 'h794d;
    543: romdata_int <= 'h468b;
    544: romdata_int <= 'h1678; // Line Descriptor
    545: romdata_int <= 'h520e;
    546: romdata_int <= 'h1937;
    547: romdata_int <= 'he34c;
    548: romdata_int <= 'h3c91;
    549: romdata_int <= 'hbd0b;
    550: romdata_int <= 'h4f3;
    551: romdata_int <= 'h6457;
    552: romdata_int <= 'h166c;
    553: romdata_int <= 'h2aee;
    554: romdata_int <= 'h66f4;
    555: romdata_int <= 'h1236;
    556: romdata_int <= 'hcf26;
    557: romdata_int <= 'h1678; // Line Descriptor
    558: romdata_int <= 'h2006;
    559: romdata_int <= 'h7c3a;
    560: romdata_int <= 'hdb60;
    561: romdata_int <= 'h2e49;
    562: romdata_int <= 'h5e38;
    563: romdata_int <= 'hde62;
    564: romdata_int <= 'h96b4;
    565: romdata_int <= 'ha56;
    566: romdata_int <= 'h3860;
    567: romdata_int <= 'h74d8;
    568: romdata_int <= 'h8e03;
    569: romdata_int <= 'haac8;
    570: romdata_int <= 'h1678; // Line Descriptor
    571: romdata_int <= 'ha10;
    572: romdata_int <= 'h5458;
    573: romdata_int <= 'h32ee;
    574: romdata_int <= 'h6465;
    575: romdata_int <= 'h487e;
    576: romdata_int <= 'ha91e;
    577: romdata_int <= 'h8e45;
    578: romdata_int <= 'h926e;
    579: romdata_int <= 'h60a8;
    580: romdata_int <= 'h5030;
    581: romdata_int <= 'he80;
    582: romdata_int <= 'h58b5;
    583: romdata_int <= 'h1678; // Line Descriptor
    584: romdata_int <= 'h9e87;
    585: romdata_int <= 'h413b;
    586: romdata_int <= 'he121;
    587: romdata_int <= 'h14b1;
    588: romdata_int <= 'he11c;
    589: romdata_int <= 'hac3d;
    590: romdata_int <= 'hb159;
    591: romdata_int <= 'hd498;
    592: romdata_int <= 'h86f3;
    593: romdata_int <= 'haed9;
    594: romdata_int <= 'h6ad4;
    595: romdata_int <= 'hb03a;
    596: romdata_int <= 'h478; // Line Descriptor
    597: romdata_int <= 'hd94c;
    598: romdata_int <= 'h3aeb;
    599: romdata_int <= 'h76cf;
    600: romdata_int <= 'h478; // Line Descriptor
    601: romdata_int <= 'h1091;
    602: romdata_int <= 'he476;
    603: romdata_int <= 'he344;
    604: romdata_int <= 'h478; // Line Descriptor
    605: romdata_int <= 'h1d43;
    606: romdata_int <= 'h1085;
    607: romdata_int <= 'h26ed;
    608: romdata_int <= 'h478; // Line Descriptor
    609: romdata_int <= 'h959;
    610: romdata_int <= 'h12e3;
    611: romdata_int <= 'h82e4;
    612: romdata_int <= 'h478; // Line Descriptor
    613: romdata_int <= 'h8b57;
    614: romdata_int <= 'ha432;
    615: romdata_int <= 'h4567;
    616: romdata_int <= 'h478; // Line Descriptor
    617: romdata_int <= 'h4a74;
    618: romdata_int <= 'h7629;
    619: romdata_int <= 'hbd52;
    620: romdata_int <= 'h478; // Line Descriptor
    621: romdata_int <= 'hba19;
    622: romdata_int <= 'h9c1c;
    623: romdata_int <= 'h9123;
    624: romdata_int <= 'h478; // Line Descriptor
    625: romdata_int <= 'h51c;
    626: romdata_int <= 'h6833;
    627: romdata_int <= 'ha0ef;
    628: romdata_int <= 'h478; // Line Descriptor
    629: romdata_int <= 'hb55f;
    630: romdata_int <= 'h7b1c;
    631: romdata_int <= 'hcb55;
    632: romdata_int <= 'h478; // Line Descriptor
    633: romdata_int <= 'h827a;
    634: romdata_int <= 'h2e94;
    635: romdata_int <= 'h6c54;
    636: romdata_int <= 'h478; // Line Descriptor
    637: romdata_int <= 'he75b;
    638: romdata_int <= 'h594c;
    639: romdata_int <= 'hbabd;
    640: romdata_int <= 'h478; // Line Descriptor
    641: romdata_int <= 'hbe79;
    642: romdata_int <= 'he281;
    643: romdata_int <= 'ha40d;
    644: romdata_int <= 'h478; // Line Descriptor
    645: romdata_int <= 'h8ef2;
    646: romdata_int <= 'hcb34;
    647: romdata_int <= 'h294c;
    648: romdata_int <= 'h478; // Line Descriptor
    649: romdata_int <= 'hc64f;
    650: romdata_int <= 'h9117;
    651: romdata_int <= 'h4205;
    652: romdata_int <= 'h478; // Line Descriptor
    653: romdata_int <= 'hde6b;
    654: romdata_int <= 'h22b0;
    655: romdata_int <= 'h114a;
    656: romdata_int <= 'h478; // Line Descriptor
    657: romdata_int <= 'ha93e;
    658: romdata_int <= 'h2e4;
    659: romdata_int <= 'h22f5;
    660: romdata_int <= 'h478; // Line Descriptor
    661: romdata_int <= 'h7618;
    662: romdata_int <= 'hb854;
    663: romdata_int <= 'hef2f;
    664: romdata_int <= 'h478; // Line Descriptor
    665: romdata_int <= 'h6cf2;
    666: romdata_int <= 'h9a2c;
    667: romdata_int <= 'h30a0;
    668: romdata_int <= 'h478; // Line Descriptor
    669: romdata_int <= 'ha44f;
    670: romdata_int <= 'h98cb;
    671: romdata_int <= 'h9aee;
    672: romdata_int <= 'h478; // Line Descriptor
    673: romdata_int <= 'hc34e;
    674: romdata_int <= 'h5c13;
    675: romdata_int <= 'h8070;
    676: romdata_int <= 'h478; // Line Descriptor
    677: romdata_int <= 'he438;
    678: romdata_int <= 'hceb3;
    679: romdata_int <= 'h4962;
    680: romdata_int <= 'h478; // Line Descriptor
    681: romdata_int <= 'hb752;
    682: romdata_int <= 'hb564;
    683: romdata_int <= 'h3ad6;
    684: romdata_int <= 'h478; // Line Descriptor
    685: romdata_int <= 'heb06;
    686: romdata_int <= 'hc50b;
    687: romdata_int <= 'hcd3d;
    688: romdata_int <= 'h478; // Line Descriptor
    689: romdata_int <= 'h309b;
    690: romdata_int <= 'hd75c;
    691: romdata_int <= 'h7147;
    692: romdata_int <= 'h478; // Line Descriptor
    693: romdata_int <= 'h139;
    694: romdata_int <= 'h1e77;
    695: romdata_int <= 'h5a87;
    696: romdata_int <= 'h478; // Line Descriptor
    697: romdata_int <= 'hca38;
    698: romdata_int <= 'h9eb4;
    699: romdata_int <= 'h1507;
    700: romdata_int <= 'h478; // Line Descriptor
    701: romdata_int <= 'h26d3;
    702: romdata_int <= 'h6d1;
    703: romdata_int <= 'h2b8;
    704: romdata_int <= 'h478; // Line Descriptor
    705: romdata_int <= 'he43;
    706: romdata_int <= 'hc205;
    707: romdata_int <= 'hd925;
    708: romdata_int <= 'h478; // Line Descriptor
    709: romdata_int <= 'h5852;
    710: romdata_int <= 'h428e;
    711: romdata_int <= 'h96a6;
    712: romdata_int <= 'h478; // Line Descriptor
    713: romdata_int <= 'hb0df;
    714: romdata_int <= 'hab25;
    715: romdata_int <= 'hdc45;
    716: romdata_int <= 'h478; // Line Descriptor
    717: romdata_int <= 'h749b;
    718: romdata_int <= 'h6c86;
    719: romdata_int <= 'h5e7b;
    720: romdata_int <= 'h478; // Line Descriptor
    721: romdata_int <= 'ha265;
    722: romdata_int <= 'h8112;
    723: romdata_int <= 'he629;
    724: romdata_int <= 'h478; // Line Descriptor
    725: romdata_int <= 'h48d2;
    726: romdata_int <= 'h200a;
    727: romdata_int <= 'hd544;
    728: romdata_int <= 'h478; // Line Descriptor
    729: romdata_int <= 'h4566;
    730: romdata_int <= 'h7cce;
    731: romdata_int <= 'h5248;
    732: romdata_int <= 'h478; // Line Descriptor
    733: romdata_int <= 'h2ec;
    734: romdata_int <= 'h1829;
    735: romdata_int <= 'h631d;
    736: romdata_int <= 'h478; // Line Descriptor
    737: romdata_int <= 'h3622;
    738: romdata_int <= 'hccf4;
    739: romdata_int <= 'ha90b;
    740: romdata_int <= 'h478; // Line Descriptor
    741: romdata_int <= 'h9ab8;
    742: romdata_int <= 'hd015;
    743: romdata_int <= 'h8878;
    744: romdata_int <= 'h478; // Line Descriptor
    745: romdata_int <= 'h3943;
    746: romdata_int <= 'ha2e1;
    747: romdata_int <= 'h2042;
    748: romdata_int <= 'h478; // Line Descriptor
    749: romdata_int <= 'h6024;
    750: romdata_int <= 'hd8d9;
    751: romdata_int <= 'h2458;
    752: romdata_int <= 'h578; // Line Descriptor
    753: romdata_int <= 'h42d3;
    754: romdata_int <= 'h5422;
    755: romdata_int <= 'h3f4b;
    756: romdata_int <= 'h166c; // Line Descriptor
    757: romdata_int <= 'hbb22;
    758: romdata_int <= 'h54ae;
    759: romdata_int <= 'h610b;
    760: romdata_int <= 'ha608;
    761: romdata_int <= 'h5cd5;
    762: romdata_int <= 'h1886;
    763: romdata_int <= 'h1a89;
    764: romdata_int <= 'h2e;
    765: romdata_int <= 'h2e04;
    766: romdata_int <= 'h8f37;
    767: romdata_int <= 'h449a;
    768: romdata_int <= 'hb0;
    769: romdata_int <= 'h166c; // Line Descriptor
    770: romdata_int <= 'hd079;
    771: romdata_int <= 'h86b8;
    772: romdata_int <= 'h8c7b;
    773: romdata_int <= 'h67f;
    774: romdata_int <= 'ha838;
    775: romdata_int <= 'hd4b9;
    776: romdata_int <= 'h293b;
    777: romdata_int <= 'h647c;
    778: romdata_int <= 'hbd02;
    779: romdata_int <= 'h929b;
    780: romdata_int <= 'h3712;
    781: romdata_int <= 'h3a99;
    782: romdata_int <= 'h166c; // Line Descriptor
    783: romdata_int <= 'hbe0d;
    784: romdata_int <= 'hd728;
    785: romdata_int <= 'h748a;
    786: romdata_int <= 'h2c6b;
    787: romdata_int <= 'ha067;
    788: romdata_int <= 'h4a55;
    789: romdata_int <= 'h1261;
    790: romdata_int <= 'h74d5;
    791: romdata_int <= 'h611e;
    792: romdata_int <= 'h90a5;
    793: romdata_int <= 'h18e0;
    794: romdata_int <= 'h5ae6;
    795: romdata_int <= 'h166c; // Line Descriptor
    796: romdata_int <= 'hb52c;
    797: romdata_int <= 'h64a7;
    798: romdata_int <= 'h9ea6;
    799: romdata_int <= 'hc22d;
    800: romdata_int <= 'h6243;
    801: romdata_int <= 'hd328;
    802: romdata_int <= 'h3cb0;
    803: romdata_int <= 'h3042;
    804: romdata_int <= 'h8473;
    805: romdata_int <= 'hb67c;
    806: romdata_int <= 'h98e5;
    807: romdata_int <= 'h66c9;
    808: romdata_int <= 'h166c; // Line Descriptor
    809: romdata_int <= 'h3b2b;
    810: romdata_int <= 'h4e64;
    811: romdata_int <= 'h8890;
    812: romdata_int <= 'h5336;
    813: romdata_int <= 'h34d5;
    814: romdata_int <= 'h7c62;
    815: romdata_int <= 'hc8f2;
    816: romdata_int <= 'hb0b6;
    817: romdata_int <= 'hac9;
    818: romdata_int <= 'h8154;
    819: romdata_int <= 'h304a;
    820: romdata_int <= 'h2277;
    821: romdata_int <= 'h166c; // Line Descriptor
    822: romdata_int <= 'h8349;
    823: romdata_int <= 'ha67;
    824: romdata_int <= 'h28a6;
    825: romdata_int <= 'h30f2;
    826: romdata_int <= 'h5288;
    827: romdata_int <= 'ha727;
    828: romdata_int <= 'h8bd;
    829: romdata_int <= 'h805c;
    830: romdata_int <= 'hd448;
    831: romdata_int <= 'h7922;
    832: romdata_int <= 'hcd01;
    833: romdata_int <= 'hb934;
    834: romdata_int <= 'h166c; // Line Descriptor
    835: romdata_int <= 'haa82;
    836: romdata_int <= 'h4670;
    837: romdata_int <= 'h274f;
    838: romdata_int <= 'h7c25;
    839: romdata_int <= 'h394d;
    840: romdata_int <= 'hb552;
    841: romdata_int <= 'h538;
    842: romdata_int <= 'h3e8f;
    843: romdata_int <= 'h6c0e;
    844: romdata_int <= 'h3cab;
    845: romdata_int <= 'hb275;
    846: romdata_int <= 'h5e41;
    847: romdata_int <= 'h166c; // Line Descriptor
    848: romdata_int <= 'h24a1;
    849: romdata_int <= 'h704d;
    850: romdata_int <= 'h1b48;
    851: romdata_int <= 'ha01a;
    852: romdata_int <= 'hd00a;
    853: romdata_int <= 'h5916;
    854: romdata_int <= 'hc4ee;
    855: romdata_int <= 'h5066;
    856: romdata_int <= 'hd632;
    857: romdata_int <= 'h8af3;
    858: romdata_int <= 'h2b2a;
    859: romdata_int <= 'ha158;
    860: romdata_int <= 'h166c; // Line Descriptor
    861: romdata_int <= 'h348d;
    862: romdata_int <= 'h9231;
    863: romdata_int <= 'h38a0;
    864: romdata_int <= 'h6ed0;
    865: romdata_int <= 'h2344;
    866: romdata_int <= 'h8c06;
    867: romdata_int <= 'h7030;
    868: romdata_int <= 'h4c9b;
    869: romdata_int <= 'h26d6;
    870: romdata_int <= 'h10df;
    871: romdata_int <= 'h86be;
    872: romdata_int <= 'h1b35;
    873: romdata_int <= 'h166c; // Line Descriptor
    874: romdata_int <= 'h2efe;
    875: romdata_int <= 'hd4a2;
    876: romdata_int <= 'h6c2a;
    877: romdata_int <= 'h76c9;
    878: romdata_int <= 'h24ce;
    879: romdata_int <= 'h42fd;
    880: romdata_int <= 'h6919;
    881: romdata_int <= 'hb850;
    882: romdata_int <= 'hb033;
    883: romdata_int <= 'h481c;
    884: romdata_int <= 'hf38;
    885: romdata_int <= 'h4021;
    886: romdata_int <= 'h166c; // Line Descriptor
    887: romdata_int <= 'h9c3f;
    888: romdata_int <= 'h1208;
    889: romdata_int <= 'hb265;
    890: romdata_int <= 'hce5;
    891: romdata_int <= 'h44c0;
    892: romdata_int <= 'h2e5d;
    893: romdata_int <= 'hbe7b;
    894: romdata_int <= 'haafd;
    895: romdata_int <= 'ha6eb;
    896: romdata_int <= 'ha218;
    897: romdata_int <= 'hac40;
    898: romdata_int <= 'h7522;
    899: romdata_int <= 'h166c; // Line Descriptor
    900: romdata_int <= 'h7a8c;
    901: romdata_int <= 'h4a7e;
    902: romdata_int <= 'h633f;
    903: romdata_int <= 'h5a1f;
    904: romdata_int <= 'h7823;
    905: romdata_int <= 'h2746;
    906: romdata_int <= 'h1490;
    907: romdata_int <= 'h8eda;
    908: romdata_int <= 'h563;
    909: romdata_int <= 'h5670;
    910: romdata_int <= 'h3eb4;
    911: romdata_int <= 'h4e8f;
    912: romdata_int <= 'h166c; // Line Descriptor
    913: romdata_int <= 'h847b;
    914: romdata_int <= 'h163e;
    915: romdata_int <= 'h72db;
    916: romdata_int <= 'h6958;
    917: romdata_int <= 'h94ee;
    918: romdata_int <= 'h2cc3;
    919: romdata_int <= 'h7645;
    920: romdata_int <= 'h1087;
    921: romdata_int <= 'h945c;
    922: romdata_int <= 'h4cca;
    923: romdata_int <= 'h9f06;
    924: romdata_int <= 'h737;
    925: romdata_int <= 'h166c; // Line Descriptor
    926: romdata_int <= 'hbc73;
    927: romdata_int <= 'h662b;
    928: romdata_int <= 'h4d58;
    929: romdata_int <= 'hcec5;
    930: romdata_int <= 'h4ead;
    931: romdata_int <= 'h9c35;
    932: romdata_int <= 'h6c42;
    933: romdata_int <= 'h5a17;
    934: romdata_int <= 'h2915;
    935: romdata_int <= 'h94c;
    936: romdata_int <= 'h5506;
    937: romdata_int <= 'h4664;
    938: romdata_int <= 'h166c; // Line Descriptor
    939: romdata_int <= 'h5f3d;
    940: romdata_int <= 'h1ced;
    941: romdata_int <= 'had31;
    942: romdata_int <= 'h2b1f;
    943: romdata_int <= 'hb6c4;
    944: romdata_int <= 'ha14;
    945: romdata_int <= 'hc6c9;
    946: romdata_int <= 'hcd5b;
    947: romdata_int <= 'hbe0a;
    948: romdata_int <= 'h9c9a;
    949: romdata_int <= 'h1ecb;
    950: romdata_int <= 'h7b1d;
    951: romdata_int <= 'h166c; // Line Descriptor
    952: romdata_int <= 'h98fc;
    953: romdata_int <= 'h4538;
    954: romdata_int <= 'h403f;
    955: romdata_int <= 'h20f5;
    956: romdata_int <= 'hd6fe;
    957: romdata_int <= 'h494b;
    958: romdata_int <= 'hcaa8;
    959: romdata_int <= 'hac97;
    960: romdata_int <= 'h16a6;
    961: romdata_int <= 'hb4d5;
    962: romdata_int <= 'hc8b1;
    963: romdata_int <= 'h58a1;
    964: romdata_int <= 'h166c; // Line Descriptor
    965: romdata_int <= 'hc66b;
    966: romdata_int <= 'h3639;
    967: romdata_int <= 'h5966;
    968: romdata_int <= 'h907;
    969: romdata_int <= 'h7345;
    970: romdata_int <= 'h329e;
    971: romdata_int <= 'h8481;
    972: romdata_int <= 'h834d;
    973: romdata_int <= 'h508b;
    974: romdata_int <= 'hba99;
    975: romdata_int <= 'h2c34;
    976: romdata_int <= 'h8951;
    977: romdata_int <= 'h166c; // Line Descriptor
    978: romdata_int <= 'h4291;
    979: romdata_int <= 'haf0b;
    980: romdata_int <= 'h2f3;
    981: romdata_int <= 'h4857;
    982: romdata_int <= 'h166c;
    983: romdata_int <= 'h20ee;
    984: romdata_int <= 'h6af4;
    985: romdata_int <= 'hc36;
    986: romdata_int <= 'hc726;
    987: romdata_int <= 'hcf9;
    988: romdata_int <= 'hc44a;
    989: romdata_int <= 'hcb56;
    990: romdata_int <= 'h166c; // Line Descriptor
    991: romdata_int <= 'h14e2;
    992: romdata_int <= 'h56ff;
    993: romdata_int <= 'h9649;
    994: romdata_int <= 'h3d49;
    995: romdata_int <= 'h9f5d;
    996: romdata_int <= 'h90a4;
    997: romdata_int <= 'h5469;
    998: romdata_int <= 'h4067;
    999: romdata_int <= 'h6f5e;
    1000: romdata_int <= 'h6a41;
    1001: romdata_int <= 'haac8;
    1002: romdata_int <= 'h7f3f;
    1003: romdata_int <= 'h166c; // Line Descriptor
    1004: romdata_int <= 'h8a65;
    1005: romdata_int <= 'h327e;
    1006: romdata_int <= 'ha31e;
    1007: romdata_int <= 'h8045;
    1008: romdata_int <= 'h7e6e;
    1009: romdata_int <= 'h6ea8;
    1010: romdata_int <= 'h5e30;
    1011: romdata_int <= 'h280;
    1012: romdata_int <= 'h52b5;
    1013: romdata_int <= 'h12db;
    1014: romdata_int <= 'h3467;
    1015: romdata_int <= 'h8d49;
    1016: romdata_int <= 'h166c; // Line Descriptor
    1017: romdata_int <= 'h10b1;
    1018: romdata_int <= 'hcd1c;
    1019: romdata_int <= 'ha43d;
    1020: romdata_int <= 'ha959;
    1021: romdata_int <= 'hbc98;
    1022: romdata_int <= 'h92f3;
    1023: romdata_int <= 'ha4d9;
    1024: romdata_int <= 'h7ad4;
    1025: romdata_int <= 'ha83a;
    1026: romdata_int <= 'h633b;
    1027: romdata_int <= 'hc251;
    1028: romdata_int <= 'haeba;
    1029: romdata_int <= 'h166c; // Line Descriptor
    1030: romdata_int <= 'hcb43;
    1031: romdata_int <= 'h9a85;
    1032: romdata_int <= 'h90ed;
    1033: romdata_int <= 'h1826;
    1034: romdata_int <= 'hce1b;
    1035: romdata_int <= 'hc2c2;
    1036: romdata_int <= 'h6159;
    1037: romdata_int <= 'h46e3;
    1038: romdata_int <= 'hcee4;
    1039: romdata_int <= 'h20ba;
    1040: romdata_int <= 'h14e6;
    1041: romdata_int <= 'h2470;
    1042: romdata_int <= 'h166c; // Line Descriptor
    1043: romdata_int <= 'h7f61;
    1044: romdata_int <= 'h1f08;
    1045: romdata_int <= 'h5079;
    1046: romdata_int <= 'h6a81;
    1047: romdata_int <= 'h2a0d;
    1048: romdata_int <= 'hbac6;
    1049: romdata_int <= 'h371d;
    1050: romdata_int <= 'ha24f;
    1051: romdata_int <= 'hd2f2;
    1052: romdata_int <= 'hd134;
    1053: romdata_int <= 'h734c;
    1054: romdata_int <= 'h9b2c;
    1055: romdata_int <= 'h166c; // Line Descriptor
    1056: romdata_int <= 'h8e36;
    1057: romdata_int <= 'h5d3e;
    1058: romdata_int <= 'h22e4;
    1059: romdata_int <= 'hc0f5;
    1060: romdata_int <= 'h6d5;
    1061: romdata_int <= 'hb2fc;
    1062: romdata_int <= 'h1f62;
    1063: romdata_int <= 'h3a18;
    1064: romdata_int <= 'h6454;
    1065: romdata_int <= 'ha52f;
    1066: romdata_int <= 'h7cc7;
    1067: romdata_int <= 'h2ad;
    1068: romdata_int <= 'h46c; // Line Descriptor
    1069: romdata_int <= 'hea0;
    1070: romdata_int <= 'h98fc;
    1071: romdata_int <= 'h32b0;
    1072: romdata_int <= 'h46c; // Line Descriptor
    1073: romdata_int <= 'hb8ee;
    1074: romdata_int <= 'h5726;
    1075: romdata_int <= 'h7070;
    1076: romdata_int <= 'h46c; // Line Descriptor
    1077: romdata_int <= 'hb070;
    1078: romdata_int <= 'hc144;
    1079: romdata_int <= 'h1d21;
    1080: romdata_int <= 'h46c; // Line Descriptor
    1081: romdata_int <= 'h3f62;
    1082: romdata_int <= 'h1d35;
    1083: romdata_int <= 'h68e6;
    1084: romdata_int <= 'h46c; // Line Descriptor
    1085: romdata_int <= 'h4d6;
    1086: romdata_int <= 'haf5f;
    1087: romdata_int <= 'hc113;
    1088: romdata_int <= 'h46c; // Line Descriptor
    1089: romdata_int <= 'hc93d;
    1090: romdata_int <= 'h9661;
    1091: romdata_int <= 'h834f;
    1092: romdata_int <= 'h46c; // Line Descriptor
    1093: romdata_int <= 'hb747;
    1094: romdata_int <= 'h8601;
    1095: romdata_int <= 'h9642;
    1096: romdata_int <= 'h46c; // Line Descriptor
    1097: romdata_int <= 'h9487;
    1098: romdata_int <= 'h9b61;
    1099: romdata_int <= 'h42d1;
    1100: romdata_int <= 'h46c; // Line Descriptor
    1101: romdata_int <= 'h107;
    1102: romdata_int <= 'he3d;
    1103: romdata_int <= 'h5c09;
    1104: romdata_int <= 'h46c; // Line Descriptor
    1105: romdata_int <= 'h78b8;
    1106: romdata_int <= 'h8820;
    1107: romdata_int <= 'h4b0f;
    1108: romdata_int <= 'h46c; // Line Descriptor
    1109: romdata_int <= 'hd325;
    1110: romdata_int <= 'h66bb;
    1111: romdata_int <= 'h384b;
    1112: romdata_int <= 'h46c; // Line Descriptor
    1113: romdata_int <= 'hc4a6;
    1114: romdata_int <= 'h8b50;
    1115: romdata_int <= 'h76f7;
    1116: romdata_int <= 'h46c; // Line Descriptor
    1117: romdata_int <= 'hb645;
    1118: romdata_int <= 'h8713;
    1119: romdata_int <= 'hb07d;
    1120: romdata_int <= 'h46c; // Line Descriptor
    1121: romdata_int <= 'h627b;
    1122: romdata_int <= 'h5af0;
    1123: romdata_int <= 'h4e4e;
    1124: romdata_int <= 'h46c; // Line Descriptor
    1125: romdata_int <= 'h4086;
    1126: romdata_int <= 'h9954;
    1127: romdata_int <= 'h6cb6;
    1128: romdata_int <= 'h46c; // Line Descriptor
    1129: romdata_int <= 'hc829;
    1130: romdata_int <= 'h36ea;
    1131: romdata_int <= 'ha443;
    1132: romdata_int <= 'h46c; // Line Descriptor
    1133: romdata_int <= 'hc744;
    1134: romdata_int <= 'h7cec;
    1135: romdata_int <= 'h489;
    1136: romdata_int <= 'h46c; // Line Descriptor
    1137: romdata_int <= 'h6048;
    1138: romdata_int <= 'hd601;
    1139: romdata_int <= 'h780b;
    1140: romdata_int <= 'h46c; // Line Descriptor
    1141: romdata_int <= 'h891d;
    1142: romdata_int <= 'h8c31;
    1143: romdata_int <= 'h16a0;
    1144: romdata_int <= 'h46c; // Line Descriptor
    1145: romdata_int <= 'hc10b;
    1146: romdata_int <= 'h1318;
    1147: romdata_int <= 'h92fa;
    1148: romdata_int <= 'h46c; // Line Descriptor
    1149: romdata_int <= 'hcc78;
    1150: romdata_int <= 'h6613;
    1151: romdata_int <= 'hc96;
    1152: romdata_int <= 'h46c; // Line Descriptor
    1153: romdata_int <= 'h242;
    1154: romdata_int <= 'hbd28;
    1155: romdata_int <= 'h80b5;
    1156: romdata_int <= 'h46c; // Line Descriptor
    1157: romdata_int <= 'h1058;
    1158: romdata_int <= 'h18cb;
    1159: romdata_int <= 'h7b67;
    1160: romdata_int <= 'h46c; // Line Descriptor
    1161: romdata_int <= 'hcb4b;
    1162: romdata_int <= 'h7538;
    1163: romdata_int <= 'h1cd9;
    1164: romdata_int <= 'h46c; // Line Descriptor
    1165: romdata_int <= 'h2aad;
    1166: romdata_int <= 'h4909;
    1167: romdata_int <= 'h96a7;
    1168: romdata_int <= 'h46c; // Line Descriptor
    1169: romdata_int <= 'h8ad2;
    1170: romdata_int <= 'h30fe;
    1171: romdata_int <= 'h72a;
    1172: romdata_int <= 'h46c; // Line Descriptor
    1173: romdata_int <= 'h5305;
    1174: romdata_int <= 'h5125;
    1175: romdata_int <= 'h3917;
    1176: romdata_int <= 'h46c; // Line Descriptor
    1177: romdata_int <= 'h828d;
    1178: romdata_int <= 'h764e;
    1179: romdata_int <= 'h3d03;
    1180: romdata_int <= 'h46c; // Line Descriptor
    1181: romdata_int <= 'ha889;
    1182: romdata_int <= 'h647b;
    1183: romdata_int <= 'h7074;
    1184: romdata_int <= 'h46c; // Line Descriptor
    1185: romdata_int <= 'h3509;
    1186: romdata_int <= 'h9417;
    1187: romdata_int <= 'h3eb6;
    1188: romdata_int <= 'h46c; // Line Descriptor
    1189: romdata_int <= 'hce39;
    1190: romdata_int <= 'h8e29;
    1191: romdata_int <= 'hb8f3;
    1192: romdata_int <= 'h46c; // Line Descriptor
    1193: romdata_int <= 'h906e;
    1194: romdata_int <= 'hb506;
    1195: romdata_int <= 'hb24d;
    1196: romdata_int <= 'h46c; // Line Descriptor
    1197: romdata_int <= 'h3262;
    1198: romdata_int <= 'hc208;
    1199: romdata_int <= 'h2c46;
    1200: romdata_int <= 'h46c; // Line Descriptor
    1201: romdata_int <= 'h6e60;
    1202: romdata_int <= 'h1e7a;
    1203: romdata_int <= 'h44f8;
    1204: romdata_int <= 'h46c; // Line Descriptor
    1205: romdata_int <= 'h5c93;
    1206: romdata_int <= 'h5553;
    1207: romdata_int <= 'h84c6;
    1208: romdata_int <= 'h46c; // Line Descriptor
    1209: romdata_int <= 'h2061;
    1210: romdata_int <= 'h280e;
    1211: romdata_int <= 'h220b;
    1212: romdata_int <= 'h46c; // Line Descriptor
    1213: romdata_int <= 'hbf1a;
    1214: romdata_int <= 'had51;
    1215: romdata_int <= 'h1acd;
    1216: romdata_int <= 'h46c; // Line Descriptor
    1217: romdata_int <= 'ha02f;
    1218: romdata_int <= 'hc468;
    1219: romdata_int <= 'hf3d;
    1220: romdata_int <= 'h46c; // Line Descriptor
    1221: romdata_int <= 'hd108;
    1222: romdata_int <= 'h6b47;
    1223: romdata_int <= 'h4c7b;
    1224: romdata_int <= 'h46c; // Line Descriptor
    1225: romdata_int <= 'hd452;
    1226: romdata_int <= 'ha20d;
    1227: romdata_int <= 'h24c4;
    1228: romdata_int <= 'h46c; // Line Descriptor
    1229: romdata_int <= 'hd2d9;
    1230: romdata_int <= 'h72a1;
    1231: romdata_int <= 'h3b49;
    1232: romdata_int <= 'h46c; // Line Descriptor
    1233: romdata_int <= 'hab32;
    1234: romdata_int <= 'h4a6b;
    1235: romdata_int <= 'h2eb8;
    1236: romdata_int <= 'h46c; // Line Descriptor
    1237: romdata_int <= 'hb3a;
    1238: romdata_int <= 'hae48;
    1239: romdata_int <= 'h7f37;
    1240: romdata_int <= 'h46c; // Line Descriptor
    1241: romdata_int <= 'ha6b9;
    1242: romdata_int <= 'h4706;
    1243: romdata_int <= 'h1463;
    1244: romdata_int <= 'h46c; // Line Descriptor
    1245: romdata_int <= 'h267a;
    1246: romdata_int <= 'h5ec3;
    1247: romdata_int <= 'h56ca;
    1248: romdata_int <= 'h46c; // Line Descriptor
    1249: romdata_int <= 'h5828;
    1250: romdata_int <= 'h4320;
    1251: romdata_int <= 'h682c;
    1252: romdata_int <= 'h46c; // Line Descriptor
    1253: romdata_int <= 'h9a33;
    1254: romdata_int <= 'hba12;
    1255: romdata_int <= 'h9c2c;
    1256: romdata_int <= 'h56c; // Line Descriptor
    1257: romdata_int <= 'h11c;
    1258: romdata_int <= 'h9e9c;
    1259: romdata_int <= 'h889;
    1260: romdata_int <= 'he5a; // Line Descriptor
    1261: romdata_int <= 'h6c00;
    1262: romdata_int <= 'h6067;
    1263: romdata_int <= 'ha49f;
    1264: romdata_int <= 'h2b32;
    1265: romdata_int <= 'hb32a;
    1266: romdata_int <= 'h6271;
    1267: romdata_int <= 'h1c1c;
    1268: romdata_int <= 'h5e5f;
    1269: romdata_int <= 'he5a; // Line Descriptor
    1270: romdata_int <= 'h7e50;
    1271: romdata_int <= 'h6e00;
    1272: romdata_int <= 'h5a33;
    1273: romdata_int <= 'h141c;
    1274: romdata_int <= 'h6538;
    1275: romdata_int <= 'h8d08;
    1276: romdata_int <= 'h6628;
    1277: romdata_int <= 'h7e21;
    1278: romdata_int <= 'he5a; // Line Descriptor
    1279: romdata_int <= 'h7000;
    1280: romdata_int <= 'h8f12;
    1281: romdata_int <= 'h706;
    1282: romdata_int <= 'h3521;
    1283: romdata_int <= 'h26c0;
    1284: romdata_int <= 'ha03f;
    1285: romdata_int <= 'h9008;
    1286: romdata_int <= 'h9e65;
    1287: romdata_int <= 'he5a; // Line Descriptor
    1288: romdata_int <= 'h7200;
    1289: romdata_int <= 'h6640;
    1290: romdata_int <= 'h6d22;
    1291: romdata_int <= 'h2ecf;
    1292: romdata_int <= 'h3e80;
    1293: romdata_int <= 'h72ab;
    1294: romdata_int <= 'ha98;
    1295: romdata_int <= 'h80b4;
    1296: romdata_int <= 'he5a; // Line Descriptor
    1297: romdata_int <= 'h7400;
    1298: romdata_int <= 'h148c;
    1299: romdata_int <= 'he7e;
    1300: romdata_int <= 'h753f;
    1301: romdata_int <= 'h41f;
    1302: romdata_int <= 'h3023;
    1303: romdata_int <= 'h3f46;
    1304: romdata_int <= 'h4a90;
    1305: romdata_int <= 'he5a; // Line Descriptor
    1306: romdata_int <= 'h7600;
    1307: romdata_int <= 'h62ba;
    1308: romdata_int <= 'hb0b1;
    1309: romdata_int <= 'h3aee;
    1310: romdata_int <= 'h5a44;
    1311: romdata_int <= 'h68eb;
    1312: romdata_int <= 'h14b0;
    1313: romdata_int <= 'h4823;
    1314: romdata_int <= 'he5a; // Line Descriptor
    1315: romdata_int <= 'h7800;
    1316: romdata_int <= 'h7158;
    1317: romdata_int <= 'h3aee;
    1318: romdata_int <= 'h88c3;
    1319: romdata_int <= 'h645;
    1320: romdata_int <= 'h2087;
    1321: romdata_int <= 'h6c5c;
    1322: romdata_int <= 'h40ca;
    1323: romdata_int <= 'he5a; // Line Descriptor
    1324: romdata_int <= 'h7a00;
    1325: romdata_int <= 'h84fd;
    1326: romdata_int <= 'ha69d;
    1327: romdata_int <= 'h9a7d;
    1328: romdata_int <= 'h5c41;
    1329: romdata_int <= 'hb007;
    1330: romdata_int <= 'h3682;
    1331: romdata_int <= 'h4c67;
    1332: romdata_int <= 'he5a; // Line Descriptor
    1333: romdata_int <= 'h7c00;
    1334: romdata_int <= 'h2a17;
    1335: romdata_int <= 'h1715;
    1336: romdata_int <= 'had4c;
    1337: romdata_int <= 'h6d06;
    1338: romdata_int <= 'h1a64;
    1339: romdata_int <= 'h22ad;
    1340: romdata_int <= 'h583c;
    1341: romdata_int <= 'he5a; // Line Descriptor
    1342: romdata_int <= 'h7e00;
    1343: romdata_int <= 'h86f6;
    1344: romdata_int <= 'h2e2c;
    1345: romdata_int <= 'h94bb;
    1346: romdata_int <= 'h93d;
    1347: romdata_int <= 'haaed;
    1348: romdata_int <= 'h9531;
    1349: romdata_int <= 'ha51f;
    1350: romdata_int <= 'he5a; // Line Descriptor
    1351: romdata_int <= 'h8000;
    1352: romdata_int <= 'h4b1d;
    1353: romdata_int <= 'h232;
    1354: romdata_int <= 'h6af6;
    1355: romdata_int <= 'haaa2;
    1356: romdata_int <= 'h4ca4;
    1357: romdata_int <= 'h60b3;
    1358: romdata_int <= 'h23d;
    1359: romdata_int <= 'he5a; // Line Descriptor
    1360: romdata_int <= 'h8200;
    1361: romdata_int <= 'h2832;
    1362: romdata_int <= 'ha8bd;
    1363: romdata_int <= 'haf03;
    1364: romdata_int <= 'h442f;
    1365: romdata_int <= 'h64f8;
    1366: romdata_int <= 'h2abc;
    1367: romdata_int <= 'h20ef;
    1368: romdata_int <= 'he5a; // Line Descriptor
    1369: romdata_int <= 'h8400;
    1370: romdata_int <= 'h6474;
    1371: romdata_int <= 'h7c44;
    1372: romdata_int <= 'h7967;
    1373: romdata_int <= 'h726a;
    1374: romdata_int <= 'h7b56;
    1375: romdata_int <= 'h4520;
    1376: romdata_int <= 'h7c1e;
    1377: romdata_int <= 'he5a; // Line Descriptor
    1378: romdata_int <= 'h8600;
    1379: romdata_int <= 'h8cf5;
    1380: romdata_int <= 'hafe;
    1381: romdata_int <= 'ha14b;
    1382: romdata_int <= 'h36a8;
    1383: romdata_int <= 'h9c97;
    1384: romdata_int <= 'h1ea6;
    1385: romdata_int <= 'h82d5;
    1386: romdata_int <= 'he5a; // Line Descriptor
    1387: romdata_int <= 'h8800;
    1388: romdata_int <= 'h3a4a;
    1389: romdata_int <= 'h60cc;
    1390: romdata_int <= 'h98cb;
    1391: romdata_int <= 'h246e;
    1392: romdata_int <= 'hd1e;
    1393: romdata_int <= 'h563c;
    1394: romdata_int <= 'h46e5;
    1395: romdata_int <= 'he5a; // Line Descriptor
    1396: romdata_int <= 'h8a00;
    1397: romdata_int <= 'h194d;
    1398: romdata_int <= 'h268b;
    1399: romdata_int <= 'hb099;
    1400: romdata_int <= 'h8434;
    1401: romdata_int <= 'h5151;
    1402: romdata_int <= 'h426f;
    1403: romdata_int <= 'h9d13;
    1404: romdata_int <= 'he5a; // Line Descriptor
    1405: romdata_int <= 'h8c00;
    1406: romdata_int <= 'h40e;
    1407: romdata_int <= 'h5537;
    1408: romdata_int <= 'h114c;
    1409: romdata_int <= 'h1a91;
    1410: romdata_int <= 'h70b;
    1411: romdata_int <= 'ha2f3;
    1412: romdata_int <= 'h4257;
    1413: romdata_int <= 'he5a; // Line Descriptor
    1414: romdata_int <= 'h8e00;
    1415: romdata_int <= 'h3049;
    1416: romdata_int <= 'h4149;
    1417: romdata_int <= 'h535d;
    1418: romdata_int <= 'h8ea4;
    1419: romdata_int <= 'h7669;
    1420: romdata_int <= 'h8267;
    1421: romdata_int <= 'h695e;
    1422: romdata_int <= 'he5a; // Line Descriptor
    1423: romdata_int <= 'h9000;
    1424: romdata_int <= 'h100f;
    1425: romdata_int <= 'h8047;
    1426: romdata_int <= 'h92b8;
    1427: romdata_int <= 'h1ce2;
    1428: romdata_int <= 'h3911;
    1429: romdata_int <= 'ha806;
    1430: romdata_int <= 'h5a3a;
    1431: romdata_int <= 'he5a; // Line Descriptor
    1432: romdata_int <= 'h9200;
    1433: romdata_int <= 'hb2d8;
    1434: romdata_int <= 'h3203;
    1435: romdata_int <= 'h16c8;
    1436: romdata_int <= 'h2822;
    1437: romdata_int <= 'h5894;
    1438: romdata_int <= 'h2c59;
    1439: romdata_int <= 'h2eaa;
    1440: romdata_int <= 'he5a; // Line Descriptor
    1441: romdata_int <= 'h9400;
    1442: romdata_int <= 'h1685;
    1443: romdata_int <= 'h8c10;
    1444: romdata_int <= 'h5058;
    1445: romdata_int <= 'h54ee;
    1446: romdata_int <= 'h4e65;
    1447: romdata_int <= 'h3c7e;
    1448: romdata_int <= 'h31e;
    1449: romdata_int <= 'he5a; // Line Descriptor
    1450: romdata_int <= 'h9600;
    1451: romdata_int <= 'hc67;
    1452: romdata_int <= 'h5d49;
    1453: romdata_int <= 'h5632;
    1454: romdata_int <= 'h1355;
    1455: romdata_int <= 'h48e5;
    1456: romdata_int <= 'h66f3;
    1457: romdata_int <= 'h7937;
    1458: romdata_int <= 'he5a; // Line Descriptor
    1459: romdata_int <= 'h9800;
    1460: romdata_int <= 'h5ab1;
    1461: romdata_int <= 'h951c;
    1462: romdata_int <= 'h3c3d;
    1463: romdata_int <= 'h8b59;
    1464: romdata_int <= 'h4698;
    1465: romdata_int <= 'h9ef3;
    1466: romdata_int <= 'h96d9;
    1467: romdata_int <= 'he5a; // Line Descriptor
    1468: romdata_int <= 'h9a00;
    1469: romdata_int <= 'h74cf;
    1470: romdata_int <= 'h2433;
    1471: romdata_int <= 'h9760;
    1472: romdata_int <= 'h1f4f;
    1473: romdata_int <= 'h6a91;
    1474: romdata_int <= 'hac76;
    1475: romdata_int <= 'h8144;
    1476: romdata_int <= 'he5a; // Line Descriptor
    1477: romdata_int <= 'h9c00;
    1478: romdata_int <= 'h8ef;
    1479: romdata_int <= 'h9b00;
    1480: romdata_int <= 'ha88;
    1481: romdata_int <= 'h3321;
    1482: romdata_int <= 'h855f;
    1483: romdata_int <= 'h8f1c;
    1484: romdata_int <= 'h1355;
    1485: romdata_int <= 'he5a; // Line Descriptor
    1486: romdata_int <= 'h9e00;
    1487: romdata_int <= 'h586b;
    1488: romdata_int <= 'h4915;
    1489: romdata_int <= 'h6f5b;
    1490: romdata_int <= 'h394c;
    1491: romdata_int <= 'h40bd;
    1492: romdata_int <= 'h2511;
    1493: romdata_int <= 'haf61;
    1494: romdata_int <= 'he5a; // Line Descriptor
    1495: romdata_int <= 'ha000;
    1496: romdata_int <= 'h98f2;
    1497: romdata_int <= 'h7334;
    1498: romdata_int <= 'h4f4c;
    1499: romdata_int <= 'h12c;
    1500: romdata_int <= 'h5ea5;
    1501: romdata_int <= 'h8a7e;
    1502: romdata_int <= 'h184f;
    1503: romdata_int <= 'he5a; // Line Descriptor
    1504: romdata_int <= 'ha200;
    1505: romdata_int <= 'h934a;
    1506: romdata_int <= 'h103;
    1507: romdata_int <= 'ha602;
    1508: romdata_int <= 'h2236;
    1509: romdata_int <= 'h53e;
    1510: romdata_int <= 'h32e4;
    1511: romdata_int <= 'h54f5;
    1512: romdata_int <= 'he5a; // Line Descriptor
    1513: romdata_int <= 'ha400;
    1514: romdata_int <= 'h46ad;
    1515: romdata_int <= 'h8e3e;
    1516: romdata_int <= 'ha8f2;
    1517: romdata_int <= 'he2c;
    1518: romdata_int <= 'h26a0;
    1519: romdata_int <= 'h9afc;
    1520: romdata_int <= 'h70b0;
    1521: romdata_int <= 'he5a; // Line Descriptor
    1522: romdata_int <= 'ha600;
    1523: romdata_int <= 'hab4e;
    1524: romdata_int <= 'h6213;
    1525: romdata_int <= 'h7670;
    1526: romdata_int <= 'h7f44;
    1527: romdata_int <= 'h9921;
    1528: romdata_int <= 'h3475;
    1529: romdata_int <= 'h7438;
    1530: romdata_int <= 'he5a; // Line Descriptor
    1531: romdata_int <= 'ha800;
    1532: romdata_int <= 'had1;
    1533: romdata_int <= 'h1eb8;
    1534: romdata_int <= 'h7020;
    1535: romdata_int <= 'h870f;
    1536: romdata_int <= 'h1129;
    1537: romdata_int <= 'h43;
    1538: romdata_int <= 'h6e05;
    1539: romdata_int <= 'he5a; // Line Descriptor
    1540: romdata_int <= 'haa00;
    1541: romdata_int <= 'had50;
    1542: romdata_int <= 'h88f7;
    1543: romdata_int <= 'h2d32;
    1544: romdata_int <= 'h7adf;
    1545: romdata_int <= 'h2925;
    1546: romdata_int <= 'h4a45;
    1547: romdata_int <= 'h5313;
    1548: romdata_int <= 'he5a; // Line Descriptor
    1549: romdata_int <= 'hac00;
    1550: romdata_int <= 'h380a;
    1551: romdata_int <= 'had44;
    1552: romdata_int <= 'hcec;
    1553: romdata_int <= 'h8c89;
    1554: romdata_int <= 'h16aa;
    1555: romdata_int <= 'hb366;
    1556: romdata_int <= 'h88ce;
    1557: romdata_int <= 'he5a; // Line Descriptor
    1558: romdata_int <= 'hae00;
    1559: romdata_int <= 'h80e1;
    1560: romdata_int <= 'haa42;
    1561: romdata_int <= 'h6328;
    1562: romdata_int <= 'h18b5;
    1563: romdata_int <= 'h5c19;
    1564: romdata_int <= 'h824;
    1565: romdata_int <= 'ha6d9;
    1566: romdata_int <= 'he5a; // Line Descriptor
    1567: romdata_int <= 'hb000;
    1568: romdata_int <= 'h3645;
    1569: romdata_int <= 'h7e84;
    1570: romdata_int <= 'ha2fd;
    1571: romdata_int <= 'h90ad;
    1572: romdata_int <= 'hf09;
    1573: romdata_int <= 'ha4a7;
    1574: romdata_int <= 'h86e8;
    1575: romdata_int <= 'he5a; // Line Descriptor
    1576: romdata_int <= 'hb200;
    1577: romdata_int <= 'h4325;
    1578: romdata_int <= 'h7517;
    1579: romdata_int <= 'h60d3;
    1580: romdata_int <= 'h30cc;
    1581: romdata_int <= 'h7c62;
    1582: romdata_int <= 'h3a8d;
    1583: romdata_int <= 'h924e;
    1584: romdata_int <= 'h45a; // Line Descriptor
    1585: romdata_int <= 'h0;
    1586: romdata_int <= 'h9aa1;
    1587: romdata_int <= 'h4715;
    1588: romdata_int <= 'h45a; // Line Descriptor
    1589: romdata_int <= 'h200;
    1590: romdata_int <= 'h4c2b;
    1591: romdata_int <= 'h1401;
    1592: romdata_int <= 'h45a; // Line Descriptor
    1593: romdata_int <= 'h400;
    1594: romdata_int <= 'h2672;
    1595: romdata_int <= 'h7802;
    1596: romdata_int <= 'h45a; // Line Descriptor
    1597: romdata_int <= 'h600;
    1598: romdata_int <= 'h910b;
    1599: romdata_int <= 'h5808;
    1600: romdata_int <= 'h45a; // Line Descriptor
    1601: romdata_int <= 'h800;
    1602: romdata_int <= 'h6a89;
    1603: romdata_int <= 'h422e;
    1604: romdata_int <= 'h45a; // Line Descriptor
    1605: romdata_int <= 'ha00;
    1606: romdata_int <= 'h29a;
    1607: romdata_int <= 'h9cb0;
    1608: romdata_int <= 'h45a; // Line Descriptor
    1609: romdata_int <= 'hc00;
    1610: romdata_int <= 'haeec;
    1611: romdata_int <= 'h700b;
    1612: romdata_int <= 'h45a; // Line Descriptor
    1613: romdata_int <= 'he00;
    1614: romdata_int <= 'h883a;
    1615: romdata_int <= 'hb2a1;
    1616: romdata_int <= 'h45a; // Line Descriptor
    1617: romdata_int <= 'h1000;
    1618: romdata_int <= 'h9d38;
    1619: romdata_int <= 'h7659;
    1620: romdata_int <= 'h45a; // Line Descriptor
    1621: romdata_int <= 'h1200;
    1622: romdata_int <= 'h2eb8;
    1623: romdata_int <= 'h387b;
    1624: romdata_int <= 'h45a; // Line Descriptor
    1625: romdata_int <= 'h1400;
    1626: romdata_int <= 'h3eb9;
    1627: romdata_int <= 'h1b3b;
    1628: romdata_int <= 'h45a; // Line Descriptor
    1629: romdata_int <= 'h1600;
    1630: romdata_int <= 'h3c9b;
    1631: romdata_int <= 'h8312;
    1632: romdata_int <= 'h45a; // Line Descriptor
    1633: romdata_int <= 'h1800;
    1634: romdata_int <= 'h4f65;
    1635: romdata_int <= 'h9ec7;
    1636: romdata_int <= 'h45a; // Line Descriptor
    1637: romdata_int <= 'h1a00;
    1638: romdata_int <= 'h2279;
    1639: romdata_int <= 'h861e;
    1640: romdata_int <= 'h45a; // Line Descriptor
    1641: romdata_int <= 'h1c00;
    1642: romdata_int <= 'h5eef;
    1643: romdata_int <= 'h4c2a;
    1644: romdata_int <= 'h45a; // Line Descriptor
    1645: romdata_int <= 'h1e00;
    1646: romdata_int <= 'h4928;
    1647: romdata_int <= 'h48a;
    1648: romdata_int <= 'h45a; // Line Descriptor
    1649: romdata_int <= 'h2000;
    1650: romdata_int <= 'h3455;
    1651: romdata_int <= 'h3061;
    1652: romdata_int <= 'h45a; // Line Descriptor
    1653: romdata_int <= 'h2200;
    1654: romdata_int <= 'h6ea5;
    1655: romdata_int <= 'h90e0;
    1656: romdata_int <= 'h45a; // Line Descriptor
    1657: romdata_int <= 'h2400;
    1658: romdata_int <= 'h76ae;
    1659: romdata_int <= 'h9911;
    1660: romdata_int <= 'h45a; // Line Descriptor
    1661: romdata_int <= 'h2600;
    1662: romdata_int <= 'ha562;
    1663: romdata_int <= 'h4e5f;
    1664: romdata_int <= 'h45a; // Line Descriptor
    1665: romdata_int <= 'h2800;
    1666: romdata_int <= 'hb0dd;
    1667: romdata_int <= 'h232e;
    1668: romdata_int <= 'h45a; // Line Descriptor
    1669: romdata_int <= 'h2a00;
    1670: romdata_int <= 'h792c;
    1671: romdata_int <= 'h52a7;
    1672: romdata_int <= 'h45a; // Line Descriptor
    1673: romdata_int <= 'h2c00;
    1674: romdata_int <= 'h5243;
    1675: romdata_int <= 'h1328;
    1676: romdata_int <= 'h45a; // Line Descriptor
    1677: romdata_int <= 'h2e00;
    1678: romdata_int <= 'h5673;
    1679: romdata_int <= 'h207c;
    1680: romdata_int <= 'h45a; // Line Descriptor
    1681: romdata_int <= 'h3000;
    1682: romdata_int <= 'h726a;
    1683: romdata_int <= 'h6494;
    1684: romdata_int <= 'h45a; // Line Descriptor
    1685: romdata_int <= 'h3200;
    1686: romdata_int <= 'h7a4e;
    1687: romdata_int <= 'h4ac4;
    1688: romdata_int <= 'h45a; // Line Descriptor
    1689: romdata_int <= 'h3400;
    1690: romdata_int <= 'ha60f;
    1691: romdata_int <= 'h92d8;
    1692: romdata_int <= 'h45a; // Line Descriptor
    1693: romdata_int <= 'h3600;
    1694: romdata_int <= 'h1f2b;
    1695: romdata_int <= 'h1c64;
    1696: romdata_int <= 'h45a; // Line Descriptor
    1697: romdata_int <= 'h3800;
    1698: romdata_int <= 'h40d5;
    1699: romdata_int <= 'ha062;
    1700: romdata_int <= 'h45a; // Line Descriptor
    1701: romdata_int <= 'h3a00;
    1702: romdata_int <= 'h7cc9;
    1703: romdata_int <= 'h5f54;
    1704: romdata_int <= 'h45a; // Line Descriptor
    1705: romdata_int <= 'h3c00;
    1706: romdata_int <= 'h1ae7;
    1707: romdata_int <= 'h3613;
    1708: romdata_int <= 'h45a; // Line Descriptor
    1709: romdata_int <= 'h3e00;
    1710: romdata_int <= 'h1c83;
    1711: romdata_int <= 'h2b18;
    1712: romdata_int <= 'h45a; // Line Descriptor
    1713: romdata_int <= 'h4000;
    1714: romdata_int <= 'h760;
    1715: romdata_int <= 'h6ac5;
    1716: romdata_int <= 'h45a; // Line Descriptor
    1717: romdata_int <= 'h4200;
    1718: romdata_int <= 'ha949;
    1719: romdata_int <= 'h9667;
    1720: romdata_int <= 'h45a; // Line Descriptor
    1721: romdata_int <= 'h4400;
    1722: romdata_int <= 'h5088;
    1723: romdata_int <= 'h7b27;
    1724: romdata_int <= 'h45a; // Line Descriptor
    1725: romdata_int <= 'h4600;
    1726: romdata_int <= 'h5c48;
    1727: romdata_int <= 'h2d22;
    1728: romdata_int <= 'h45a; // Line Descriptor
    1729: romdata_int <= 'h4800;
    1730: romdata_int <= 'h8322;
    1731: romdata_int <= 'ha27c;
    1732: romdata_int <= 'h45a; // Line Descriptor
    1733: romdata_int <= 'h4a00;
    1734: romdata_int <= 'h2055;
    1735: romdata_int <= 'h692b;
    1736: romdata_int <= 'h45a; // Line Descriptor
    1737: romdata_int <= 'h4c00;
    1738: romdata_int <= 'hb5;
    1739: romdata_int <= 'h285e;
    1740: romdata_int <= 'h45a; // Line Descriptor
    1741: romdata_int <= 'h4e00;
    1742: romdata_int <= 'h9482;
    1743: romdata_int <= 'h5070;
    1744: romdata_int <= 'h45a; // Line Descriptor
    1745: romdata_int <= 'h5000;
    1746: romdata_int <= 'ha34d;
    1747: romdata_int <= 'hd52;
    1748: romdata_int <= 'h45a; // Line Descriptor
    1749: romdata_int <= 'h5200;
    1750: romdata_int <= 'h960e;
    1751: romdata_int <= 'h44ab;
    1752: romdata_int <= 'h45a; // Line Descriptor
    1753: romdata_int <= 'h5400;
    1754: romdata_int <= 'h324c;
    1755: romdata_int <= 'h18c5;
    1756: romdata_int <= 'h45a; // Line Descriptor
    1757: romdata_int <= 'h5600;
    1758: romdata_int <= 'h1361;
    1759: romdata_int <= 'h8a8a;
    1760: romdata_int <= 'h45a; // Line Descriptor
    1761: romdata_int <= 'h5800;
    1762: romdata_int <= 'ha164;
    1763: romdata_int <= 'h3ee9;
    1764: romdata_int <= 'h45a; // Line Descriptor
    1765: romdata_int <= 'h5a00;
    1766: romdata_int <= 'h24a1;
    1767: romdata_int <= 'h844d;
    1768: romdata_int <= 'h45a; // Line Descriptor
    1769: romdata_int <= 'h5c00;
    1770: romdata_int <= 'h9e0a;
    1771: romdata_int <= 'h916;
    1772: romdata_int <= 'h45a; // Line Descriptor
    1773: romdata_int <= 'h5e00;
    1774: romdata_int <= 'h6c32;
    1775: romdata_int <= 'h34f3;
    1776: romdata_int <= 'h45a; // Line Descriptor
    1777: romdata_int <= 'h6000;
    1778: romdata_int <= 'h8a58;
    1779: romdata_int <= 'haef1;
    1780: romdata_int <= 'h45a; // Line Descriptor
    1781: romdata_int <= 'h6200;
    1782: romdata_int <= 'h2c37;
    1783: romdata_int <= 'h66e5;
    1784: romdata_int <= 'h45a; // Line Descriptor
    1785: romdata_int <= 'h6400;
    1786: romdata_int <= 'h5449;
    1787: romdata_int <= 'h3c1e;
    1788: romdata_int <= 'h45a; // Line Descriptor
    1789: romdata_int <= 'h6600;
    1790: romdata_int <= 'h688d;
    1791: romdata_int <= 'h1031;
    1792: romdata_int <= 'h45a; // Line Descriptor
    1793: romdata_int <= 'h6800;
    1794: romdata_int <= 'h4544;
    1795: romdata_int <= 'h6e06;
    1796: romdata_int <= 'h55a; // Line Descriptor
    1797: romdata_int <= 'h6a00;
    1798: romdata_int <= 'hed6;
    1799: romdata_int <= 'h56df;
    1800: romdata_int <= 'h1648; // Line Descriptor
    1801: romdata_int <= 'h3d37;
    1802: romdata_int <= 'h748e;
    1803: romdata_int <= 'h44a1;
    1804: romdata_int <= 'h6b15;
    1805: romdata_int <= 'h29b;
    1806: romdata_int <= 'h5428;
    1807: romdata_int <= 'h342b;
    1808: romdata_int <= 'h3601;
    1809: romdata_int <= 'h124e;
    1810: romdata_int <= 'hed;
    1811: romdata_int <= 'h7c72;
    1812: romdata_int <= 'h4602;
    1813: romdata_int <= 'h1648; // Line Descriptor
    1814: romdata_int <= 'h3f5c;
    1815: romdata_int <= 'h24e1;
    1816: romdata_int <= 'h2eec;
    1817: romdata_int <= 'h480b;
    1818: romdata_int <= 'h3316;
    1819: romdata_int <= 'h3164;
    1820: romdata_int <= 'h143a;
    1821: romdata_int <= 'h4aa1;
    1822: romdata_int <= 'h7f39;
    1823: romdata_int <= 'h32f0;
    1824: romdata_int <= 'h6738;
    1825: romdata_int <= 'h6e59;
    1826: romdata_int <= 'h1648; // Line Descriptor
    1827: romdata_int <= 'h4299;
    1828: romdata_int <= 'h3b3d;
    1829: romdata_int <= 'h565;
    1830: romdata_int <= 'h78c7;
    1831: romdata_int <= 'h384c;
    1832: romdata_int <= 'h2b0b;
    1833: romdata_int <= 'h2879;
    1834: romdata_int <= 'h221e;
    1835: romdata_int <= 'h26bc;
    1836: romdata_int <= 'h549d;
    1837: romdata_int <= 'h72ef;
    1838: romdata_int <= 'h5a2a;
    1839: romdata_int <= 'h1648; // Line Descriptor
    1840: romdata_int <= 'h2ae6;
    1841: romdata_int <= 'h6334;
    1842: romdata_int <= 'h46ae;
    1843: romdata_int <= 'h7b11;
    1844: romdata_int <= 'h4347;
    1845: romdata_int <= 'h46a0;
    1846: romdata_int <= 'h1162;
    1847: romdata_int <= 'h1a5f;
    1848: romdata_int <= 'h7760;
    1849: romdata_int <= 'h4448;
    1850: romdata_int <= 'h1add;
    1851: romdata_int <= 'h2d2e;
    1852: romdata_int <= 'h1648; // Line Descriptor
    1853: romdata_int <= 'h52e5;
    1854: romdata_int <= 'h1ec9;
    1855: romdata_int <= 'h166a;
    1856: romdata_int <= 'h7694;
    1857: romdata_int <= 'h24f2;
    1858: romdata_int <= 'h3e9a;
    1859: romdata_int <= 'h7e4e;
    1860: romdata_int <= 'h56c4;
    1861: romdata_int <= 'h2b50;
    1862: romdata_int <= 'h6123;
    1863: romdata_int <= 'h480f;
    1864: romdata_int <= 'h88d8;
    1865: romdata_int <= 'h1648; // Line Descriptor
    1866: romdata_int <= 'h184a;
    1867: romdata_int <= 'h8877;
    1868: romdata_int <= 'h7ae7;
    1869: romdata_int <= 'h8413;
    1870: romdata_int <= 'h264e;
    1871: romdata_int <= 'h485a;
    1872: romdata_int <= 'h6483;
    1873: romdata_int <= 'h3b18;
    1874: romdata_int <= 'h740e;
    1875: romdata_int <= 'h4ad0;
    1876: romdata_int <= 'h2360;
    1877: romdata_int <= 'h76c5;
    1878: romdata_int <= 'h1648; // Line Descriptor
    1879: romdata_int <= 'h501;
    1880: romdata_int <= 'h7934;
    1881: romdata_int <= 'h4122;
    1882: romdata_int <= 'h307c;
    1883: romdata_int <= 'h2a4b;
    1884: romdata_int <= 'h86d9;
    1885: romdata_int <= 'hc55;
    1886: romdata_int <= 'h872b;
    1887: romdata_int <= 'h8806;
    1888: romdata_int <= 'h805f;
    1889: romdata_int <= 'h36b5;
    1890: romdata_int <= 'h445e;
    1891: romdata_int <= 'h1648; // Line Descriptor
    1892: romdata_int <= 'h1275;
    1893: romdata_int <= 'h1c41;
    1894: romdata_int <= 'h684c;
    1895: romdata_int <= 'h40c5;
    1896: romdata_int <= 'h1a33;
    1897: romdata_int <= 'h8311;
    1898: romdata_int <= 'h961;
    1899: romdata_int <= 'h28a;
    1900: romdata_int <= 'h6b4a;
    1901: romdata_int <= 'h5e7d;
    1902: romdata_int <= 'h2764;
    1903: romdata_int <= 'h64e9;
    1904: romdata_int <= 'h1648; // Line Descriptor
    1905: romdata_int <= 'h592a;
    1906: romdata_int <= 'h5d58;
    1907: romdata_int <= 'h1058;
    1908: romdata_int <= 'h3cf1;
    1909: romdata_int <= 'h1062;
    1910: romdata_int <= 'h42c1;
    1911: romdata_int <= 'h5837;
    1912: romdata_int <= 'h80e5;
    1913: romdata_int <= 'h4b2;
    1914: romdata_int <= 'h1079;
    1915: romdata_int <= 'h3c49;
    1916: romdata_int <= 'h5c1e;
    1917: romdata_int <= 'h1648; // Line Descriptor
    1918: romdata_int <= 'h6b38;
    1919: romdata_int <= 'h6a21;
    1920: romdata_int <= 'h7308;
    1921: romdata_int <= 'h5228;
    1922: romdata_int <= 'h172c;
    1923: romdata_int <= 'h21a;
    1924: romdata_int <= 'h2668;
    1925: romdata_int <= 'h5a4e;
    1926: romdata_int <= 'h4d3f;
    1927: romdata_int <= 'h2141;
    1928: romdata_int <= 'h2f1d;
    1929: romdata_int <= 'h6312;
    1930: romdata_int <= 'h1648; // Line Descriptor
    1931: romdata_int <= 'h5418;
    1932: romdata_int <= 'h3840;
    1933: romdata_int <= 'h2922;
    1934: romdata_int <= 'h36cf;
    1935: romdata_int <= 'h3e80;
    1936: romdata_int <= 'h38ab;
    1937: romdata_int <= 'h8098;
    1938: romdata_int <= 'hcb4;
    1939: romdata_int <= 'he3e;
    1940: romdata_int <= 'h8625;
    1941: romdata_int <= 'h3ae4;
    1942: romdata_int <= 'h8e0a;
    1943: romdata_int <= 'h1648; // Line Descriptor
    1944: romdata_int <= 'h165c;
    1945: romdata_int <= 'h18ca;
    1946: romdata_int <= 'h306;
    1947: romdata_int <= 'h3b37;
    1948: romdata_int <= 'h2933;
    1949: romdata_int <= 'h32b0;
    1950: romdata_int <= 'h1688;
    1951: romdata_int <= 'h8b61;
    1952: romdata_int <= 'h506b;
    1953: romdata_int <= 'h4cfd;
    1954: romdata_int <= 'h129d;
    1955: romdata_int <= 'h87d;
    1956: romdata_int <= 'h1648; // Line Descriptor
    1957: romdata_int <= 'h4d15;
    1958: romdata_int <= 'h774c;
    1959: romdata_int <= 'h6106;
    1960: romdata_int <= 'hc64;
    1961: romdata_int <= 'h58ad;
    1962: romdata_int <= 'h7c3c;
    1963: romdata_int <= 'h6716;
    1964: romdata_int <= 'h7255;
    1965: romdata_int <= 'h6f23;
    1966: romdata_int <= 'h5610;
    1967: romdata_int <= 'h747;
    1968: romdata_int <= 'h8b58;
    1969: romdata_int <= 'h1648; // Line Descriptor
    1970: romdata_int <= 'h480a;
    1971: romdata_int <= 'h8c9a;
    1972: romdata_int <= 'h3ccb;
    1973: romdata_int <= 'h1d1d;
    1974: romdata_int <= 'h5e32;
    1975: romdata_int <= 'h20f6;
    1976: romdata_int <= 'h18a2;
    1977: romdata_int <= 'h46a4;
    1978: romdata_int <= 'h62b3;
    1979: romdata_int <= 'h143d;
    1980: romdata_int <= 'h6a72;
    1981: romdata_int <= 'h613e;
    1982: romdata_int <= 'h1648; // Line Descriptor
    1983: romdata_int <= 'h2481;
    1984: romdata_int <= 'h434d;
    1985: romdata_int <= 'h88b;
    1986: romdata_int <= 'h8299;
    1987: romdata_int <= 'h434;
    1988: romdata_int <= 'h7b51;
    1989: romdata_int <= 'h886f;
    1990: romdata_int <= 'h3513;
    1991: romdata_int <= 'h640b;
    1992: romdata_int <= 'h687a;
    1993: romdata_int <= 'h2428;
    1994: romdata_int <= 'h6645;
    1995: romdata_int <= 'h1648; // Line Descriptor
    1996: romdata_int <= 'h1e69;
    1997: romdata_int <= 'h4e67;
    1998: romdata_int <= 'h595e;
    1999: romdata_int <= 'h7041;
    2000: romdata_int <= 'hc8;
    2001: romdata_int <= 'h1b3f;
    2002: romdata_int <= 'h8e4c;
    2003: romdata_int <= 'h1c6f;
    2004: romdata_int <= 'h1750;
    2005: romdata_int <= 'h2ab5;
    2006: romdata_int <= 'h500f;
    2007: romdata_int <= 'h2047;
    2008: romdata_int <= 'h1648; // Line Descriptor
    2009: romdata_int <= 'h3430;
    2010: romdata_int <= 'h6c80;
    2011: romdata_int <= 'h36b5;
    2012: romdata_int <= 'h72db;
    2013: romdata_int <= 'h4a67;
    2014: romdata_int <= 'h7749;
    2015: romdata_int <= 'h7032;
    2016: romdata_int <= 'h4355;
    2017: romdata_int <= 'h6ce5;
    2018: romdata_int <= 'h16f3;
    2019: romdata_int <= 'h8d37;
    2020: romdata_int <= 'h6ccb;
    2021: romdata_int <= 'h1648; // Line Descriptor
    2022: romdata_int <= 'h6d9;
    2023: romdata_int <= 'h34d4;
    2024: romdata_int <= 'h2c3a;
    2025: romdata_int <= 'h893b;
    2026: romdata_int <= 'h1451;
    2027: romdata_int <= 'h6ba;
    2028: romdata_int <= 'h1d4c;
    2029: romdata_int <= 'h82eb;
    2030: romdata_int <= 'h32cf;
    2031: romdata_int <= 'h6c33;
    2032: romdata_int <= 'hd60;
    2033: romdata_int <= 'h4b4f;
    2034: romdata_int <= 'h1648; // Line Descriptor
    2035: romdata_int <= 'h7159;
    2036: romdata_int <= 'h2ae3;
    2037: romdata_int <= 'hee4;
    2038: romdata_int <= 'h8aba;
    2039: romdata_int <= 'h6ee6;
    2040: romdata_int <= 'h5670;
    2041: romdata_int <= 'h5b57;
    2042: romdata_int <= 'h832;
    2043: romdata_int <= 'h7167;
    2044: romdata_int <= 'h879;
    2045: romdata_int <= 'h3885;
    2046: romdata_int <= 'h7b1a;
    2047: romdata_int <= 'h1648; // Line Descriptor
    2048: romdata_int <= 'h7233;
    2049: romdata_int <= 'h4aef;
    2050: romdata_int <= 'h2100;
    2051: romdata_int <= 'h8c88;
    2052: romdata_int <= 'h2f21;
    2053: romdata_int <= 'h6d5f;
    2054: romdata_int <= 'h8b1c;
    2055: romdata_int <= 'h8555;
    2056: romdata_int <= 'h44b8;
    2057: romdata_int <= 'h7646;
    2058: romdata_int <= 'h8ec4;
    2059: romdata_int <= 'h287a;
    2060: romdata_int <= 'h1648; // Line Descriptor
    2061: romdata_int <= 'h4ee4;
    2062: romdata_int <= 'hcf5;
    2063: romdata_int <= 'h50d5;
    2064: romdata_int <= 'h64fc;
    2065: romdata_int <= 'h5162;
    2066: romdata_int <= 'h6218;
    2067: romdata_int <= 'h2454;
    2068: romdata_int <= 'h4f2f;
    2069: romdata_int <= 'h58c7;
    2070: romdata_int <= 'h7aad;
    2071: romdata_int <= 'h303e;
    2072: romdata_int <= 'h84f2;
    2073: romdata_int <= 'h1648; // Line Descriptor
    2074: romdata_int <= 'h4013;
    2075: romdata_int <= 'h8e70;
    2076: romdata_int <= 'h5f44;
    2077: romdata_int <= 'h8f21;
    2078: romdata_int <= 'h6875;
    2079: romdata_int <= 'h6838;
    2080: romdata_int <= 'h60b3;
    2081: romdata_int <= 'h6162;
    2082: romdata_int <= 'h7b35;
    2083: romdata_int <= 'h2ce6;
    2084: romdata_int <= 'h8458;
    2085: romdata_int <= 'h3152;
    2086: romdata_int <= 'h1648; // Line Descriptor
    2087: romdata_int <= 'h7f5c;
    2088: romdata_int <= 'h5547;
    2089: romdata_int <= 'h7001;
    2090: romdata_int <= 'h1242;
    2091: romdata_int <= 'h691;
    2092: romdata_int <= 'h139;
    2093: romdata_int <= 'h4e77;
    2094: romdata_int <= 'h4087;
    2095: romdata_int <= 'h3d61;
    2096: romdata_int <= 'had1;
    2097: romdata_int <= 'h7019;
    2098: romdata_int <= 'h1038;
    2099: romdata_int <= 'h1648; // Line Descriptor
    2100: romdata_int <= 'h2205;
    2101: romdata_int <= 'h8125;
    2102: romdata_int <= 'h14bb;
    2103: romdata_int <= 'h664b;
    2104: romdata_int <= 'h44ee;
    2105: romdata_int <= 'h4452;
    2106: romdata_int <= 'h408e;
    2107: romdata_int <= 'h28a6;
    2108: romdata_int <= 'h2550;
    2109: romdata_int <= 'h62f7;
    2110: romdata_int <= 'h1f32;
    2111: romdata_int <= 'h68df;
    2112: romdata_int <= 'h1648; // Line Descriptor
    2113: romdata_int <= 'h56b5;
    2114: romdata_int <= 'h86;
    2115: romdata_int <= 'h8554;
    2116: romdata_int <= 'h5cb6;
    2117: romdata_int <= 'h474b;
    2118: romdata_int <= 'h4a65;
    2119: romdata_int <= 'h8d12;
    2120: romdata_int <= 'h4829;
    2121: romdata_int <= 'h14ea;
    2122: romdata_int <= 'h243;
    2123: romdata_int <= 'h5d4c;
    2124: romdata_int <= 'had2;
    2125: romdata_int <= 'h1648; // Line Descriptor
    2126: romdata_int <= 'hd1d;
    2127: romdata_int <= 'h3231;
    2128: romdata_int <= 'haa0;
    2129: romdata_int <= 'h4d44;
    2130: romdata_int <= 'h822;
    2131: romdata_int <= 'h74f4;
    2132: romdata_int <= 'h530b;
    2133: romdata_int <= 'h1918;
    2134: romdata_int <= 'h78fa;
    2135: romdata_int <= 'h5355;
    2136: romdata_int <= 'heb8;
    2137: romdata_int <= 'h5015;
    2138: romdata_int <= 'h1648; // Line Descriptor
    2139: romdata_int <= 'h5f05;
    2140: romdata_int <= 'h4925;
    2141: romdata_int <= 'h3f17;
    2142: romdata_int <= 'h2cd3;
    2143: romdata_int <= 'h22cc;
    2144: romdata_int <= 'h5062;
    2145: romdata_int <= 'h2c8d;
    2146: romdata_int <= 'h5e4e;
    2147: romdata_int <= 'h703;
    2148: romdata_int <= 'h5911;
    2149: romdata_int <= 'h88ad;
    2150: romdata_int <= 'h82c2;
    2151: romdata_int <= 'h1648; // Line Descriptor
    2152: romdata_int <= 'h2e39;
    2153: romdata_int <= 'h2629;
    2154: romdata_int <= 'h6f3;
    2155: romdata_int <= 'h1ee2;
    2156: romdata_int <= 'h6136;
    2157: romdata_int <= 'hf2a;
    2158: romdata_int <= 'h2e6e;
    2159: romdata_int <= 'h2106;
    2160: romdata_int <= 'h2e4d;
    2161: romdata_int <= 'h6e6f;
    2162: romdata_int <= 'h4744;
    2163: romdata_int <= 'h3a5e;
    2164: romdata_int <= 'h1648; // Line Descriptor
    2165: romdata_int <= 'h8693;
    2166: romdata_int <= 'h7f53;
    2167: romdata_int <= 'h8ac6;
    2168: romdata_int <= 'h6238;
    2169: romdata_int <= 'h7464;
    2170: romdata_int <= 'h6a44;
    2171: romdata_int <= 'h7861;
    2172: romdata_int <= 'h8c0e;
    2173: romdata_int <= 'ha0b;
    2174: romdata_int <= 'h1d3e;
    2175: romdata_int <= 'h351c;
    2176: romdata_int <= 'h8c3b;
    2177: romdata_int <= 'h1648; // Line Descriptor
    2178: romdata_int <= 'h7d28;
    2179: romdata_int <= 'h6eb7;
    2180: romdata_int <= 'h233f;
    2181: romdata_int <= 'h2046;
    2182: romdata_int <= 'ha35;
    2183: romdata_int <= 'h3d49;
    2184: romdata_int <= 'h84c4;
    2185: romdata_int <= 'h548a;
    2186: romdata_int <= 'h2d08;
    2187: romdata_int <= 'h6547;
    2188: romdata_int <= 'h4e7b;
    2189: romdata_int <= 'h1d60;
    2190: romdata_int <= 'h1648; // Line Descriptor
    2191: romdata_int <= 'he56;
    2192: romdata_int <= 'h3132;
    2193: romdata_int <= 'h5a6b;
    2194: romdata_int <= 'h7cb8;
    2195: romdata_int <= 'h4e37;
    2196: romdata_int <= 'h1349;
    2197: romdata_int <= 'h3ae4;
    2198: romdata_int <= 'h393a;
    2199: romdata_int <= 'h5248;
    2200: romdata_int <= 'h5b37;
    2201: romdata_int <= 'h434f;
    2202: romdata_int <= 'h1483;
    2203: romdata_int <= 'h1648; // Line Descriptor
    2204: romdata_int <= 'h746e;
    2205: romdata_int <= 'h12a9;
    2206: romdata_int <= 'h1a28;
    2207: romdata_int <= 'h5520;
    2208: romdata_int <= 'he2c;
    2209: romdata_int <= 'ha78;
    2210: romdata_int <= 'h6ea4;
    2211: romdata_int <= 'h8f55;
    2212: romdata_int <= 'h1e8f;
    2213: romdata_int <= 'h7f65;
    2214: romdata_int <= 'h82ec;
    2215: romdata_int <= 'h2633;
    2216: romdata_int <= 'h1648; // Line Descriptor
    2217: romdata_int <= 'h331c;
    2218: romdata_int <= 'h7c9c;
    2219: romdata_int <= 'h6489;
    2220: romdata_int <= 'h7f3c;
    2221: romdata_int <= 'h6c23;
    2222: romdata_int <= 'h1e75;
    2223: romdata_int <= 'h3633;
    2224: romdata_int <= 'h3e4b;
    2225: romdata_int <= 'h159;
    2226: romdata_int <= 'h2930;
    2227: romdata_int <= 'h40df;
    2228: romdata_int <= 'h38fd;
    2229: romdata_int <= 'h1648; // Line Descriptor
    2230: romdata_int <= 'h72;
    2231: romdata_int <= 'h864f;
    2232: romdata_int <= 'h6708;
    2233: romdata_int <= 'h5a76;
    2234: romdata_int <= 'h195a;
    2235: romdata_int <= 'h5c59;
    2236: romdata_int <= 'h49c;
    2237: romdata_int <= 'h6891;
    2238: romdata_int <= 'h7ce3;
    2239: romdata_int <= 'h3e96;
    2240: romdata_int <= 'h789e;
    2241: romdata_int <= 'h286;
    2242: romdata_int <= 'h1648; // Line Descriptor
    2243: romdata_int <= 'h80e1;
    2244: romdata_int <= 'h569c;
    2245: romdata_int <= 'h535a;
    2246: romdata_int <= 'h5620;
    2247: romdata_int <= 'h86af;
    2248: romdata_int <= 'h4d0a;
    2249: romdata_int <= 'h7264;
    2250: romdata_int <= 'h5c63;
    2251: romdata_int <= 'h6758;
    2252: romdata_int <= 'h7428;
    2253: romdata_int <= 'h423;
    2254: romdata_int <= 'h1aa3;
    2255: romdata_int <= 'h1648; // Line Descriptor
    2256: romdata_int <= 'h3632;
    2257: romdata_int <= 'h8252;
    2258: romdata_int <= 'h4cc0;
    2259: romdata_int <= 'h3415;
    2260: romdata_int <= 'h8141;
    2261: romdata_int <= 'h2258;
    2262: romdata_int <= 'h5e27;
    2263: romdata_int <= 'h10f6;
    2264: romdata_int <= 'h3022;
    2265: romdata_int <= 'h1867;
    2266: romdata_int <= 'h8a07;
    2267: romdata_int <= 'h78d0;
    2268: romdata_int <= 'h448; // Line Descriptor
    2269: romdata_int <= 'h0;
    2270: romdata_int <= 'h4701;
    2271: romdata_int <= 'h1b03;
    2272: romdata_int <= 'h448; // Line Descriptor
    2273: romdata_int <= 'h200;
    2274: romdata_int <= 'h7c91;
    2275: romdata_int <= 'h6429;
    2276: romdata_int <= 'h448; // Line Descriptor
    2277: romdata_int <= 'h400;
    2278: romdata_int <= 'h1082;
    2279: romdata_int <= 'h4295;
    2280: romdata_int <= 'h448; // Line Descriptor
    2281: romdata_int <= 'h600;
    2282: romdata_int <= 'h76aa;
    2283: romdata_int <= 'h686c;
    2284: romdata_int <= 'h448; // Line Descriptor
    2285: romdata_int <= 'h800;
    2286: romdata_int <= 'hd1;
    2287: romdata_int <= 'h54b9;
    2288: romdata_int <= 'h448; // Line Descriptor
    2289: romdata_int <= 'ha00;
    2290: romdata_int <= 'h1900;
    2291: romdata_int <= 'h2156;
    2292: romdata_int <= 'h448; // Line Descriptor
    2293: romdata_int <= 'hc00;
    2294: romdata_int <= 'h4f20;
    2295: romdata_int <= 'h2f0a;
    2296: romdata_int <= 'h448; // Line Descriptor
    2297: romdata_int <= 'he00;
    2298: romdata_int <= 'h4507;
    2299: romdata_int <= 'h3698;
    2300: romdata_int <= 'h448; // Line Descriptor
    2301: romdata_int <= 'h1000;
    2302: romdata_int <= 'h24a;
    2303: romdata_int <= 'h4d15;
    2304: romdata_int <= 'h448; // Line Descriptor
    2305: romdata_int <= 'h1200;
    2306: romdata_int <= 'h809c;
    2307: romdata_int <= 'hf03;
    2308: romdata_int <= 'h448; // Line Descriptor
    2309: romdata_int <= 'h1400;
    2310: romdata_int <= 'h8cd0;
    2311: romdata_int <= 'h871e;
    2312: romdata_int <= 'h448; // Line Descriptor
    2313: romdata_int <= 'h1600;
    2314: romdata_int <= 'h3865;
    2315: romdata_int <= 'h4933;
    2316: romdata_int <= 'h448; // Line Descriptor
    2317: romdata_int <= 'h1800;
    2318: romdata_int <= 'h8b31;
    2319: romdata_int <= 'hac9;
    2320: romdata_int <= 'h448; // Line Descriptor
    2321: romdata_int <= 'h1a00;
    2322: romdata_int <= 'h529a;
    2323: romdata_int <= 'h2c0a;
    2324: romdata_int <= 'h448; // Line Descriptor
    2325: romdata_int <= 'h1c00;
    2326: romdata_int <= 'hcb8;
    2327: romdata_int <= 'h7abf;
    2328: romdata_int <= 'h448; // Line Descriptor
    2329: romdata_int <= 'h1e00;
    2330: romdata_int <= 'h150b;
    2331: romdata_int <= 'h32b8;
    2332: romdata_int <= 'h448; // Line Descriptor
    2333: romdata_int <= 'h2000;
    2334: romdata_int <= 'h3e54;
    2335: romdata_int <= 'h3525;
    2336: romdata_int <= 'h448; // Line Descriptor
    2337: romdata_int <= 'h2200;
    2338: romdata_int <= 'h3d3c;
    2339: romdata_int <= 'h8850;
    2340: romdata_int <= 'h448; // Line Descriptor
    2341: romdata_int <= 'h2400;
    2342: romdata_int <= 'h5f12;
    2343: romdata_int <= 'h8e3a;
    2344: romdata_int <= 'h448; // Line Descriptor
    2345: romdata_int <= 'h2600;
    2346: romdata_int <= 'h817;
    2347: romdata_int <= 'h5b0d;
    2348: romdata_int <= 'h448; // Line Descriptor
    2349: romdata_int <= 'h2800;
    2350: romdata_int <= 'h163d;
    2351: romdata_int <= 'h6232;
    2352: romdata_int <= 'h448; // Line Descriptor
    2353: romdata_int <= 'h2a00;
    2354: romdata_int <= 'h66b9;
    2355: romdata_int <= 'h767;
    2356: romdata_int <= 'h448; // Line Descriptor
    2357: romdata_int <= 'h2c00;
    2358: romdata_int <= 'h253c;
    2359: romdata_int <= 'h512e;
    2360: romdata_int <= 'h448; // Line Descriptor
    2361: romdata_int <= 'h2e00;
    2362: romdata_int <= 'h3a95;
    2363: romdata_int <= 'h26c4;
    2364: romdata_int <= 'h448; // Line Descriptor
    2365: romdata_int <= 'h3000;
    2366: romdata_int <= 'h1edf;
    2367: romdata_int <= 'h232c;
    2368: romdata_int <= 'h448; // Line Descriptor
    2369: romdata_int <= 'h3200;
    2370: romdata_int <= 'h7258;
    2371: romdata_int <= 'h6a33;
    2372: romdata_int <= 'h448; // Line Descriptor
    2373: romdata_int <= 'h3400;
    2374: romdata_int <= 'h2a08;
    2375: romdata_int <= 'h3115;
    2376: romdata_int <= 'h448; // Line Descriptor
    2377: romdata_int <= 'h3600;
    2378: romdata_int <= 'h6e4f;
    2379: romdata_int <= 'h2870;
    2380: romdata_int <= 'h448; // Line Descriptor
    2381: romdata_int <= 'h3800;
    2382: romdata_int <= 'h45e;
    2383: romdata_int <= 'h5884;
    2384: romdata_int <= 'h448; // Line Descriptor
    2385: romdata_int <= 'h3a00;
    2386: romdata_int <= 'h4a3b;
    2387: romdata_int <= 'h5cf3;
    2388: romdata_int <= 'h448; // Line Descriptor
    2389: romdata_int <= 'h3c00;
    2390: romdata_int <= 'h40bc;
    2391: romdata_int <= 'h7f39;
    2392: romdata_int <= 'h448; // Line Descriptor
    2393: romdata_int <= 'h3e00;
    2394: romdata_int <= 'h7418;
    2395: romdata_int <= 'h1240;
    2396: romdata_int <= 'h448; // Line Descriptor
    2397: romdata_int <= 'h4000;
    2398: romdata_int <= 'h6d42;
    2399: romdata_int <= 'h70a1;
    2400: romdata_int <= 'h448; // Line Descriptor
    2401: romdata_int <= 'h4200;
    2402: romdata_int <= 'h5710;
    2403: romdata_int <= 'h1c1c;
    2404: romdata_int <= 'h448; // Line Descriptor
    2405: romdata_int <= 'h4400;
    2406: romdata_int <= 'h82bc;
    2407: romdata_int <= 'h84ba;
    2408: romdata_int <= 'h448; // Line Descriptor
    2409: romdata_int <= 'h4600;
    2410: romdata_int <= 'h78be;
    2411: romdata_int <= 'h60f0;
    2412: romdata_int <= 'h448; // Line Descriptor
    2413: romdata_int <= 'h4800;
    2414: romdata_int <= 'h395b;
    2415: romdata_int <= 'h60c1;
    2416: romdata_int <= 'h448; // Line Descriptor
    2417: romdata_int <= 'h4a00;
    2418: romdata_int <= 'h6338;
    2419: romdata_int <= 'h7e5c;
    2420: romdata_int <= 'h448; // Line Descriptor
    2421: romdata_int <= 'h4c00;
    2422: romdata_int <= 'h4c44;
    2423: romdata_int <= 'h76ae;
    2424: romdata_int <= 'h448; // Line Descriptor
    2425: romdata_int <= 'h4e00;
    2426: romdata_int <= 'h3b26;
    2427: romdata_int <= 'h2a47;
    2428: romdata_int <= 'h448; // Line Descriptor
    2429: romdata_int <= 'h5000;
    2430: romdata_int <= 'h333b;
    2431: romdata_int <= 'h3460;
    2432: romdata_int <= 'h448; // Line Descriptor
    2433: romdata_int <= 'h5200;
    2434: romdata_int <= 'h5c68;
    2435: romdata_int <= 'h1356;
    2436: romdata_int <= 'h448; // Line Descriptor
    2437: romdata_int <= 'h5400;
    2438: romdata_int <= 'h8152;
    2439: romdata_int <= 'h6ab1;
    2440: romdata_int <= 'h448; // Line Descriptor
    2441: romdata_int <= 'h5600;
    2442: romdata_int <= 'h2f30;
    2443: romdata_int <= 'h1165;
    2444: romdata_int <= 'h448; // Line Descriptor
    2445: romdata_int <= 'h5800;
    2446: romdata_int <= 'h1ea7;
    2447: romdata_int <= 'h780f;
    2448: romdata_int <= 'h448; // Line Descriptor
    2449: romdata_int <= 'h5a00;
    2450: romdata_int <= 'h5551;
    2451: romdata_int <= 'h1a0e;
    2452: romdata_int <= 'h448; // Line Descriptor
    2453: romdata_int <= 'h5c00;
    2454: romdata_int <= 'h58c2;
    2455: romdata_int <= 'h1720;
    2456: romdata_int <= 'h448; // Line Descriptor
    2457: romdata_int <= 'h5e00;
    2458: romdata_int <= 'h429c;
    2459: romdata_int <= 'h36d3;
    2460: romdata_int <= 'h448; // Line Descriptor
    2461: romdata_int <= 'h6000;
    2462: romdata_int <= 'h7c40;
    2463: romdata_int <= 'h66d7;
    2464: romdata_int <= 'h448; // Line Descriptor
    2465: romdata_int <= 'h6200;
    2466: romdata_int <= 'h7282;
    2467: romdata_int <= 'h3ec7;
    2468: romdata_int <= 'h448; // Line Descriptor
    2469: romdata_int <= 'h6400;
    2470: romdata_int <= 'h4e21;
    2471: romdata_int <= 'h305a;
    2472: romdata_int <= 'h448; // Line Descriptor
    2473: romdata_int <= 'h6600;
    2474: romdata_int <= 'h695a;
    2475: romdata_int <= 'h8556;
    2476: romdata_int <= 'h448; // Line Descriptor
    2477: romdata_int <= 'h6800;
    2478: romdata_int <= 'h56c8;
    2479: romdata_int <= 'h407a;
    2480: romdata_int <= 'h448; // Line Descriptor
    2481: romdata_int <= 'h6a00;
    2482: romdata_int <= 'h1c60;
    2483: romdata_int <= 'h8611;
    2484: romdata_int <= 'h448; // Line Descriptor
    2485: romdata_int <= 'h6c00;
    2486: romdata_int <= 'h2256;
    2487: romdata_int <= 'h8d20;
    2488: romdata_int <= 'h448; // Line Descriptor
    2489: romdata_int <= 'h6e00;
    2490: romdata_int <= 'h26c1;
    2491: romdata_int <= 'h5e38;
    2492: romdata_int <= 'h448; // Line Descriptor
    2493: romdata_int <= 'h7000;
    2494: romdata_int <= 'h553;
    2495: romdata_int <= 'h28b7;
    2496: romdata_int <= 'h448; // Line Descriptor
    2497: romdata_int <= 'h7200;
    2498: romdata_int <= 'h52bb;
    2499: romdata_int <= 'h8a54;
    2500: romdata_int <= 'h448; // Line Descriptor
    2501: romdata_int <= 'h7400;
    2502: romdata_int <= 'ha89;
    2503: romdata_int <= 'h1872;
    2504: romdata_int <= 'h448; // Line Descriptor
    2505: romdata_int <= 'h7600;
    2506: romdata_int <= 'h7415;
    2507: romdata_int <= 'h8853;
    2508: romdata_int <= 'h448; // Line Descriptor
    2509: romdata_int <= 'h7800;
    2510: romdata_int <= 'h966;
    2511: romdata_int <= 'h46f1;
    2512: romdata_int <= 'h448; // Line Descriptor
    2513: romdata_int <= 'h7a00;
    2514: romdata_int <= 'hf1f;
    2515: romdata_int <= 'h35a;
    2516: romdata_int <= 'h448; // Line Descriptor
    2517: romdata_int <= 'h7c00;
    2518: romdata_int <= 'hd55;
    2519: romdata_int <= 'h8f1d;
    2520: romdata_int <= 'h448; // Line Descriptor
    2521: romdata_int <= 'h7e00;
    2522: romdata_int <= 'h24ac;
    2523: romdata_int <= 'h3c33;
    2524: romdata_int <= 'h448; // Line Descriptor
    2525: romdata_int <= 'h8000;
    2526: romdata_int <= 'h4473;
    2527: romdata_int <= 'h7a12;
    2528: romdata_int <= 'h448; // Line Descriptor
    2529: romdata_int <= 'h8200;
    2530: romdata_int <= 'h6f16;
    2531: romdata_int <= 'hcb;
    2532: romdata_int <= 'h448; // Line Descriptor
    2533: romdata_int <= 'h8400;
    2534: romdata_int <= 'h2cec;
    2535: romdata_int <= 'h2033;
    2536: romdata_int <= 'h448; // Line Descriptor
    2537: romdata_int <= 'h8600;
    2538: romdata_int <= 'h4b13;
    2539: romdata_int <= 'h140d;
    2540: romdata_int <= 'h448; // Line Descriptor
    2541: romdata_int <= 'h8800;
    2542: romdata_int <= 'h6d3;
    2543: romdata_int <= 'h50a8;
    2544: romdata_int <= 'h448; // Line Descriptor
    2545: romdata_int <= 'h8a00;
    2546: romdata_int <= 'h6c6b;
    2547: romdata_int <= 'h713c;
    2548: romdata_int <= 'h448; // Line Descriptor
    2549: romdata_int <= 'h8c00;
    2550: romdata_int <= 'h4831;
    2551: romdata_int <= 'h5a28;
    2552: romdata_int <= 'h548; // Line Descriptor
    2553: romdata_int <= 'h8e00;
    2554: romdata_int <= 'h642f;
    2555: romdata_int <= 'h826b;
    2556: romdata_int <= 'h183c; // Line Descriptor
    2557: romdata_int <= 'h0;
    2558: romdata_int <= 'h66ae;
    2559: romdata_int <= 'h2f0b;
    2560: romdata_int <= 'h3408;
    2561: romdata_int <= 'h5cd5;
    2562: romdata_int <= 'h3286;
    2563: romdata_int <= 'hc89;
    2564: romdata_int <= 'he2e;
    2565: romdata_int <= 'h4;
    2566: romdata_int <= 'h1b37;
    2567: romdata_int <= 'h4e9a;
    2568: romdata_int <= 'h26b0;
    2569: romdata_int <= 'h615c;
    2570: romdata_int <= 'h183c; // Line Descriptor
    2571: romdata_int <= 'h200;
    2572: romdata_int <= 'h7728;
    2573: romdata_int <= 'h428a;
    2574: romdata_int <= 'h1a6b;
    2575: romdata_int <= 'h5867;
    2576: romdata_int <= 'h2855;
    2577: romdata_int <= 'h861;
    2578: romdata_int <= 'h40d5;
    2579: romdata_int <= 'h371e;
    2580: romdata_int <= 'h50a5;
    2581: romdata_int <= 'hee0;
    2582: romdata_int <= 'h32e6;
    2583: romdata_int <= 'h734;
    2584: romdata_int <= 'h183c; // Line Descriptor
    2585: romdata_int <= 'h400;
    2586: romdata_int <= 'h232b;
    2587: romdata_int <= 'h3064;
    2588: romdata_int <= 'h5290;
    2589: romdata_int <= 'h3936;
    2590: romdata_int <= 'h1cd5;
    2591: romdata_int <= 'h4662;
    2592: romdata_int <= 'h70f2;
    2593: romdata_int <= 'h64b6;
    2594: romdata_int <= 'h8c9;
    2595: romdata_int <= 'h4b54;
    2596: romdata_int <= 'h1e4a;
    2597: romdata_int <= 'h1677;
    2598: romdata_int <= 'h183c; // Line Descriptor
    2599: romdata_int <= 'h600;
    2600: romdata_int <= 'h4b49;
    2601: romdata_int <= 'h667;
    2602: romdata_int <= 'h18a6;
    2603: romdata_int <= 'h20f2;
    2604: romdata_int <= 'h2c88;
    2605: romdata_int <= 'h6327;
    2606: romdata_int <= 'h2bd;
    2607: romdata_int <= 'h485c;
    2608: romdata_int <= 'h7648;
    2609: romdata_int <= 'h4522;
    2610: romdata_int <= 'h7301;
    2611: romdata_int <= 'h6934;
    2612: romdata_int <= 'h183c; // Line Descriptor
    2613: romdata_int <= 'h800;
    2614: romdata_int <= 'h3e4d;
    2615: romdata_int <= 'h1348;
    2616: romdata_int <= 'h601a;
    2617: romdata_int <= 'h760a;
    2618: romdata_int <= 'h3716;
    2619: romdata_int <= 'h6eee;
    2620: romdata_int <= 'h2e66;
    2621: romdata_int <= 'h7432;
    2622: romdata_int <= 'h4cf3;
    2623: romdata_int <= 'h1d2a;
    2624: romdata_int <= 'h5958;
    2625: romdata_int <= 'h3458;
    2626: romdata_int <= 'h183c; // Line Descriptor
    2627: romdata_int <= 'ha00;
    2628: romdata_int <= 'h74a2;
    2629: romdata_int <= 'h402a;
    2630: romdata_int <= 'h48c9;
    2631: romdata_int <= 'h12ce;
    2632: romdata_int <= 'h24fd;
    2633: romdata_int <= 'h3d19;
    2634: romdata_int <= 'h6650;
    2635: romdata_int <= 'h6233;
    2636: romdata_int <= 'h281c;
    2637: romdata_int <= 'hb38;
    2638: romdata_int <= 'h2221;
    2639: romdata_int <= 'h5508;
    2640: romdata_int <= 'h183c; // Line Descriptor
    2641: romdata_int <= 'hc00;
    2642: romdata_int <= 'hc08;
    2643: romdata_int <= 'h6665;
    2644: romdata_int <= 'h6e5;
    2645: romdata_int <= 'h22c0;
    2646: romdata_int <= 'h165d;
    2647: romdata_int <= 'h6a7b;
    2648: romdata_int <= 'h5efd;
    2649: romdata_int <= 'h5aeb;
    2650: romdata_int <= 'h5618;
    2651: romdata_int <= 'h5e40;
    2652: romdata_int <= 'h3f22;
    2653: romdata_int <= 'h14cf;
    2654: romdata_int <= 'h183c; // Line Descriptor
    2655: romdata_int <= 'he00;
    2656: romdata_int <= 'hf58;
    2657: romdata_int <= 'h3eee;
    2658: romdata_int <= 'h44c3;
    2659: romdata_int <= 'h5045;
    2660: romdata_int <= 'h1487;
    2661: romdata_int <= 'ha5c;
    2662: romdata_int <= 'h2aca;
    2663: romdata_int <= 'h5306;
    2664: romdata_int <= 'h337;
    2665: romdata_int <= 'h2b33;
    2666: romdata_int <= 'h12b0;
    2667: romdata_int <= 'h4088;
    2668: romdata_int <= 'h183c; // Line Descriptor
    2669: romdata_int <= 'h1000;
    2670: romdata_int <= 'h163f;
    2671: romdata_int <= 'h76f5;
    2672: romdata_int <= 'h30fe;
    2673: romdata_int <= 'h754b;
    2674: romdata_int <= 'h68a8;
    2675: romdata_int <= 'h497;
    2676: romdata_int <= 'h64a6;
    2677: romdata_int <= 'hcd5;
    2678: romdata_int <= 'h6eb1;
    2679: romdata_int <= 'h2ca1;
    2680: romdata_int <= 'h5d40;
    2681: romdata_int <= 'h6c5a;
    2682: romdata_int <= 'h183c; // Line Descriptor
    2683: romdata_int <= 'h1200;
    2684: romdata_int <= 'h3345;
    2685: romdata_int <= 'ha9e;
    2686: romdata_int <= 'h4a81;
    2687: romdata_int <= 'h274d;
    2688: romdata_int <= 'h4c8b;
    2689: romdata_int <= 'h3a99;
    2690: romdata_int <= 'h5634;
    2691: romdata_int <= 'h1951;
    2692: romdata_int <= 'h3c6f;
    2693: romdata_int <= 'h2513;
    2694: romdata_int <= 'h700b;
    2695: romdata_int <= 'h427a;
    2696: romdata_int <= 'h183c; // Line Descriptor
    2697: romdata_int <= 'h1400;
    2698: romdata_int <= 'h384c;
    2699: romdata_int <= 'h626f;
    2700: romdata_int <= 'h5550;
    2701: romdata_int <= 'h5ab5;
    2702: romdata_int <= 'h1e0f;
    2703: romdata_int <= 'h7247;
    2704: romdata_int <= 'h42b8;
    2705: romdata_int <= 'h20e2;
    2706: romdata_int <= 'h6b11;
    2707: romdata_int <= 'h1006;
    2708: romdata_int <= 'h383a;
    2709: romdata_int <= 'h6760;
    2710: romdata_int <= 'h183c; // Line Descriptor
    2711: romdata_int <= 'h1600;
    2712: romdata_int <= 'h40ea;
    2713: romdata_int <= 'h1a43;
    2714: romdata_int <= 'h4f4c;
    2715: romdata_int <= 'h10d2;
    2716: romdata_int <= 'h3e0a;
    2717: romdata_int <= 'h6d44;
    2718: romdata_int <= 'hec;
    2719: romdata_int <= 'h3a89;
    2720: romdata_int <= 'h2eaa;
    2721: romdata_int <= 'h3166;
    2722: romdata_int <= 'h46ce;
    2723: romdata_int <= 'h448;
    2724: romdata_int <= 'h43c; // Line Descriptor
    2725: romdata_int <= 'h1800;
    2726: romdata_int <= 'he6;
    2727: romdata_int <= 'h2ec;
    2728: romdata_int <= 'h43c; // Line Descriptor
    2729: romdata_int <= 'h1a00;
    2730: romdata_int <= 'h1031;
    2731: romdata_int <= 'h5ea0;
    2732: romdata_int <= 'h43c; // Line Descriptor
    2733: romdata_int <= 'h1c00;
    2734: romdata_int <= 'h6af4;
    2735: romdata_int <= 'hf0b;
    2736: romdata_int <= 'h43c; // Line Descriptor
    2737: romdata_int <= 'h1e00;
    2738: romdata_int <= 'h5d55;
    2739: romdata_int <= 'h54b8;
    2740: romdata_int <= 'h43c; // Line Descriptor
    2741: romdata_int <= 'h2000;
    2742: romdata_int <= 'h613;
    2743: romdata_int <= 'h2896;
    2744: romdata_int <= 'h43c; // Line Descriptor
    2745: romdata_int <= 'h2200;
    2746: romdata_int <= 'h2e1;
    2747: romdata_int <= 'h6c42;
    2748: romdata_int <= 'h43c; // Line Descriptor
    2749: romdata_int <= 'h2400;
    2750: romdata_int <= 'h6019;
    2751: romdata_int <= 'h3c24;
    2752: romdata_int <= 'h43c; // Line Descriptor
    2753: romdata_int <= 'h2600;
    2754: romdata_int <= 'h48cb;
    2755: romdata_int <= 'h2167;
    2756: romdata_int <= 'h43c; // Line Descriptor
    2757: romdata_int <= 'h2800;
    2758: romdata_int <= 'h6e22;
    2759: romdata_int <= 'h4b4b;
    2760: romdata_int <= 'h43c; // Line Descriptor
    2761: romdata_int <= 'h2a00;
    2762: romdata_int <= 'h6245;
    2763: romdata_int <= 'h4c84;
    2764: romdata_int <= 'h43c; // Line Descriptor
    2765: romdata_int <= 'h2c00;
    2766: romdata_int <= 'h5109;
    2767: romdata_int <= 'h38a7;
    2768: romdata_int <= 'h43c; // Line Descriptor
    2769: romdata_int <= 'h2e00;
    2770: romdata_int <= 'h4608;
    2771: romdata_int <= 'h1cd2;
    2772: romdata_int <= 'h43c; // Line Descriptor
    2773: romdata_int <= 'h3000;
    2774: romdata_int <= 'h528d;
    2775: romdata_int <= 'h648c;
    2776: romdata_int <= 'h43c; // Line Descriptor
    2777: romdata_int <= 'h3200;
    2778: romdata_int <= 'h1f25;
    2779: romdata_int <= 'h5917;
    2780: romdata_int <= 'h43c; // Line Descriptor
    2781: romdata_int <= 'h3400;
    2782: romdata_int <= 'h4262;
    2783: romdata_int <= 'h468d;
    2784: romdata_int <= 'h43c; // Line Descriptor
    2785: romdata_int <= 'h3600;
    2786: romdata_int <= 'h1d11;
    2787: romdata_int <= 'h56ad;
    2788: romdata_int <= 'h43c; // Line Descriptor
    2789: romdata_int <= 'h3800;
    2790: romdata_int <= 'h3a7b;
    2791: romdata_int <= 'h2a74;
    2792: romdata_int <= 'h43c; // Line Descriptor
    2793: romdata_int <= 'h3a00;
    2794: romdata_int <= 'h246f;
    2795: romdata_int <= 'h4f09;
    2796: romdata_int <= 'h43c; // Line Descriptor
    2797: romdata_int <= 'h3c00;
    2798: romdata_int <= 'h953;
    2799: romdata_int <= 'h36d8;
    2800: romdata_int <= 'h43c; // Line Descriptor
    2801: romdata_int <= 'h3e00;
    2802: romdata_int <= 'h6429;
    2803: romdata_int <= 'h10f3;
    2804: romdata_int <= 'h43c; // Line Descriptor
    2805: romdata_int <= 'h4000;
    2806: romdata_int <= 'h4d2a;
    2807: romdata_int <= 'h6e6e;
    2808: romdata_int <= 'h43c; // Line Descriptor
    2809: romdata_int <= 'h4200;
    2810: romdata_int <= 'h566f;
    2811: romdata_int <= 'h1744;
    2812: romdata_int <= 'h43c; // Line Descriptor
    2813: romdata_int <= 'h4400;
    2814: romdata_int <= 'h2008;
    2815: romdata_int <= 'h2246;
    2816: romdata_int <= 'h43c; // Line Descriptor
    2817: romdata_int <= 'h4600;
    2818: romdata_int <= 'h3c79;
    2819: romdata_int <= 'hc60;
    2820: romdata_int <= 'h43c; // Line Descriptor
    2821: romdata_int <= 'h4800;
    2822: romdata_int <= 'h2aaf;
    2823: romdata_int <= 'h5a94;
    2824: romdata_int <= 'h43c; // Line Descriptor
    2825: romdata_int <= 'h4a00;
    2826: romdata_int <= 'h4f53;
    2827: romdata_int <= 'h32c6;
    2828: romdata_int <= 'h43c; // Line Descriptor
    2829: romdata_int <= 'h4c00;
    2830: romdata_int <= 'h1444;
    2831: romdata_int <= 'h2461;
    2832: romdata_int <= 'h43c; // Line Descriptor
    2833: romdata_int <= 'h4e00;
    2834: romdata_int <= 'h53e;
    2835: romdata_int <= 'h11c;
    2836: romdata_int <= 'h43c; // Line Descriptor
    2837: romdata_int <= 'h5000;
    2838: romdata_int <= 'h1b51;
    2839: romdata_int <= 'h68cd;
    2840: romdata_int <= 'h43c; // Line Descriptor
    2841: romdata_int <= 'h5200;
    2842: romdata_int <= 'h5b42;
    2843: romdata_int <= 'h5d45;
    2844: romdata_int <= 'h43c; // Line Descriptor
    2845: romdata_int <= 'h5400;
    2846: romdata_int <= 'h1268;
    2847: romdata_int <= 'h153d;
    2848: romdata_int <= 'h43c; // Line Descriptor
    2849: romdata_int <= 'h5600;
    2850: romdata_int <= 'h72b7;
    2851: romdata_int <= 'h6b3f;
    2852: romdata_int <= 'h43c; // Line Descriptor
    2853: romdata_int <= 'h5800;
    2854: romdata_int <= 'h2949;
    2855: romdata_int <= 'h18c4;
    2856: romdata_int <= 'h43c; // Line Descriptor
    2857: romdata_int <= 'h5a00;
    2858: romdata_int <= 'h3147;
    2859: romdata_int <= 'h607b;
    2860: romdata_int <= 'h43c; // Line Descriptor
    2861: romdata_int <= 'h5c00;
    2862: romdata_int <= 'h710b;
    2863: romdata_int <= 'h523a;
    2864: romdata_int <= 'h43c; // Line Descriptor
    2865: romdata_int <= 'h5e00;
    2866: romdata_int <= 'h26c4;
    2867: romdata_int <= 'h55f;
    2868: romdata_int <= 'h43c; // Line Descriptor
    2869: romdata_int <= 'h6000;
    2870: romdata_int <= 'h54d9;
    2871: romdata_int <= 'h2ca1;
    2872: romdata_int <= 'h43c; // Line Descriptor
    2873: romdata_int <= 'h6200;
    2874: romdata_int <= 'h6c94;
    2875: romdata_int <= 'h7256;
    2876: romdata_int <= 'h43c; // Line Descriptor
    2877: romdata_int <= 'h6400;
    2878: romdata_int <= 'h5eb8;
    2879: romdata_int <= 'h2637;
    2880: romdata_int <= 'h43c; // Line Descriptor
    2881: romdata_int <= 'h6600;
    2882: romdata_int <= 'h693a;
    2883: romdata_int <= 'h4848;
    2884: romdata_int <= 'h43c; // Line Descriptor
    2885: romdata_int <= 'h6800;
    2886: romdata_int <= 'h4483;
    2887: romdata_int <= 'h7440;
    2888: romdata_int <= 'h43c; // Line Descriptor
    2889: romdata_int <= 'h6a00;
    2890: romdata_int <= 'h2e63;
    2891: romdata_int <= 'h5048;
    2892: romdata_int <= 'h43c; // Line Descriptor
    2893: romdata_int <= 'h6c00;
    2894: romdata_int <= 'h347a;
    2895: romdata_int <= 'h34c3;
    2896: romdata_int <= 'h43c; // Line Descriptor
    2897: romdata_int <= 'h6e00;
    2898: romdata_int <= 'h2c56;
    2899: romdata_int <= 'h3a5d;
    2900: romdata_int <= 'h43c; // Line Descriptor
    2901: romdata_int <= 'h7000;
    2902: romdata_int <= 'h1828;
    2903: romdata_int <= 'h1f20;
    2904: romdata_int <= 'h43c; // Line Descriptor
    2905: romdata_int <= 'h7200;
    2906: romdata_int <= 'haa4;
    2907: romdata_int <= 'h4555;
    2908: romdata_int <= 'h43c; // Line Descriptor
    2909: romdata_int <= 'h7400;
    2910: romdata_int <= 'h366f;
    2911: romdata_int <= 'h81f;
    2912: romdata_int <= 'h43c; // Line Descriptor
    2913: romdata_int <= 'h7600;
    2914: romdata_int <= 'h5956;
    2915: romdata_int <= 'h7056;
    2916: romdata_int <= 'h43c; // Line Descriptor
    2917: romdata_int <= 'h0;
    2918: romdata_int <= 'h5d2f;
    2919: romdata_int <= 'h5f1e;
    2920: romdata_int <= 'h43c; // Line Descriptor
    2921: romdata_int <= 'h200;
    2922: romdata_int <= 'h289c;
    2923: romdata_int <= 'h5c89;
    2924: romdata_int <= 'h43c; // Line Descriptor
    2925: romdata_int <= 'h400;
    2926: romdata_int <= 'h6a75;
    2927: romdata_int <= 'ha33;
    2928: romdata_int <= 'h43c; // Line Descriptor
    2929: romdata_int <= 'h600;
    2930: romdata_int <= 'h1930;
    2931: romdata_int <= 'h72df;
    2932: romdata_int <= 'h43c; // Line Descriptor
    2933: romdata_int <= 'h800;
    2934: romdata_int <= 'h5298;
    2935: romdata_int <= 'h5504;
    2936: romdata_int <= 'h43c; // Line Descriptor
    2937: romdata_int <= 'ha00;
    2938: romdata_int <= 'h44b2;
    2939: romdata_int <= 'h1aa9;
    2940: romdata_int <= 'h43c; // Line Descriptor
    2941: romdata_int <= 'hc00;
    2942: romdata_int <= 'hac1;
    2943: romdata_int <= 'h2497;
    2944: romdata_int <= 'h43c; // Line Descriptor
    2945: romdata_int <= 'he00;
    2946: romdata_int <= 'h2659;
    2947: romdata_int <= 'h749c;
    2948: romdata_int <= 'h43c; // Line Descriptor
    2949: romdata_int <= 'h1000;
    2950: romdata_int <= 'h3096;
    2951: romdata_int <= 'h469e;
    2952: romdata_int <= 'h43c; // Line Descriptor
    2953: romdata_int <= 'h1200;
    2954: romdata_int <= 'hc14;
    2955: romdata_int <= 'h4510;
    2956: romdata_int <= 'h43c; // Line Descriptor
    2957: romdata_int <= 'h1400;
    2958: romdata_int <= 'h6cf9;
    2959: romdata_int <= 'h2c12;
    2960: romdata_int <= 'h43c; // Line Descriptor
    2961: romdata_int <= 'h1600;
    2962: romdata_int <= 'h1e9c;
    2963: romdata_int <= 'h495a;
    2964: romdata_int <= 'h43c; // Line Descriptor
    2965: romdata_int <= 'h1800;
    2966: romdata_int <= 'h90a;
    2967: romdata_int <= 'h3664;
    2968: romdata_int <= 'h43c; // Line Descriptor
    2969: romdata_int <= 'h1a00;
    2970: romdata_int <= 'h3af6;
    2971: romdata_int <= 'h406b;
    2972: romdata_int <= 'h43c; // Line Descriptor
    2973: romdata_int <= 'h1c00;
    2974: romdata_int <= 'h2c85;
    2975: romdata_int <= 'h6735;
    2976: romdata_int <= 'h43c; // Line Descriptor
    2977: romdata_int <= 'h1e00;
    2978: romdata_int <= 'h54f5;
    2979: romdata_int <= 'h62ea;
    2980: romdata_int <= 'h43c; // Line Descriptor
    2981: romdata_int <= 'h2000;
    2982: romdata_int <= 'h1a04;
    2983: romdata_int <= 'h5a32;
    2984: romdata_int <= 'h43c; // Line Descriptor
    2985: romdata_int <= 'h2200;
    2986: romdata_int <= 'h1c15;
    2987: romdata_int <= 'h3541;
    2988: romdata_int <= 'h43c; // Line Descriptor
    2989: romdata_int <= 'h2400;
    2990: romdata_int <= 'h22f6;
    2991: romdata_int <= 'h822;
    2992: romdata_int <= 'h43c; // Line Descriptor
    2993: romdata_int <= 'h2600;
    2994: romdata_int <= 'he8;
    2995: romdata_int <= 'ha5;
    2996: romdata_int <= 'h43c; // Line Descriptor
    2997: romdata_int <= 'h2800;
    2998: romdata_int <= 'h4007;
    2999: romdata_int <= 'h6c7a;
    3000: romdata_int <= 'h43c; // Line Descriptor
    3001: romdata_int <= 'h2a00;
    3002: romdata_int <= 'h352f;
    3003: romdata_int <= 'h2aa5;
    3004: romdata_int <= 'h43c; // Line Descriptor
    3005: romdata_int <= 'h2c00;
    3006: romdata_int <= 'h1666;
    3007: romdata_int <= 'h1c5a;
    3008: romdata_int <= 'h43c; // Line Descriptor
    3009: romdata_int <= 'h2e00;
    3010: romdata_int <= 'h72a7;
    3011: romdata_int <= 'hca2;
    3012: romdata_int <= 'h43c; // Line Descriptor
    3013: romdata_int <= 'h3000;
    3014: romdata_int <= 'h5ac8;
    3015: romdata_int <= 'h265b;
    3016: romdata_int <= 'h43c; // Line Descriptor
    3017: romdata_int <= 'h3200;
    3018: romdata_int <= 'h448;
    3019: romdata_int <= 'h1485;
    3020: romdata_int <= 'h43c; // Line Descriptor
    3021: romdata_int <= 'h3400;
    3022: romdata_int <= 'h2104;
    3023: romdata_int <= 'h3c5c;
    3024: romdata_int <= 'h43c; // Line Descriptor
    3025: romdata_int <= 'h3600;
    3026: romdata_int <= 'h2b03;
    3027: romdata_int <= 'h52b1;
    3028: romdata_int <= 'h43c; // Line Descriptor
    3029: romdata_int <= 'h3800;
    3030: romdata_int <= 'h2559;
    3031: romdata_int <= 'he7b;
    3032: romdata_int <= 'h43c; // Line Descriptor
    3033: romdata_int <= 'h3a00;
    3034: romdata_int <= 'h7429;
    3035: romdata_int <= 'h3139;
    3036: romdata_int <= 'h43c; // Line Descriptor
    3037: romdata_int <= 'h3c00;
    3038: romdata_int <= 'h5895;
    3039: romdata_int <= 'h282b;
    3040: romdata_int <= 'h43c; // Line Descriptor
    3041: romdata_int <= 'h3e00;
    3042: romdata_int <= 'h486c;
    3043: romdata_int <= 'h3b2a;
    3044: romdata_int <= 'h43c; // Line Descriptor
    3045: romdata_int <= 'h4000;
    3046: romdata_int <= 'h60b9;
    3047: romdata_int <= 'h4c01;
    3048: romdata_int <= 'h43c; // Line Descriptor
    3049: romdata_int <= 'h4200;
    3050: romdata_int <= 'h4f56;
    3051: romdata_int <= 'h583d;
    3052: romdata_int <= 'h43c; // Line Descriptor
    3053: romdata_int <= 'h4400;
    3054: romdata_int <= 'h147d;
    3055: romdata_int <= 'h121a;
    3056: romdata_int <= 'h43c; // Line Descriptor
    3057: romdata_int <= 'h4600;
    3058: romdata_int <= 'h510a;
    3059: romdata_int <= 'h68c2;
    3060: romdata_int <= 'h43c; // Line Descriptor
    3061: romdata_int <= 'h4800;
    3062: romdata_int <= 'h3698;
    3063: romdata_int <= 'h56ab;
    3064: romdata_int <= 'h43c; // Line Descriptor
    3065: romdata_int <= 'h4a00;
    3066: romdata_int <= 'h3d15;
    3067: romdata_int <= 'h1603;
    3068: romdata_int <= 'h43c; // Line Descriptor
    3069: romdata_int <= 'h4c00;
    3070: romdata_int <= 'h4b03;
    3071: romdata_int <= 'h3337;
    3072: romdata_int <= 'h43c; // Line Descriptor
    3073: romdata_int <= 'h4e00;
    3074: romdata_int <= 'hf1e;
    3075: romdata_int <= 'h4b5c;
    3076: romdata_int <= 'h43c; // Line Descriptor
    3077: romdata_int <= 'h5000;
    3078: romdata_int <= 'h7046;
    3079: romdata_int <= 'h3e38;
    3080: romdata_int <= 'h43c; // Line Descriptor
    3081: romdata_int <= 'h5200;
    3082: romdata_int <= 'h694e;
    3083: romdata_int <= 'h771e;
    3084: romdata_int <= 'h43c; // Line Descriptor
    3085: romdata_int <= 'h5400;
    3086: romdata_int <= 'h4c99;
    3087: romdata_int <= 'h2054;
    3088: romdata_int <= 'h43c; // Line Descriptor
    3089: romdata_int <= 'h5600;
    3090: romdata_int <= 'h1333;
    3091: romdata_int <= 'h188d;
    3092: romdata_int <= 'h43c; // Line Descriptor
    3093: romdata_int <= 'h5800;
    3094: romdata_int <= 'h42c9;
    3095: romdata_int <= 'h6b59;
    3096: romdata_int <= 'h43c; // Line Descriptor
    3097: romdata_int <= 'h5a00;
    3098: romdata_int <= 'h3310;
    3099: romdata_int <= 'h38d4;
    3100: romdata_int <= 'h43c; // Line Descriptor
    3101: romdata_int <= 'h5c00;
    3102: romdata_int <= 'h70b;
    3103: romdata_int <= 'h6eb8;
    3104: romdata_int <= 'h43c; // Line Descriptor
    3105: romdata_int <= 'h5e00;
    3106: romdata_int <= 'h1054;
    3107: romdata_int <= 'h1f25;
    3108: romdata_int <= 'h43c; // Line Descriptor
    3109: romdata_int <= 'h6000;
    3110: romdata_int <= 'h473c;
    3111: romdata_int <= 'h2250;
    3112: romdata_int <= 'h43c; // Line Descriptor
    3113: romdata_int <= 'h6200;
    3114: romdata_int <= 'h5712;
    3115: romdata_int <= 'h703a;
    3116: romdata_int <= 'h43c; // Line Descriptor
    3117: romdata_int <= 'h6400;
    3118: romdata_int <= 'h7617;
    3119: romdata_int <= 'h110d;
    3120: romdata_int <= 'h43c; // Line Descriptor
    3121: romdata_int <= 'h6600;
    3122: romdata_int <= 'h23d;
    3123: romdata_int <= 'h4e32;
    3124: romdata_int <= 'h43c; // Line Descriptor
    3125: romdata_int <= 'h6800;
    3126: romdata_int <= 'h653c;
    3127: romdata_int <= 'h32e;
    3128: romdata_int <= 'h43c; // Line Descriptor
    3129: romdata_int <= 'h6a00;
    3130: romdata_int <= 'h3895;
    3131: romdata_int <= 'h42c4;
    3132: romdata_int <= 'h43c; // Line Descriptor
    3133: romdata_int <= 'h6c00;
    3134: romdata_int <= 'h5edf;
    3135: romdata_int <= 'h72c;
    3136: romdata_int <= 'h43c; // Line Descriptor
    3137: romdata_int <= 'h6e00;
    3138: romdata_int <= 'h2e58;
    3139: romdata_int <= 'h2e33;
    3140: romdata_int <= 'h43c; // Line Descriptor
    3141: romdata_int <= 'h7000;
    3142: romdata_int <= 'h6608;
    3143: romdata_int <= 'h6115;
    3144: romdata_int <= 'h43c; // Line Descriptor
    3145: romdata_int <= 'h7200;
    3146: romdata_int <= 'h3e4f;
    3147: romdata_int <= 'h470;
    3148: romdata_int <= 'h43c; // Line Descriptor
    3149: romdata_int <= 'h7400;
    3150: romdata_int <= 'h6e5e;
    3151: romdata_int <= 'h5084;
    3152: romdata_int <= 'h53c; // Line Descriptor
    3153: romdata_int <= 'h7600;
    3154: romdata_int <= 'h623b;
    3155: romdata_int <= 'h64f3;
    3156: romdata_int <= 'h162d; // Line Descriptor
    3157: romdata_int <= 'h0;
    3158: romdata_int <= 'h508d;
    3159: romdata_int <= 'h34af;
    3160: romdata_int <= 'h3f44;
    3161: romdata_int <= 'h3129;
    3162: romdata_int <= 'h50f8;
    3163: romdata_int <= 'h1848;
    3164: romdata_int <= 'h2e74;
    3165: romdata_int <= 'h3a37;
    3166: romdata_int <= 'h2c3c;
    3167: romdata_int <= 'h1612;
    3168: romdata_int <= 'h4ea3;
    3169: romdata_int <= 'h162d; // Line Descriptor
    3170: romdata_int <= 'h200;
    3171: romdata_int <= 'h26fc;
    3172: romdata_int <= 'h563b;
    3173: romdata_int <= 'h5407;
    3174: romdata_int <= 'h1333;
    3175: romdata_int <= 'h4b1b;
    3176: romdata_int <= 'h58a0;
    3177: romdata_int <= 'h496;
    3178: romdata_int <= 'h1554;
    3179: romdata_int <= 'h5412;
    3180: romdata_int <= 'h2a2c;
    3181: romdata_int <= 'h40fd;
    3182: romdata_int <= 'h162d; // Line Descriptor
    3183: romdata_int <= 'h400;
    3184: romdata_int <= 'h40ae;
    3185: romdata_int <= 'h18b1;
    3186: romdata_int <= 'h2a8c;
    3187: romdata_int <= 'h2d2e;
    3188: romdata_int <= 'h50f;
    3189: romdata_int <= 'h941;
    3190: romdata_int <= 'h2350;
    3191: romdata_int <= 'h134;
    3192: romdata_int <= 'h5625;
    3193: romdata_int <= 'h128e;
    3194: romdata_int <= 'h452a;
    3195: romdata_int <= 'h162d; // Line Descriptor
    3196: romdata_int <= 'h600;
    3197: romdata_int <= 'h3c22;
    3198: romdata_int <= 'h1d06;
    3199: romdata_int <= 'h9b;
    3200: romdata_int <= 'h2327;
    3201: romdata_int <= 'h251;
    3202: romdata_int <= 'h4054;
    3203: romdata_int <= 'h54c2;
    3204: romdata_int <= 'h20a2;
    3205: romdata_int <= 'h4680;
    3206: romdata_int <= 'h233e;
    3207: romdata_int <= 'h48ae;
    3208: romdata_int <= 'h162d; // Line Descriptor
    3209: romdata_int <= 'h800;
    3210: romdata_int <= 'h2aa9;
    3211: romdata_int <= 'h2cfd;
    3212: romdata_int <= 'h2744;
    3213: romdata_int <= 'h1cd7;
    3214: romdata_int <= 'h1024;
    3215: romdata_int <= 'h562e;
    3216: romdata_int <= 'h12f0;
    3217: romdata_int <= 'h1ace;
    3218: romdata_int <= 'h1e1b;
    3219: romdata_int <= 'h3f52;
    3220: romdata_int <= 'h146c;
    3221: romdata_int <= 'h162d; // Line Descriptor
    3222: romdata_int <= 'ha00;
    3223: romdata_int <= 'h4623;
    3224: romdata_int <= 'h3a7e;
    3225: romdata_int <= 'h4960;
    3226: romdata_int <= 'h52d1;
    3227: romdata_int <= 'hb16;
    3228: romdata_int <= 'ha1f;
    3229: romdata_int <= 'h68c;
    3230: romdata_int <= 'h1678;
    3231: romdata_int <= 'hd3b;
    3232: romdata_int <= 'h2935;
    3233: romdata_int <= 'h2ea3;
    3234: romdata_int <= 'h162d; // Line Descriptor
    3235: romdata_int <= 'hc00;
    3236: romdata_int <= 'h125a;
    3237: romdata_int <= 'h20c4;
    3238: romdata_int <= 'h3c4b;
    3239: romdata_int <= 'h2eae;
    3240: romdata_int <= 'h36b1;
    3241: romdata_int <= 'h4954;
    3242: romdata_int <= 'h3c84;
    3243: romdata_int <= 'h24e6;
    3244: romdata_int <= 'h24e4;
    3245: romdata_int <= 'hd7;
    3246: romdata_int <= 'h2067;
    3247: romdata_int <= 'h162d; // Line Descriptor
    3248: romdata_int <= 'he00;
    3249: romdata_int <= 'h3e62;
    3250: romdata_int <= 'h658;
    3251: romdata_int <= 'h24cb;
    3252: romdata_int <= 'h4e2e;
    3253: romdata_int <= 'h4d19;
    3254: romdata_int <= 'h44a5;
    3255: romdata_int <= 'h1f0b;
    3256: romdata_int <= 'h350f;
    3257: romdata_int <= 'h580d;
    3258: romdata_int <= 'h552;
    3259: romdata_int <= 'h209;
    3260: romdata_int <= 'h162d; // Line Descriptor
    3261: romdata_int <= 'h1000;
    3262: romdata_int <= 'h2c85;
    3263: romdata_int <= 'h52ba;
    3264: romdata_int <= 'h1680;
    3265: romdata_int <= 'h404d;
    3266: romdata_int <= 'h60c;
    3267: romdata_int <= 'h373b;
    3268: romdata_int <= 'h2813;
    3269: romdata_int <= 'hccc;
    3270: romdata_int <= 'h328a;
    3271: romdata_int <= 'h735;
    3272: romdata_int <= 'h104f;
    3273: romdata_int <= 'h162d; // Line Descriptor
    3274: romdata_int <= 'h1200;
    3275: romdata_int <= 'h4a47;
    3276: romdata_int <= 'h1493;
    3277: romdata_int <= 'h326a;
    3278: romdata_int <= 'hc0c;
    3279: romdata_int <= 'h20d9;
    3280: romdata_int <= 'h22e;
    3281: romdata_int <= 'h2ca2;
    3282: romdata_int <= 'h304b;
    3283: romdata_int <= 'haa1;
    3284: romdata_int <= 'h366d;
    3285: romdata_int <= 'hf19;
    3286: romdata_int <= 'h162d; // Line Descriptor
    3287: romdata_int <= 'h1400;
    3288: romdata_int <= 'hc4;
    3289: romdata_int <= 'h10e0;
    3290: romdata_int <= 'h28f6;
    3291: romdata_int <= 'h89d;
    3292: romdata_int <= 'h1e92;
    3293: romdata_int <= 'h4f23;
    3294: romdata_int <= 'h42e1;
    3295: romdata_int <= 'h389f;
    3296: romdata_int <= 'h4c0a;
    3297: romdata_int <= 'h3ca5;
    3298: romdata_int <= 'h1acd;
    3299: romdata_int <= 'h162d; // Line Descriptor
    3300: romdata_int <= 'h1600;
    3301: romdata_int <= 'h1a2a;
    3302: romdata_int <= 'h24f0;
    3303: romdata_int <= 'h3a02;
    3304: romdata_int <= 'h4604;
    3305: romdata_int <= 'h56a7;
    3306: romdata_int <= 'h2af5;
    3307: romdata_int <= 'h50eb;
    3308: romdata_int <= 'h3300;
    3309: romdata_int <= 'h3148;
    3310: romdata_int <= 'h52b0;
    3311: romdata_int <= 'h95b;
    3312: romdata_int <= 'h162d; // Line Descriptor
    3313: romdata_int <= 'h1800;
    3314: romdata_int <= 'h1451;
    3315: romdata_int <= 'hcc2;
    3316: romdata_int <= 'h186d;
    3317: romdata_int <= 'h4560;
    3318: romdata_int <= 'h5871;
    3319: romdata_int <= 'h262f;
    3320: romdata_int <= 'h1d62;
    3321: romdata_int <= 'h1148;
    3322: romdata_int <= 'h509e;
    3323: romdata_int <= 'h4a3b;
    3324: romdata_int <= 'h3a20;
    3325: romdata_int <= 'h162d; // Line Descriptor
    3326: romdata_int <= 'h1a00;
    3327: romdata_int <= 'h48b8;
    3328: romdata_int <= 'h5054;
    3329: romdata_int <= 'h140b;
    3330: romdata_int <= 'h1ac6;
    3331: romdata_int <= 'he96;
    3332: romdata_int <= 'h5211;
    3333: romdata_int <= 'h4ab0;
    3334: romdata_int <= 'h3e5d;
    3335: romdata_int <= 'h275a;
    3336: romdata_int <= 'h1d26;
    3337: romdata_int <= 'h183a;
    3338: romdata_int <= 'h162d; // Line Descriptor
    3339: romdata_int <= 'h1c00;
    3340: romdata_int <= 'h2541;
    3341: romdata_int <= 'h4a6b;
    3342: romdata_int <= 'h395d;
    3343: romdata_int <= 'h3443;
    3344: romdata_int <= 'h42f8;
    3345: romdata_int <= 'h471d;
    3346: romdata_int <= 'h4d2f;
    3347: romdata_int <= 'heb5;
    3348: romdata_int <= 'h3491;
    3349: romdata_int <= 'h434f;
    3350: romdata_int <= 'h38c2;
    3351: romdata_int <= 'h42d; // Line Descriptor
    3352: romdata_int <= 'h1e00;
    3353: romdata_int <= 'h5845;
    3354: romdata_int <= 'h170a;
    3355: romdata_int <= 'h42d; // Line Descriptor
    3356: romdata_int <= 'h2000;
    3357: romdata_int <= 'hd2a;
    3358: romdata_int <= 'h2a99;
    3359: romdata_int <= 'h42d; // Line Descriptor
    3360: romdata_int <= 'h2200;
    3361: romdata_int <= 'h723;
    3362: romdata_int <= 'h4128;
    3363: romdata_int <= 'h42d; // Line Descriptor
    3364: romdata_int <= 'h2400;
    3365: romdata_int <= 'h3a2c;
    3366: romdata_int <= 'h1f41;
    3367: romdata_int <= 'h42d; // Line Descriptor
    3368: romdata_int <= 'h2600;
    3369: romdata_int <= 'hea0;
    3370: romdata_int <= 'h4e5f;
    3371: romdata_int <= 'h42d; // Line Descriptor
    3372: romdata_int <= 'h2800;
    3373: romdata_int <= 'h3649;
    3374: romdata_int <= 'h3c57;
    3375: romdata_int <= 'h42d; // Line Descriptor
    3376: romdata_int <= 'h2a00;
    3377: romdata_int <= 'h1062;
    3378: romdata_int <= 'h4c8a;
    3379: romdata_int <= 'h42d; // Line Descriptor
    3380: romdata_int <= 'h2c00;
    3381: romdata_int <= 'h1c3b;
    3382: romdata_int <= 'h3336;
    3383: romdata_int <= 'h42d; // Line Descriptor
    3384: romdata_int <= 'h2e00;
    3385: romdata_int <= 'h16a8;
    3386: romdata_int <= 'h2ec8;
    3387: romdata_int <= 'h42d; // Line Descriptor
    3388: romdata_int <= 'h3000;
    3389: romdata_int <= 'h553a;
    3390: romdata_int <= 'h5441;
    3391: romdata_int <= 'h42d; // Line Descriptor
    3392: romdata_int <= 'h3200;
    3393: romdata_int <= 'h34a1;
    3394: romdata_int <= 'h389e;
    3395: romdata_int <= 'h42d; // Line Descriptor
    3396: romdata_int <= 'h3400;
    3397: romdata_int <= 'h1e88;
    3398: romdata_int <= 'h472f;
    3399: romdata_int <= 'h42d; // Line Descriptor
    3400: romdata_int <= 'h3600;
    3401: romdata_int <= 'h28a6;
    3402: romdata_int <= 'h3143;
    3403: romdata_int <= 'h42d; // Line Descriptor
    3404: romdata_int <= 'h3800;
    3405: romdata_int <= 'h22c0;
    3406: romdata_int <= 'h4836;
    3407: romdata_int <= 'h42d; // Line Descriptor
    3408: romdata_int <= 'h3a00;
    3409: romdata_int <= 'h8bf;
    3410: romdata_int <= 'h131d;
    3411: romdata_int <= 'h42d; // Line Descriptor
    3412: romdata_int <= 'h3c00;
    3413: romdata_int <= 'ha4d;
    3414: romdata_int <= 'h446;
    3415: romdata_int <= 'h42d; // Line Descriptor
    3416: romdata_int <= 'h3e00;
    3417: romdata_int <= 'h1935;
    3418: romdata_int <= 'h61;
    3419: romdata_int <= 'h42d; // Line Descriptor
    3420: romdata_int <= 'h4000;
    3421: romdata_int <= 'h4e85;
    3422: romdata_int <= 'hb31;
    3423: romdata_int <= 'h42d; // Line Descriptor
    3424: romdata_int <= 'h4200;
    3425: romdata_int <= 'h4cf3;
    3426: romdata_int <= 'hf3b;
    3427: romdata_int <= 'h42d; // Line Descriptor
    3428: romdata_int <= 'h4400;
    3429: romdata_int <= 'h4436;
    3430: romdata_int <= 'h3724;
    3431: romdata_int <= 'h42d; // Line Descriptor
    3432: romdata_int <= 'h4600;
    3433: romdata_int <= 'h2075;
    3434: romdata_int <= 'h274e;
    3435: romdata_int <= 'h42d; // Line Descriptor
    3436: romdata_int <= 'h4800;
    3437: romdata_int <= 'h2e18;
    3438: romdata_int <= 'h829;
    3439: romdata_int <= 'h42d; // Line Descriptor
    3440: romdata_int <= 'h4a00;
    3441: romdata_int <= 'h422d;
    3442: romdata_int <= 'h4417;
    3443: romdata_int <= 'h42d; // Line Descriptor
    3444: romdata_int <= 'h4c00;
    3445: romdata_int <= 'h30d6;
    3446: romdata_int <= 'h2887;
    3447: romdata_int <= 'h42d; // Line Descriptor
    3448: romdata_int <= 'h4e00;
    3449: romdata_int <= 'h33e;
    3450: romdata_int <= 'h22aa;
    3451: romdata_int <= 'h42d; // Line Descriptor
    3452: romdata_int <= 'h5000;
    3453: romdata_int <= 'h55b;
    3454: romdata_int <= 'h2b5;
    3455: romdata_int <= 'h42d; // Line Descriptor
    3456: romdata_int <= 'h5200;
    3457: romdata_int <= 'h5665;
    3458: romdata_int <= 'h1af9;
    3459: romdata_int <= 'h42d; // Line Descriptor
    3460: romdata_int <= 'h5400;
    3461: romdata_int <= 'h332f;
    3462: romdata_int <= 'h428a;
    3463: romdata_int <= 'h42d; // Line Descriptor
    3464: romdata_int <= 'h5600;
    3465: romdata_int <= 'h38be;
    3466: romdata_int <= 'h58ae;
    3467: romdata_int <= 'h42d; // Line Descriptor
    3468: romdata_int <= 'h5800;
    3469: romdata_int <= 'h5304;
    3470: romdata_int <= 'h3e3b;
    3471: romdata_int <= 'h42d; // Line Descriptor
    3472: romdata_int <= 'h0;
    3473: romdata_int <= 'h4016;
    3474: romdata_int <= 'h81c;
    3475: romdata_int <= 'h42d; // Line Descriptor
    3476: romdata_int <= 'h200;
    3477: romdata_int <= 'h918;
    3478: romdata_int <= 'h28dd;
    3479: romdata_int <= 'h42d; // Line Descriptor
    3480: romdata_int <= 'h400;
    3481: romdata_int <= 'h36b6;
    3482: romdata_int <= 'he3c;
    3483: romdata_int <= 'h42d; // Line Descriptor
    3484: romdata_int <= 'h600;
    3485: romdata_int <= 'hc46;
    3486: romdata_int <= 'h706;
    3487: romdata_int <= 'h42d; // Line Descriptor
    3488: romdata_int <= 'h800;
    3489: romdata_int <= 'h4e07;
    3490: romdata_int <= 'h3a21;
    3491: romdata_int <= 'h42d; // Line Descriptor
    3492: romdata_int <= 'ha00;
    3493: romdata_int <= 'h69b;
    3494: romdata_int <= 'h2538;
    3495: romdata_int <= 'h42d; // Line Descriptor
    3496: romdata_int <= 'hc00;
    3497: romdata_int <= 'h4b0;
    3498: romdata_int <= 'h1d65;
    3499: romdata_int <= 'h42d; // Line Descriptor
    3500: romdata_int <= 'he00;
    3501: romdata_int <= 'h194f;
    3502: romdata_int <= 'h430d;
    3503: romdata_int <= 'h42d; // Line Descriptor
    3504: romdata_int <= 'h1000;
    3505: romdata_int <= 'h1a70;
    3506: romdata_int <= 'h468f;
    3507: romdata_int <= 'h42d; // Line Descriptor
    3508: romdata_int <= 'h1200;
    3509: romdata_int <= 'h5519;
    3510: romdata_int <= 'h4b4b;
    3511: romdata_int <= 'h42d; // Line Descriptor
    3512: romdata_int <= 'h1400;
    3513: romdata_int <= 'h2f57;
    3514: romdata_int <= 'h1027;
    3515: romdata_int <= 'h42d; // Line Descriptor
    3516: romdata_int <= 'h1600;
    3517: romdata_int <= 'h2ab4;
    3518: romdata_int <= 'h1626;
    3519: romdata_int <= 'h42d; // Line Descriptor
    3520: romdata_int <= 'h1800;
    3521: romdata_int <= 'h1714;
    3522: romdata_int <= 'h120c;
    3523: romdata_int <= 'h42d; // Line Descriptor
    3524: romdata_int <= 'h1a00;
    3525: romdata_int <= 'h445b;
    3526: romdata_int <= 'h349d;
    3527: romdata_int <= 'h42d; // Line Descriptor
    3528: romdata_int <= 'h1c00;
    3529: romdata_int <= 'h3e1f;
    3530: romdata_int <= 'hbb;
    3531: romdata_int <= 'h42d; // Line Descriptor
    3532: romdata_int <= 'h1e00;
    3533: romdata_int <= 'h24d9;
    3534: romdata_int <= 'h58a8;
    3535: romdata_int <= 'h42d; // Line Descriptor
    3536: romdata_int <= 'h2000;
    3537: romdata_int <= 'h508b;
    3538: romdata_int <= 'h44fb;
    3539: romdata_int <= 'h42d; // Line Descriptor
    3540: romdata_int <= 'h2200;
    3541: romdata_int <= 'h1c1f;
    3542: romdata_int <= 'h30c;
    3543: romdata_int <= 'h42d; // Line Descriptor
    3544: romdata_int <= 'h2400;
    3545: romdata_int <= 'h14b3;
    3546: romdata_int <= 'h54c9;
    3547: romdata_int <= 'h42d; // Line Descriptor
    3548: romdata_int <= 'h2600;
    3549: romdata_int <= 'h4c40;
    3550: romdata_int <= 'h2ebb;
    3551: romdata_int <= 'h42d; // Line Descriptor
    3552: romdata_int <= 'h2800;
    3553: romdata_int <= 'h421c;
    3554: romdata_int <= 'h3d39;
    3555: romdata_int <= 'h42d; // Line Descriptor
    3556: romdata_int <= 'h2a00;
    3557: romdata_int <= 'he57;
    3558: romdata_int <= 'h4933;
    3559: romdata_int <= 'h42d; // Line Descriptor
    3560: romdata_int <= 'h2c00;
    3561: romdata_int <= 'h3455;
    3562: romdata_int <= 'h5058;
    3563: romdata_int <= 'h42d; // Line Descriptor
    3564: romdata_int <= 'h2e00;
    3565: romdata_int <= 'h1e82;
    3566: romdata_int <= 'h1a27;
    3567: romdata_int <= 'h42d; // Line Descriptor
    3568: romdata_int <= 'h3000;
    3569: romdata_int <= 'h3b;
    3570: romdata_int <= 'h234c;
    3571: romdata_int <= 'h42d; // Line Descriptor
    3572: romdata_int <= 'h3200;
    3573: romdata_int <= 'h3c7b;
    3574: romdata_int <= 'h408c;
    3575: romdata_int <= 'h42d; // Line Descriptor
    3576: romdata_int <= 'h3400;
    3577: romdata_int <= 'h385f;
    3578: romdata_int <= 'h3f18;
    3579: romdata_int <= 'h42d; // Line Descriptor
    3580: romdata_int <= 'h3600;
    3581: romdata_int <= 'h5702;
    3582: romdata_int <= 'h530f;
    3583: romdata_int <= 'h42d; // Line Descriptor
    3584: romdata_int <= 'h3800;
    3585: romdata_int <= 'hb64;
    3586: romdata_int <= 'h36a9;
    3587: romdata_int <= 'h42d; // Line Descriptor
    3588: romdata_int <= 'h3a00;
    3589: romdata_int <= 'h2867;
    3590: romdata_int <= 'h5739;
    3591: romdata_int <= 'h42d; // Line Descriptor
    3592: romdata_int <= 'h3c00;
    3593: romdata_int <= 'h58d4;
    3594: romdata_int <= 'h3923;
    3595: romdata_int <= 'h42d; // Line Descriptor
    3596: romdata_int <= 'h3e00;
    3597: romdata_int <= 'h4b36;
    3598: romdata_int <= 'h18d5;
    3599: romdata_int <= 'h42d; // Line Descriptor
    3600: romdata_int <= 'h4000;
    3601: romdata_int <= 'h2756;
    3602: romdata_int <= 'hb0d;
    3603: romdata_int <= 'h42d; // Line Descriptor
    3604: romdata_int <= 'h4200;
    3605: romdata_int <= 'h30c2;
    3606: romdata_int <= 'h1558;
    3607: romdata_int <= 'h42d; // Line Descriptor
    3608: romdata_int <= 'h4400;
    3609: romdata_int <= 'h48a4;
    3610: romdata_int <= 'h3354;
    3611: romdata_int <= 'h42d; // Line Descriptor
    3612: romdata_int <= 'h4600;
    3613: romdata_int <= 'h3a40;
    3614: romdata_int <= 'h3159;
    3615: romdata_int <= 'h42d; // Line Descriptor
    3616: romdata_int <= 'h4800;
    3617: romdata_int <= 'h3242;
    3618: romdata_int <= 'h2cb7;
    3619: romdata_int <= 'h42d; // Line Descriptor
    3620: romdata_int <= 'h4a00;
    3621: romdata_int <= 'h2d1;
    3622: romdata_int <= 'h2a6a;
    3623: romdata_int <= 'h42d; // Line Descriptor
    3624: romdata_int <= 'h4c00;
    3625: romdata_int <= 'h52f6;
    3626: romdata_int <= 'h4e6b;
    3627: romdata_int <= 'h42d; // Line Descriptor
    3628: romdata_int <= 'h4e00;
    3629: romdata_int <= 'h2c3e;
    3630: romdata_int <= 'h20bd;
    3631: romdata_int <= 'h42d; // Line Descriptor
    3632: romdata_int <= 'h5000;
    3633: romdata_int <= 'h20bc;
    3634: romdata_int <= 'h547;
    3635: romdata_int <= 'h42d; // Line Descriptor
    3636: romdata_int <= 'h5200;
    3637: romdata_int <= 'h46ad;
    3638: romdata_int <= 'h1f55;
    3639: romdata_int <= 'h42d; // Line Descriptor
    3640: romdata_int <= 'h5400;
    3641: romdata_int <= 'h121a;
    3642: romdata_int <= 'h26b0;
    3643: romdata_int <= 'h42d; // Line Descriptor
    3644: romdata_int <= 'h5600;
    3645: romdata_int <= 'h2234;
    3646: romdata_int <= 'h4cc0;
    3647: romdata_int <= 'h42d; // Line Descriptor
    3648: romdata_int <= 'h5800;
    3649: romdata_int <= 'h10ab;
    3650: romdata_int <= 'hc8a;
    3651: romdata_int <= 'h42d; // Line Descriptor
    3652: romdata_int <= 'h0;
    3653: romdata_int <= 'h184d;
    3654: romdata_int <= 'h49d;
    3655: romdata_int <= 'h42d; // Line Descriptor
    3656: romdata_int <= 'h200;
    3657: romdata_int <= 'h2057;
    3658: romdata_int <= 'h3d33;
    3659: romdata_int <= 'h42d; // Line Descriptor
    3660: romdata_int <= 'h400;
    3661: romdata_int <= 'h32aa;
    3662: romdata_int <= 'h3b1e;
    3663: romdata_int <= 'h42d; // Line Descriptor
    3664: romdata_int <= 'h600;
    3665: romdata_int <= 'h5826;
    3666: romdata_int <= 'h54b5;
    3667: romdata_int <= 'h42d; // Line Descriptor
    3668: romdata_int <= 'h800;
    3669: romdata_int <= 'had;
    3670: romdata_int <= 'ha1f;
    3671: romdata_int <= 'h42d; // Line Descriptor
    3672: romdata_int <= 'ha00;
    3673: romdata_int <= 'h42cc;
    3674: romdata_int <= 'h5282;
    3675: romdata_int <= 'h42d; // Line Descriptor
    3676: romdata_int <= 'hc00;
    3677: romdata_int <= 'h2637;
    3678: romdata_int <= 'h10ab;
    3679: romdata_int <= 'h42d; // Line Descriptor
    3680: romdata_int <= 'he00;
    3681: romdata_int <= 'h1639;
    3682: romdata_int <= 'h36af;
    3683: romdata_int <= 'h42d; // Line Descriptor
    3684: romdata_int <= 'h1000;
    3685: romdata_int <= 'hc6b;
    3686: romdata_int <= 'h2d5c;
    3687: romdata_int <= 'h42d; // Line Descriptor
    3688: romdata_int <= 'h1200;
    3689: romdata_int <= 'h3ee7;
    3690: romdata_int <= 'h1509;
    3691: romdata_int <= 'h42d; // Line Descriptor
    3692: romdata_int <= 'h1400;
    3693: romdata_int <= 'h1428;
    3694: romdata_int <= 'h814;
    3695: romdata_int <= 'h42d; // Line Descriptor
    3696: romdata_int <= 'h1600;
    3697: romdata_int <= 'h4afb;
    3698: romdata_int <= 'h4ecd;
    3699: romdata_int <= 'h42d; // Line Descriptor
    3700: romdata_int <= 'h1800;
    3701: romdata_int <= 'h22fb;
    3702: romdata_int <= 'h1e4f;
    3703: romdata_int <= 'h42d; // Line Descriptor
    3704: romdata_int <= 'h1a00;
    3705: romdata_int <= 'h2b4b;
    3706: romdata_int <= 'h503a;
    3707: romdata_int <= 'h42d; // Line Descriptor
    3708: romdata_int <= 'h1c00;
    3709: romdata_int <= 'h3aaa;
    3710: romdata_int <= 'h18ae;
    3711: romdata_int <= 'h42d; // Line Descriptor
    3712: romdata_int <= 'h1e00;
    3713: romdata_int <= 'h1c87;
    3714: romdata_int <= 'h4522;
    3715: romdata_int <= 'h42d; // Line Descriptor
    3716: romdata_int <= 'h2000;
    3717: romdata_int <= 'h2e57;
    3718: romdata_int <= 'hc3d;
    3719: romdata_int <= 'h42d; // Line Descriptor
    3720: romdata_int <= 'h2200;
    3721: romdata_int <= 'h8bd;
    3722: romdata_int <= 'h1a67;
    3723: romdata_int <= 'h42d; // Line Descriptor
    3724: romdata_int <= 'h2400;
    3725: romdata_int <= 'h130f;
    3726: romdata_int <= 'hec6;
    3727: romdata_int <= 'h42d; // Line Descriptor
    3728: romdata_int <= 'h2600;
    3729: romdata_int <= 'h447f;
    3730: romdata_int <= 'h2f14;
    3731: romdata_int <= 'h42d; // Line Descriptor
    3732: romdata_int <= 'h2800;
    3733: romdata_int <= 'h1b18;
    3734: romdata_int <= 'h2a62;
    3735: romdata_int <= 'h42d; // Line Descriptor
    3736: romdata_int <= 'h2a00;
    3737: romdata_int <= 'h4e1d;
    3738: romdata_int <= 'h1259;
    3739: romdata_int <= 'h42d; // Line Descriptor
    3740: romdata_int <= 'h2c00;
    3741: romdata_int <= 'h38bc;
    3742: romdata_int <= 'h4733;
    3743: romdata_int <= 'h42d; // Line Descriptor
    3744: romdata_int <= 'h2e00;
    3745: romdata_int <= 'h2826;
    3746: romdata_int <= 'h34b;
    3747: romdata_int <= 'h42d; // Line Descriptor
    3748: romdata_int <= 'h3000;
    3749: romdata_int <= 'h54c;
    3750: romdata_int <= 'h209e;
    3751: romdata_int <= 'h42d; // Line Descriptor
    3752: romdata_int <= 'h3200;
    3753: romdata_int <= 'h574c;
    3754: romdata_int <= 'h56c4;
    3755: romdata_int <= 'h42d; // Line Descriptor
    3756: romdata_int <= 'h3400;
    3757: romdata_int <= 'h1092;
    3758: romdata_int <= 'h1cbe;
    3759: romdata_int <= 'h42d; // Line Descriptor
    3760: romdata_int <= 'h3600;
    3761: romdata_int <= 'h546d;
    3762: romdata_int <= 'h4808;
    3763: romdata_int <= 'h42d; // Line Descriptor
    3764: romdata_int <= 'h3800;
    3765: romdata_int <= 'h3606;
    3766: romdata_int <= 'h331c;
    3767: romdata_int <= 'h42d; // Line Descriptor
    3768: romdata_int <= 'h3a00;
    3769: romdata_int <= 'h2534;
    3770: romdata_int <= 'h4094;
    3771: romdata_int <= 'h42d; // Line Descriptor
    3772: romdata_int <= 'h3c00;
    3773: romdata_int <= 'h2d07;
    3774: romdata_int <= 'h34f8;
    3775: romdata_int <= 'h42d; // Line Descriptor
    3776: romdata_int <= 'h3e00;
    3777: romdata_int <= 'h513f;
    3778: romdata_int <= 'h24ff;
    3779: romdata_int <= 'h42d; // Line Descriptor
    3780: romdata_int <= 'h4000;
    3781: romdata_int <= 'h4766;
    3782: romdata_int <= 'h1710;
    3783: romdata_int <= 'h42d; // Line Descriptor
    3784: romdata_int <= 'h4200;
    3785: romdata_int <= 'hf2b;
    3786: romdata_int <= 'h6a5;
    3787: romdata_int <= 'h42d; // Line Descriptor
    3788: romdata_int <= 'h4400;
    3789: romdata_int <= 'h4942;
    3790: romdata_int <= 'h3123;
    3791: romdata_int <= 'h42d; // Line Descriptor
    3792: romdata_int <= 'h4600;
    3793: romdata_int <= 'h1e38;
    3794: romdata_int <= 'h4cf9;
    3795: romdata_int <= 'h42d; // Line Descriptor
    3796: romdata_int <= 'h4800;
    3797: romdata_int <= 'h3c8f;
    3798: romdata_int <= 'h11a;
    3799: romdata_int <= 'h42d; // Line Descriptor
    3800: romdata_int <= 'h4a00;
    3801: romdata_int <= 'h4098;
    3802: romdata_int <= 'h26cf;
    3803: romdata_int <= 'h42d; // Line Descriptor
    3804: romdata_int <= 'h4c00;
    3805: romdata_int <= 'h3555;
    3806: romdata_int <= 'h3937;
    3807: romdata_int <= 'h42d; // Line Descriptor
    3808: romdata_int <= 'h4e00;
    3809: romdata_int <= 'h2b4;
    3810: romdata_int <= 'h22e2;
    3811: romdata_int <= 'h42d; // Line Descriptor
    3812: romdata_int <= 'h5000;
    3813: romdata_int <= 'h4d09;
    3814: romdata_int <= 'h426b;
    3815: romdata_int <= 'h42d; // Line Descriptor
    3816: romdata_int <= 'h5200;
    3817: romdata_int <= 'hb50;
    3818: romdata_int <= 'h5887;
    3819: romdata_int <= 'h42d; // Line Descriptor
    3820: romdata_int <= 'h5400;
    3821: romdata_int <= 'h52b2;
    3822: romdata_int <= 'h2941;
    3823: romdata_int <= 'h42d; // Line Descriptor
    3824: romdata_int <= 'h5600;
    3825: romdata_int <= 'h30f7;
    3826: romdata_int <= 'h4a72;
    3827: romdata_int <= 'h52d; // Line Descriptor
    3828: romdata_int <= 'h5800;
    3829: romdata_int <= 'h640;
    3830: romdata_int <= 'h3f42;
    3831: romdata_int <= 'h1424; // Line Descriptor
    3832: romdata_int <= 'h0;
    3833: romdata_int <= 'ha04;
    3834: romdata_int <= 'h2137;
    3835: romdata_int <= 'h3e9a;
    3836: romdata_int <= 'h30b0;
    3837: romdata_int <= 'h3f5c;
    3838: romdata_int <= 'h10e1;
    3839: romdata_int <= 'h12ec;
    3840: romdata_int <= 'h180b;
    3841: romdata_int <= 'h2516;
    3842: romdata_int <= 'h1964;
    3843: romdata_int <= 'h1424; // Line Descriptor
    3844: romdata_int <= 'h200;
    3845: romdata_int <= 'h2291;
    3846: romdata_int <= 'h2c0d;
    3847: romdata_int <= 'h2b28;
    3848: romdata_int <= 'h3c8a;
    3849: romdata_int <= 'h226b;
    3850: romdata_int <= 'h3467;
    3851: romdata_int <= 'h4055;
    3852: romdata_int <= 'h2261;
    3853: romdata_int <= 'h46d5;
    3854: romdata_int <= 'h131e;
    3855: romdata_int <= 'h1424; // Line Descriptor
    3856: romdata_int <= 'h400;
    3857: romdata_int <= 'h3cf2;
    3858: romdata_int <= 'h129a;
    3859: romdata_int <= 'h184e;
    3860: romdata_int <= 'h3ac4;
    3861: romdata_int <= 'h2950;
    3862: romdata_int <= 'h1323;
    3863: romdata_int <= 'h300f;
    3864: romdata_int <= 'h26d8;
    3865: romdata_int <= 'h2852;
    3866: romdata_int <= 'h423b;
    3867: romdata_int <= 'h1424; // Line Descriptor
    3868: romdata_int <= 'h600;
    3869: romdata_int <= 'h464a;
    3870: romdata_int <= 'h2877;
    3871: romdata_int <= 'h44e7;
    3872: romdata_int <= 'h3813;
    3873: romdata_int <= 'h424e;
    3874: romdata_int <= 'h145a;
    3875: romdata_int <= 'h1e83;
    3876: romdata_int <= 'h3318;
    3877: romdata_int <= 'h1a0e;
    3878: romdata_int <= 'h38d0;
    3879: romdata_int <= 'h1424; // Line Descriptor
    3880: romdata_int <= 'h800;
    3881: romdata_int <= 'hf4f;
    3882: romdata_int <= 'h2625;
    3883: romdata_int <= 'h94d;
    3884: romdata_int <= 'h2f52;
    3885: romdata_int <= 'h4738;
    3886: romdata_int <= 'h1a8f;
    3887: romdata_int <= 'h420e;
    3888: romdata_int <= 'h14ab;
    3889: romdata_int <= 'h4475;
    3890: romdata_int <= 'h2e41;
    3891: romdata_int <= 'h1424; // Line Descriptor
    3892: romdata_int <= 'ha00;
    3893: romdata_int <= 'h30bd;
    3894: romdata_int <= 'h1ec5;
    3895: romdata_int <= 'h63b;
    3896: romdata_int <= 'h2067;
    3897: romdata_int <= 'h269f;
    3898: romdata_int <= 'h3132;
    3899: romdata_int <= 'h392a;
    3900: romdata_int <= 'ha71;
    3901: romdata_int <= 'h61c;
    3902: romdata_int <= 'h45f;
    3903: romdata_int <= 'h1424; // Line Descriptor
    3904: romdata_int <= 'hc00;
    3905: romdata_int <= 'h3738;
    3906: romdata_int <= 'h3821;
    3907: romdata_int <= 'h2d08;
    3908: romdata_int <= 'h3428;
    3909: romdata_int <= 'h212c;
    3910: romdata_int <= 'h81a;
    3911: romdata_int <= 'h68;
    3912: romdata_int <= 'he4e;
    3913: romdata_int <= 'h2d3f;
    3914: romdata_int <= 'h2341;
    3915: romdata_int <= 'h1424; // Line Descriptor
    3916: romdata_int <= 'he00;
    3917: romdata_int <= 'h1a7e;
    3918: romdata_int <= 'h2f3f;
    3919: romdata_int <= 'h41f;
    3920: romdata_int <= 'h1c23;
    3921: romdata_int <= 'h1f46;
    3922: romdata_int <= 'h2e90;
    3923: romdata_int <= 'hcda;
    3924: romdata_int <= 'h2f63;
    3925: romdata_int <= 'h1e70;
    3926: romdata_int <= 'h8b4;
    3927: romdata_int <= 'h1424; // Line Descriptor
    3928: romdata_int <= 'h1000;
    3929: romdata_int <= 'hcea;
    3930: romdata_int <= 'h1672;
    3931: romdata_int <= 'h1106;
    3932: romdata_int <= 'h220b;
    3933: romdata_int <= 'h367b;
    3934: romdata_int <= 'h3c3e;
    3935: romdata_int <= 'h3edb;
    3936: romdata_int <= 'h2558;
    3937: romdata_int <= 'h16ee;
    3938: romdata_int <= 'h40c3;
    3939: romdata_int <= 'h1424; // Line Descriptor
    3940: romdata_int <= 'h1200;
    3941: romdata_int <= 'h426b;
    3942: romdata_int <= 'h24fd;
    3943: romdata_int <= 'h1a9d;
    3944: romdata_int <= 'ha7d;
    3945: romdata_int <= 'h641;
    3946: romdata_int <= 'h207;
    3947: romdata_int <= 'h3682;
    3948: romdata_int <= 'h4467;
    3949: romdata_int <= 'h3473;
    3950: romdata_int <= 'h102b;
    3951: romdata_int <= 'h1424; // Line Descriptor
    3952: romdata_int <= 'h1400;
    3953: romdata_int <= 'h182f;
    3954: romdata_int <= 'h10f8;
    3955: romdata_int <= 'hebc;
    3956: romdata_int <= 'h46ef;
    3957: romdata_int <= 'hee3;
    3958: romdata_int <= 'h44dc;
    3959: romdata_int <= 'h34e4;
    3960: romdata_int <= 'h4da;
    3961: romdata_int <= 'h36f6;
    3962: romdata_int <= 'h2f2;
    3963: romdata_int <= 'h1424; // Line Descriptor
    3964: romdata_int <= 'h1600;
    3965: romdata_int <= 'h2145;
    3966: romdata_int <= 'h3078;
    3967: romdata_int <= 'h1efc;
    3968: romdata_int <= 'h4138;
    3969: romdata_int <= 'hc3f;
    3970: romdata_int <= 'h18f5;
    3971: romdata_int <= 'h6fe;
    3972: romdata_int <= 'h1d4b;
    3973: romdata_int <= 'hca8;
    3974: romdata_int <= 'h2697;
    3975: romdata_int <= 'h1424; // Line Descriptor
    3976: romdata_int <= 'h1800;
    3977: romdata_int <= 'h1ecb;
    3978: romdata_int <= 'h146e;
    3979: romdata_int <= 'h431e;
    3980: romdata_int <= 'h143c;
    3981: romdata_int <= 'h24e5;
    3982: romdata_int <= 'h46b;
    3983: romdata_int <= 'h4639;
    3984: romdata_int <= 'h1766;
    3985: romdata_int <= 'h3b07;
    3986: romdata_int <= 'h145;
    3987: romdata_int <= 'h1424; // Line Descriptor
    3988: romdata_int <= 'h1a00;
    3989: romdata_int <= 'h347a;
    3990: romdata_int <= 'h3628;
    3991: romdata_int <= 'hc45;
    3992: romdata_int <= 'h12a2;
    3993: romdata_int <= 'h3216;
    3994: romdata_int <= 'hb3e;
    3995: romdata_int <= 'h3a0e;
    3996: romdata_int <= 'h2b37;
    3997: romdata_int <= 'h154c;
    3998: romdata_int <= 'h3e91;
    3999: romdata_int <= 'h1424; // Line Descriptor
    4000: romdata_int <= 'h1c00;
    4001: romdata_int <= 'h3a2a;
    4002: romdata_int <= 'h327d;
    4003: romdata_int <= 'h28dd;
    4004: romdata_int <= 'h260;
    4005: romdata_int <= 'h4108;
    4006: romdata_int <= 'h2ad6;
    4007: romdata_int <= 'h1069;
    4008: romdata_int <= 'h3c52;
    4009: romdata_int <= 'heaf;
    4010: romdata_int <= 'h2aa6;
    4011: romdata_int <= 'h1424; // Line Descriptor
    4012: romdata_int <= 'h1e00;
    4013: romdata_int <= 'h13f;
    4014: romdata_int <= 'h64c;
    4015: romdata_int <= 'h366f;
    4016: romdata_int <= 'h1750;
    4017: romdata_int <= 'hb5;
    4018: romdata_int <= 'h160f;
    4019: romdata_int <= 'h2047;
    4020: romdata_int <= 'h8b8;
    4021: romdata_int <= 'h1ce2;
    4022: romdata_int <= 'h3111;
    4023: romdata_int <= 'h1424; // Line Descriptor
    4024: romdata_int <= 'h2000;
    4025: romdata_int <= 'h2ca8;
    4026: romdata_int <= 'h4230;
    4027: romdata_int <= 'h2680;
    4028: romdata_int <= 'h24b5;
    4029: romdata_int <= 'h3adb;
    4030: romdata_int <= 'h2c67;
    4031: romdata_int <= 'h2d49;
    4032: romdata_int <= 'h1a32;
    4033: romdata_int <= 'h3d55;
    4034: romdata_int <= 'hae5;
    4035: romdata_int <= 'h1424; // Line Descriptor
    4036: romdata_int <= 'h2200;
    4037: romdata_int <= 'h2b59;
    4038: romdata_int <= 'h2298;
    4039: romdata_int <= 'hf3;
    4040: romdata_int <= 'h32d9;
    4041: romdata_int <= 'h38d4;
    4042: romdata_int <= 'h1c3a;
    4043: romdata_int <= 'h33b;
    4044: romdata_int <= 'h2851;
    4045: romdata_int <= 'h20ba;
    4046: romdata_int <= 'h334c;
    4047: romdata_int <= 'h424; // Line Descriptor
    4048: romdata_int <= 'h2400;
    4049: romdata_int <= 'h71a;
    4050: romdata_int <= 'h4474;
    4051: romdata_int <= 'h424; // Line Descriptor
    4052: romdata_int <= 'h2600;
    4053: romdata_int <= 'h41c;
    4054: romdata_int <= 'hf23;
    4055: romdata_int <= 'h424; // Line Descriptor
    4056: romdata_int <= 'h2800;
    4057: romdata_int <= 'h10f7;
    4058: romdata_int <= 'h351c;
    4059: romdata_int <= 'h424; // Line Descriptor
    4060: romdata_int <= 'h2a00;
    4061: romdata_int <= 'h271c;
    4062: romdata_int <= 'h555;
    4063: romdata_int <= 'h424; // Line Descriptor
    4064: romdata_int <= 'h2c00;
    4065: romdata_int <= 'h1cc4;
    4066: romdata_int <= 'ha7a;
    4067: romdata_int <= 'h424; // Line Descriptor
    4068: romdata_int <= 'h2e00;
    4069: romdata_int <= 'h3f54;
    4070: romdata_int <= 'h466b;
    4071: romdata_int <= 'h424; // Line Descriptor
    4072: romdata_int <= 'h3000;
    4073: romdata_int <= 'h394c;
    4074: romdata_int <= 'h40bd;
    4075: romdata_int <= 'h424; // Line Descriptor
    4076: romdata_int <= 'h3200;
    4077: romdata_int <= 'h1508;
    4078: romdata_int <= 'h79;
    4079: romdata_int <= 'h424; // Line Descriptor
    4080: romdata_int <= 'h3400;
    4081: romdata_int <= 'h12c6;
    4082: romdata_int <= 'h2b1d;
    4083: romdata_int <= 'h424; // Line Descriptor
    4084: romdata_int <= 'h3600;
    4085: romdata_int <= 'h34a;
    4086: romdata_int <= 'hc46;
    4087: romdata_int <= 'h424; // Line Descriptor
    4088: romdata_int <= 'h3800;
    4089: romdata_int <= 'h3236;
    4090: romdata_int <= 'h3b3e;
    4091: romdata_int <= 'h424; // Line Descriptor
    4092: romdata_int <= 'h3a00;
    4093: romdata_int <= 'h2854;
    4094: romdata_int <= 'h1b2f;
    4095: romdata_int <= 'h424; // Line Descriptor
    4096: romdata_int <= 'h3c00;
    4097: romdata_int <= 'h83e;
    4098: romdata_int <= 'h18f2;
    4099: romdata_int <= 'h424; // Line Descriptor
    4100: romdata_int <= 'h3e00;
    4101: romdata_int <= 'h40fc;
    4102: romdata_int <= 'h8b0;
    4103: romdata_int <= 'h424; // Line Descriptor
    4104: romdata_int <= 'h4000;
    4105: romdata_int <= 'h44cb;
    4106: romdata_int <= 'h1cee;
    4107: romdata_int <= 'h424; // Line Descriptor
    4108: romdata_int <= 'h4200;
    4109: romdata_int <= 'h1744;
    4110: romdata_int <= 'h321;
    4111: romdata_int <= 'h424; // Line Descriptor
    4112: romdata_int <= 'h4400;
    4113: romdata_int <= 'h2eb3;
    4114: romdata_int <= 'h3f62;
    4115: romdata_int <= 'h424; // Line Descriptor
    4116: romdata_int <= 'h4600;
    4117: romdata_int <= 'h2458;
    4118: romdata_int <= 'h3d52;
    4119: romdata_int <= 'h424; // Line Descriptor
    4120: romdata_int <= 'h0;
    4121: romdata_int <= 'h130b;
    4122: romdata_int <= 'h433d;
    4123: romdata_int <= 'h424; // Line Descriptor
    4124: romdata_int <= 'h200;
    4125: romdata_int <= 'h44cf;
    4126: romdata_int <= 'h3e9b;
    4127: romdata_int <= 'h424; // Line Descriptor
    4128: romdata_int <= 'h400;
    4129: romdata_int <= 'h4677;
    4130: romdata_int <= 'h2687;
    4131: romdata_int <= 'h424; // Line Descriptor
    4132: romdata_int <= 'h600;
    4133: romdata_int <= 'h3d;
    4134: romdata_int <= 'h2809;
    4135: romdata_int <= 'h424; // Line Descriptor
    4136: romdata_int <= 'h800;
    4137: romdata_int <= 'h6d1;
    4138: romdata_int <= 'h34b8;
    4139: romdata_int <= 'h424; // Line Descriptor
    4140: romdata_int <= 'ha00;
    4141: romdata_int <= 'h329;
    4142: romdata_int <= 'h3843;
    4143: romdata_int <= 'h424; // Line Descriptor
    4144: romdata_int <= 'hc00;
    4145: romdata_int <= 'h2ebb;
    4146: romdata_int <= 'hc4b;
    4147: romdata_int <= 'h424; // Line Descriptor
    4148: romdata_int <= 'he00;
    4149: romdata_int <= 'h408e;
    4150: romdata_int <= 'h2ca6;
    4151: romdata_int <= 'h424; // Line Descriptor
    4152: romdata_int <= 'h1000;
    4153: romdata_int <= 'h3732;
    4154: romdata_int <= 'hadf;
    4155: romdata_int <= 'h424; // Line Descriptor
    4156: romdata_int <= 'h1200;
    4157: romdata_int <= 'h2c86;
    4158: romdata_int <= 'he7b;
    4159: romdata_int <= 'h424; // Line Descriptor
    4160: romdata_int <= 'h1400;
    4161: romdata_int <= 'h2273;
    4162: romdata_int <= 'h1900;
    4163: romdata_int <= 'h424; // Line Descriptor
    4164: romdata_int <= 'h1600;
    4165: romdata_int <= 'h3d54;
    4166: romdata_int <= 'h14b6;
    4167: romdata_int <= 'h424; // Line Descriptor
    4168: romdata_int <= 'h1800;
    4169: romdata_int <= 'h54c;
    4170: romdata_int <= 'h40d2;
    4171: romdata_int <= 'h424; // Line Descriptor
    4172: romdata_int <= 'h1a00;
    4173: romdata_int <= 'h8ce;
    4174: romdata_int <= 'h48;
    4175: romdata_int <= 'h424; // Line Descriptor
    4176: romdata_int <= 'h1c00;
    4177: romdata_int <= 'h34f4;
    4178: romdata_int <= 'h310b;
    4179: romdata_int <= 'h424; // Line Descriptor
    4180: romdata_int <= 'h1e00;
    4181: romdata_int <= 'ha13;
    4182: romdata_int <= 'h3c96;
    4183: romdata_int <= 'h424; // Line Descriptor
    4184: romdata_int <= 'h2000;
    4185: romdata_int <= 'h2819;
    4186: romdata_int <= 'h1024;
    4187: romdata_int <= 'h424; // Line Descriptor
    4188: romdata_int <= 'h2200;
    4189: romdata_int <= 'h3a22;
    4190: romdata_int <= 'h254b;
    4191: romdata_int <= 'h424; // Line Descriptor
    4192: romdata_int <= 'h2400;
    4193: romdata_int <= 'h2709;
    4194: romdata_int <= 'h8a7;
    4195: romdata_int <= 'h424; // Line Descriptor
    4196: romdata_int <= 'h2600;
    4197: romdata_int <= 'h3008;
    4198: romdata_int <= 'h3ad2;
    4199: romdata_int <= 'h424; // Line Descriptor
    4200: romdata_int <= 'h2800;
    4201: romdata_int <= 'h167b;
    4202: romdata_int <= 'h2a74;
    4203: romdata_int <= 'h424; // Line Descriptor
    4204: romdata_int <= 'h2a00;
    4205: romdata_int <= 'hc6f;
    4206: romdata_int <= 'h1f09;
    4207: romdata_int <= 'h424; // Line Descriptor
    4208: romdata_int <= 'h2c00;
    4209: romdata_int <= 'h3953;
    4210: romdata_int <= 'h6d8;
    4211: romdata_int <= 'h424; // Line Descriptor
    4212: romdata_int <= 'h2e00;
    4213: romdata_int <= 'h2429;
    4214: romdata_int <= 'h44f3;
    4215: romdata_int <= 'h424; // Line Descriptor
    4216: romdata_int <= 'h3000;
    4217: romdata_int <= 'h2b2a;
    4218: romdata_int <= 'h126e;
    4219: romdata_int <= 'h424; // Line Descriptor
    4220: romdata_int <= 'h3200;
    4221: romdata_int <= 'h1879;
    4222: romdata_int <= 'h2e60;
    4223: romdata_int <= 'h424; // Line Descriptor
    4224: romdata_int <= 'h3400;
    4225: romdata_int <= 'h20af;
    4226: romdata_int <= 'h1c94;
    4227: romdata_int <= 'h424; // Line Descriptor
    4228: romdata_int <= 'h3600;
    4229: romdata_int <= 'he44;
    4230: romdata_int <= 'h261;
    4231: romdata_int <= 'h424; // Line Descriptor
    4232: romdata_int <= 'h3800;
    4233: romdata_int <= 'h3351;
    4234: romdata_int <= 'h32cd;
    4235: romdata_int <= 'h424; // Line Descriptor
    4236: romdata_int <= 'h3a00;
    4237: romdata_int <= 'h14b7;
    4238: romdata_int <= 'h173f;
    4239: romdata_int <= 'h424; // Line Descriptor
    4240: romdata_int <= 'h3c00;
    4241: romdata_int <= 'h4347;
    4242: romdata_int <= 'h367b;
    4243: romdata_int <= 'h424; // Line Descriptor
    4244: romdata_int <= 'h3e00;
    4245: romdata_int <= 'h1b0b;
    4246: romdata_int <= 'h43a;
    4247: romdata_int <= 'h424; // Line Descriptor
    4248: romdata_int <= 'h4000;
    4249: romdata_int <= 'h1e83;
    4250: romdata_int <= 'h2240;
    4251: romdata_int <= 'h424; // Line Descriptor
    4252: romdata_int <= 'h4200;
    4253: romdata_int <= 'h1c63;
    4254: romdata_int <= 'h2048;
    4255: romdata_int <= 'h424; // Line Descriptor
    4256: romdata_int <= 'h4400;
    4257: romdata_int <= 'h10ec;
    4258: romdata_int <= 'h1a33;
    4259: romdata_int <= 'h424; // Line Descriptor
    4260: romdata_int <= 'h4600;
    4261: romdata_int <= 'h3e6f;
    4262: romdata_int <= 'h461f;
    4263: romdata_int <= 'h424; // Line Descriptor
    4264: romdata_int <= 'h0;
    4265: romdata_int <= 'h3e9c;
    4266: romdata_int <= 'h689;
    4267: romdata_int <= 'h424; // Line Descriptor
    4268: romdata_int <= 'h200;
    4269: romdata_int <= 'he75;
    4270: romdata_int <= 'h4433;
    4271: romdata_int <= 'h424; // Line Descriptor
    4272: romdata_int <= 'h400;
    4273: romdata_int <= 'h3130;
    4274: romdata_int <= 'h34df;
    4275: romdata_int <= 'h424; // Line Descriptor
    4276: romdata_int <= 'h600;
    4277: romdata_int <= 'h2cc1;
    4278: romdata_int <= 'h1697;
    4279: romdata_int <= 'h424; // Line Descriptor
    4280: romdata_int <= 'h800;
    4281: romdata_int <= 'h1a59;
    4282: romdata_int <= 'h2c9c;
    4283: romdata_int <= 'h424; // Line Descriptor
    4284: romdata_int <= 'ha00;
    4285: romdata_int <= 'h10f9;
    4286: romdata_int <= 'h2a12;
    4287: romdata_int <= 'h424; // Line Descriptor
    4288: romdata_int <= 'hc00;
    4289: romdata_int <= 'h49c;
    4290: romdata_int <= 'h215a;
    4291: romdata_int <= 'h424; // Line Descriptor
    4292: romdata_int <= 'he00;
    4293: romdata_int <= 'h2228;
    4294: romdata_int <= 'h2823;
    4295: romdata_int <= 'h424; // Line Descriptor
    4296: romdata_int <= 'h1000;
    4297: romdata_int <= 'h18f6;
    4298: romdata_int <= 'h3e6b;
    4299: romdata_int <= 'h424; // Line Descriptor
    4300: romdata_int <= 'h1200;
    4301: romdata_int <= 'h14f6;
    4302: romdata_int <= 'h22;
    4303: romdata_int <= 'h424; // Line Descriptor
    4304: romdata_int <= 'h1400;
    4305: romdata_int <= 'h26e8;
    4306: romdata_int <= 'h40a5;
    4307: romdata_int <= 'h424; // Line Descriptor
    4308: romdata_int <= 'h1600;
    4309: romdata_int <= 'h1c07;
    4310: romdata_int <= 'h1a7a;
    4311: romdata_int <= 'h424; // Line Descriptor
    4312: romdata_int <= 'h1800;
    4313: romdata_int <= 'h4466;
    4314: romdata_int <= 'h85a;
    4315: romdata_int <= 'h424; // Line Descriptor
    4316: romdata_int <= 'h1a00;
    4317: romdata_int <= 'h36a7;
    4318: romdata_int <= 'h18a2;
    4319: romdata_int <= 'h424; // Line Descriptor
    4320: romdata_int <= 'h1c00;
    4321: romdata_int <= 'hc8;
    4322: romdata_int <= 'he5b;
    4323: romdata_int <= 'h424; // Line Descriptor
    4324: romdata_int <= 'h1e00;
    4325: romdata_int <= 'h3429;
    4326: romdata_int <= 'h1d39;
    4327: romdata_int <= 'h424; // Line Descriptor
    4328: romdata_int <= 'h2000;
    4329: romdata_int <= 'hd56;
    4330: romdata_int <= 'hc3d;
    4331: romdata_int <= 'h424; // Line Descriptor
    4332: romdata_int <= 'h2200;
    4333: romdata_int <= 'h2e7d;
    4334: romdata_int <= 'h3a1a;
    4335: romdata_int <= 'h424; // Line Descriptor
    4336: romdata_int <= 'h2400;
    4337: romdata_int <= 'h170a;
    4338: romdata_int <= 'h36c2;
    4339: romdata_int <= 'h424; // Line Descriptor
    4340: romdata_int <= 'h2600;
    4341: romdata_int <= 'h4046;
    4342: romdata_int <= 'h4638;
    4343: romdata_int <= 'h424; // Line Descriptor
    4344: romdata_int <= 'h2800;
    4345: romdata_int <= 'h2b4e;
    4346: romdata_int <= 'h151e;
    4347: romdata_int <= 'h424; // Line Descriptor
    4348: romdata_int <= 'h2a00;
    4349: romdata_int <= 'h2533;
    4350: romdata_int <= 'h388d;
    4351: romdata_int <= 'h424; // Line Descriptor
    4352: romdata_int <= 'h2c00;
    4353: romdata_int <= 'h6b8;
    4354: romdata_int <= 'h3cbf;
    4355: romdata_int <= 'h424; // Line Descriptor
    4356: romdata_int <= 'h2e00;
    4357: romdata_int <= 'h3312;
    4358: romdata_int <= 'h423a;
    4359: romdata_int <= 'h424; // Line Descriptor
    4360: romdata_int <= 'h3000;
    4361: romdata_int <= 'h217;
    4362: romdata_int <= 'h230d;
    4363: romdata_int <= 'h424; // Line Descriptor
    4364: romdata_int <= 'h3200;
    4365: romdata_int <= 'ha3d;
    4366: romdata_int <= 'h2632;
    4367: romdata_int <= 'h424; // Line Descriptor
    4368: romdata_int <= 'h3400;
    4369: romdata_int <= 'h3ab9;
    4370: romdata_int <= 'h367;
    4371: romdata_int <= 'h424; // Line Descriptor
    4372: romdata_int <= 'h3600;
    4373: romdata_int <= 'h1e3b;
    4374: romdata_int <= 'h12f3;
    4375: romdata_int <= 'h424; // Line Descriptor
    4376: romdata_int <= 'h3800;
    4377: romdata_int <= 'h214d;
    4378: romdata_int <= 'h10a5;
    4379: romdata_int <= 'h424; // Line Descriptor
    4380: romdata_int <= 'h3a00;
    4381: romdata_int <= 'h38f1;
    4382: romdata_int <= 'h2e58;
    4383: romdata_int <= 'h424; // Line Descriptor
    4384: romdata_int <= 'h3c00;
    4385: romdata_int <= 'h46e2;
    4386: romdata_int <= 'h332f;
    4387: romdata_int <= 'h424; // Line Descriptor
    4388: romdata_int <= 'h3e00;
    4389: romdata_int <= 'h42ae;
    4390: romdata_int <= 'h30c5;
    4391: romdata_int <= 'h424; // Line Descriptor
    4392: romdata_int <= 'h4000;
    4393: romdata_int <= 'h811;
    4394: romdata_int <= 'h24c6;
    4395: romdata_int <= 'h424; // Line Descriptor
    4396: romdata_int <= 'h4200;
    4397: romdata_int <= 'h3c8e;
    4398: romdata_int <= 'hb0f;
    4399: romdata_int <= 'h424; // Line Descriptor
    4400: romdata_int <= 'h4400;
    4401: romdata_int <= 'h1320;
    4402: romdata_int <= 'h4e2;
    4403: romdata_int <= 'h424; // Line Descriptor
    4404: romdata_int <= 'h4600;
    4405: romdata_int <= 'h28d3;
    4406: romdata_int <= 'h1ea1;
    4407: romdata_int <= 'h424; // Line Descriptor
    4408: romdata_int <= 'h0;
    4409: romdata_int <= 'h1aca;
    4410: romdata_int <= 'h4711;
    4411: romdata_int <= 'h424; // Line Descriptor
    4412: romdata_int <= 'h200;
    4413: romdata_int <= 'h30d7;
    4414: romdata_int <= 'h3f2d;
    4415: romdata_int <= 'h424; // Line Descriptor
    4416: romdata_int <= 'h400;
    4417: romdata_int <= 'h3f56;
    4418: romdata_int <= 'h26fa;
    4419: romdata_int <= 'h424; // Line Descriptor
    4420: romdata_int <= 'h600;
    4421: romdata_int <= 'h2c7a;
    4422: romdata_int <= 'h1ee7;
    4423: romdata_int <= 'h424; // Line Descriptor
    4424: romdata_int <= 'h800;
    4425: romdata_int <= 'h1060;
    4426: romdata_int <= 'h3c11;
    4427: romdata_int <= 'h424; // Line Descriptor
    4428: romdata_int <= 'ha00;
    4429: romdata_int <= 'h18c1;
    4430: romdata_int <= 'h2e38;
    4431: romdata_int <= 'h424; // Line Descriptor
    4432: romdata_int <= 'hc00;
    4433: romdata_int <= 'h3c15;
    4434: romdata_int <= 'h4253;
    4435: romdata_int <= 'h424; // Line Descriptor
    4436: romdata_int <= 'he00;
    4437: romdata_int <= 'h3413;
    4438: romdata_int <= 'h4439;
    4439: romdata_int <= 'h424; // Line Descriptor
    4440: romdata_int <= 'h1000;
    4441: romdata_int <= 'hece;
    4442: romdata_int <= 'h2a9b;
    4443: romdata_int <= 'h424; // Line Descriptor
    4444: romdata_int <= 'h1200;
    4445: romdata_int <= 'h28e1;
    4446: romdata_int <= 'h3287;
    4447: romdata_int <= 'h424; // Line Descriptor
    4448: romdata_int <= 'h1400;
    4449: romdata_int <= 'h358;
    4450: romdata_int <= 'h54d;
    4451: romdata_int <= 'h424; // Line Descriptor
    4452: romdata_int <= 'h1600;
    4453: romdata_int <= 'h270e;
    4454: romdata_int <= 'h3516;
    4455: romdata_int <= 'h424; // Line Descriptor
    4456: romdata_int <= 'h1800;
    4457: romdata_int <= 'h380b;
    4458: romdata_int <= 'h151a;
    4459: romdata_int <= 'h424; // Line Descriptor
    4460: romdata_int <= 'h1a00;
    4461: romdata_int <= 'h1e25;
    4462: romdata_int <= 'h2d3;
    4463: romdata_int <= 'h424; // Line Descriptor
    4464: romdata_int <= 'h1c00;
    4465: romdata_int <= 'h1428;
    4466: romdata_int <= 'h803;
    4467: romdata_int <= 'h424; // Line Descriptor
    4468: romdata_int <= 'h1e00;
    4469: romdata_int <= 'h12dd;
    4470: romdata_int <= 'h24eb;
    4471: romdata_int <= 'h424; // Line Descriptor
    4472: romdata_int <= 'h2000;
    4473: romdata_int <= 'h22f8;
    4474: romdata_int <= 'h22cd;
    4475: romdata_int <= 'h424; // Line Descriptor
    4476: romdata_int <= 'h2200;
    4477: romdata_int <= 'h4b7;
    4478: romdata_int <= 'he7;
    4479: romdata_int <= 'h424; // Line Descriptor
    4480: romdata_int <= 'h2400;
    4481: romdata_int <= 'h44bd;
    4482: romdata_int <= 'h16fa;
    4483: romdata_int <= 'h424; // Line Descriptor
    4484: romdata_int <= 'h2600;
    4485: romdata_int <= 'h24ab;
    4486: romdata_int <= 'h1d05;
    4487: romdata_int <= 'h424; // Line Descriptor
    4488: romdata_int <= 'h2800;
    4489: romdata_int <= 'h607;
    4490: romdata_int <= 'ha03;
    4491: romdata_int <= 'h424; // Line Descriptor
    4492: romdata_int <= 'h2a00;
    4493: romdata_int <= 'haac;
    4494: romdata_int <= 'h6a2;
    4495: romdata_int <= 'h424; // Line Descriptor
    4496: romdata_int <= 'h2c00;
    4497: romdata_int <= 'h1d66;
    4498: romdata_int <= 'h386a;
    4499: romdata_int <= 'h424; // Line Descriptor
    4500: romdata_int <= 'h2e00;
    4501: romdata_int <= 'h2a79;
    4502: romdata_int <= 'h1a61;
    4503: romdata_int <= 'h424; // Line Descriptor
    4504: romdata_int <= 'h3000;
    4505: romdata_int <= 'hc98;
    4506: romdata_int <= 'h40f0;
    4507: romdata_int <= 'h424; // Line Descriptor
    4508: romdata_int <= 'h3200;
    4509: romdata_int <= 'h327b;
    4510: romdata_int <= 'h103b;
    4511: romdata_int <= 'h424; // Line Descriptor
    4512: romdata_int <= 'h3400;
    4513: romdata_int <= 'h90e;
    4514: romdata_int <= 'h1826;
    4515: romdata_int <= 'h424; // Line Descriptor
    4516: romdata_int <= 'h3600;
    4517: romdata_int <= 'h4750;
    4518: romdata_int <= 'hd40;
    4519: romdata_int <= 'h424; // Line Descriptor
    4520: romdata_int <= 'h3800;
    4521: romdata_int <= 'h1756;
    4522: romdata_int <= 'hf08;
    4523: romdata_int <= 'h424; // Line Descriptor
    4524: romdata_int <= 'h3a00;
    4525: romdata_int <= 'h2ee4;
    4526: romdata_int <= 'h3030;
    4527: romdata_int <= 'h424; // Line Descriptor
    4528: romdata_int <= 'h3c00;
    4529: romdata_int <= 'h3a0d;
    4530: romdata_int <= 'h2cfa;
    4531: romdata_int <= 'h424; // Line Descriptor
    4532: romdata_int <= 'h3e00;
    4533: romdata_int <= 'h102;
    4534: romdata_int <= 'h2855;
    4535: romdata_int <= 'h424; // Line Descriptor
    4536: romdata_int <= 'h4000;
    4537: romdata_int <= 'h4244;
    4538: romdata_int <= 'h36d0;
    4539: romdata_int <= 'h424; // Line Descriptor
    4540: romdata_int <= 'h4200;
    4541: romdata_int <= 'h404a;
    4542: romdata_int <= 'h2007;
    4543: romdata_int <= 'h424; // Line Descriptor
    4544: romdata_int <= 'h4400;
    4545: romdata_int <= 'h366f;
    4546: romdata_int <= 'h3b56;
    4547: romdata_int <= 'h524; // Line Descriptor
    4548: romdata_int <= 'h4600;
    4549: romdata_int <= 'h20c5;
    4550: romdata_int <= 'h129a;
    4551: romdata_int <= 'h181e; // Line Descriptor
    4552: romdata_int <= 'h0;
    4553: romdata_int <= 'h1891;
    4554: romdata_int <= 'h340d;
    4555: romdata_int <= 'h3b28;
    4556: romdata_int <= 'h208a;
    4557: romdata_int <= 'hc6b;
    4558: romdata_int <= 'h2c67;
    4559: romdata_int <= 'h1455;
    4560: romdata_int <= 'h461;
    4561: romdata_int <= 'h1ed5;
    4562: romdata_int <= 'h1b1e;
    4563: romdata_int <= 'h26a5;
    4564: romdata_int <= 'h6e0;
    4565: romdata_int <= 'h181e; // Line Descriptor
    4566: romdata_int <= 'h200;
    4567: romdata_int <= 'h2652;
    4568: romdata_int <= 'h203b;
    4569: romdata_int <= 'h112b;
    4570: romdata_int <= 'h1664;
    4571: romdata_int <= 'h2690;
    4572: romdata_int <= 'h1b36;
    4573: romdata_int <= 'hed5;
    4574: romdata_int <= 'h2262;
    4575: romdata_int <= 'h38f2;
    4576: romdata_int <= 'h30b6;
    4577: romdata_int <= 'h2c9;
    4578: romdata_int <= 'h2354;
    4579: romdata_int <= 'h181e; // Line Descriptor
    4580: romdata_int <= 'h400;
    4581: romdata_int <= 'hb53;
    4582: romdata_int <= 'h132c;
    4583: romdata_int <= 'h2749;
    4584: romdata_int <= 'h267;
    4585: romdata_int <= 'haa6;
    4586: romdata_int <= 'hef2;
    4587: romdata_int <= 'h1888;
    4588: romdata_int <= 'h3127;
    4589: romdata_int <= 'h2bd;
    4590: romdata_int <= 'h225c;
    4591: romdata_int <= 'h3a48;
    4592: romdata_int <= 'h2122;
    4593: romdata_int <= 'h181e; // Line Descriptor
    4594: romdata_int <= 'h600;
    4595: romdata_int <= 'h2d2d;
    4596: romdata_int <= 'h329f;
    4597: romdata_int <= 'h3082;
    4598: romdata_int <= 'h1470;
    4599: romdata_int <= 'h114f;
    4600: romdata_int <= 'h2425;
    4601: romdata_int <= 'hd4d;
    4602: romdata_int <= 'h3352;
    4603: romdata_int <= 'h138;
    4604: romdata_int <= 'he8f;
    4605: romdata_int <= 'h1c0e;
    4606: romdata_int <= 'h10ab;
    4607: romdata_int <= 'h181e; // Line Descriptor
    4608: romdata_int <= 'h800;
    4609: romdata_int <= 'h124f;
    4610: romdata_int <= 'h905;
    4611: romdata_int <= 'haa1;
    4612: romdata_int <= 'h224d;
    4613: romdata_int <= 'h748;
    4614: romdata_int <= 'h301a;
    4615: romdata_int <= 'h3a0a;
    4616: romdata_int <= 'h1b16;
    4617: romdata_int <= 'h36ee;
    4618: romdata_int <= 'h1466;
    4619: romdata_int <= 'h3832;
    4620: romdata_int <= 'h2af3;
    4621: romdata_int <= 'h181e; // Line Descriptor
    4622: romdata_int <= 'ha00;
    4623: romdata_int <= 'h1e72;
    4624: romdata_int <= 'h1706;
    4625: romdata_int <= 'h240b;
    4626: romdata_int <= 'h67b;
    4627: romdata_int <= 'h203e;
    4628: romdata_int <= 'h1edb;
    4629: romdata_int <= 'h2958;
    4630: romdata_int <= 'h8ee;
    4631: romdata_int <= 'h28c3;
    4632: romdata_int <= 'h1c45;
    4633: romdata_int <= 'h487;
    4634: romdata_int <= 'h285c;
    4635: romdata_int <= 'h181e; // Line Descriptor
    4636: romdata_int <= 'hc00;
    4637: romdata_int <= 'h2282;
    4638: romdata_int <= 'h2a67;
    4639: romdata_int <= 'h3473;
    4640: romdata_int <= 'h1c2b;
    4641: romdata_int <= 'h1758;
    4642: romdata_int <= 'h3ac5;
    4643: romdata_int <= 'h12ad;
    4644: romdata_int <= 'h2a35;
    4645: romdata_int <= 'h1642;
    4646: romdata_int <= 'h1217;
    4647: romdata_int <= 'hd15;
    4648: romdata_int <= 'h14c;
    4649: romdata_int <= 'h181e; // Line Descriptor
    4650: romdata_int <= 'he00;
    4651: romdata_int <= 'h1ae5;
    4652: romdata_int <= 'h366b;
    4653: romdata_int <= 'he39;
    4654: romdata_int <= 'h1966;
    4655: romdata_int <= 'h307;
    4656: romdata_int <= 'h1d45;
    4657: romdata_int <= 'ha9e;
    4658: romdata_int <= 'h2481;
    4659: romdata_int <= 'h274d;
    4660: romdata_int <= 'hc8b;
    4661: romdata_int <= 'h3099;
    4662: romdata_int <= 'he34;
    4663: romdata_int <= 'h181e; // Line Descriptor
    4664: romdata_int <= 'h1000;
    4665: romdata_int <= 'h3760;
    4666: romdata_int <= 'ha49;
    4667: romdata_int <= 'h1238;
    4668: romdata_int <= 'h3862;
    4669: romdata_int <= 'h28b4;
    4670: romdata_int <= 'h56;
    4671: romdata_int <= 'h660;
    4672: romdata_int <= 'h20d8;
    4673: romdata_int <= 'h2a03;
    4674: romdata_int <= 'h2ec8;
    4675: romdata_int <= 'h822;
    4676: romdata_int <= 'h1294;
    4677: romdata_int <= 'h181e; // Line Descriptor
    4678: romdata_int <= 'h1200;
    4679: romdata_int <= 'hc7e;
    4680: romdata_int <= 'h1b1e;
    4681: romdata_int <= 'h845;
    4682: romdata_int <= 'h2a6e;
    4683: romdata_int <= 'h22a8;
    4684: romdata_int <= 'h1430;
    4685: romdata_int <= 'h80;
    4686: romdata_int <= 'h1cb5;
    4687: romdata_int <= 'h4db;
    4688: romdata_int <= 'h867;
    4689: romdata_int <= 'h2d49;
    4690: romdata_int <= 'h1832;
    4691: romdata_int <= 'h181e; // Line Descriptor
    4692: romdata_int <= 'h1400;
    4693: romdata_int <= 'h391c;
    4694: romdata_int <= 'h243d;
    4695: romdata_int <= 'h2d59;
    4696: romdata_int <= 'h3298;
    4697: romdata_int <= 'h2ef3;
    4698: romdata_int <= 'h34d9;
    4699: romdata_int <= 'h26d4;
    4700: romdata_int <= 'h343a;
    4701: romdata_int <= 'h193b;
    4702: romdata_int <= 'h3451;
    4703: romdata_int <= 'h34ba;
    4704: romdata_int <= 'h1f4c;
    4705: romdata_int <= 'h181e; // Line Descriptor
    4706: romdata_int <= 'h1600;
    4707: romdata_int <= 'h1d11;
    4708: romdata_int <= 'h761;
    4709: romdata_int <= 'h1f08;
    4710: romdata_int <= 'hc79;
    4711: romdata_int <= 'h1881;
    4712: romdata_int <= 'h80d;
    4713: romdata_int <= 'h38c6;
    4714: romdata_int <= 'h171d;
    4715: romdata_int <= 'h324f;
    4716: romdata_int <= 'h3af2;
    4717: romdata_int <= 'h3734;
    4718: romdata_int <= 'h254c;
    4719: romdata_int <= 'h181e; // Line Descriptor
    4720: romdata_int <= 'h1800;
    4721: romdata_int <= 'h3303;
    4722: romdata_int <= 'h1c02;
    4723: romdata_int <= 'h1a36;
    4724: romdata_int <= 'h53e;
    4725: romdata_int <= 'h36e4;
    4726: romdata_int <= 'h4f5;
    4727: romdata_int <= 'h36d5;
    4728: romdata_int <= 'h10fc;
    4729: romdata_int <= 'h762;
    4730: romdata_int <= 'ha18;
    4731: romdata_int <= 'h1654;
    4732: romdata_int <= 'h332f;
    4733: romdata_int <= 'h181e; // Line Descriptor
    4734: romdata_int <= 'h1a00;
    4735: romdata_int <= 'h16ee;
    4736: romdata_int <= 'h2c52;
    4737: romdata_int <= 'h8e;
    4738: romdata_int <= 'h2ea6;
    4739: romdata_int <= 'h3350;
    4740: romdata_int <= 'h12f7;
    4741: romdata_int <= 'h2f32;
    4742: romdata_int <= 'h2df;
    4743: romdata_int <= 'h1125;
    4744: romdata_int <= 'h2c45;
    4745: romdata_int <= 'h1b13;
    4746: romdata_int <= 'ha7d;
    4747: romdata_int <= 'h181e; // Line Descriptor
    4748: romdata_int <= 'h1c00;
    4749: romdata_int <= 'h78;
    4750: romdata_int <= 'h13;
    4751: romdata_int <= 'h3696;
    4752: romdata_int <= 'h2806;
    4753: romdata_int <= 'h3943;
    4754: romdata_int <= 'h2ae1;
    4755: romdata_int <= 'h1e42;
    4756: romdata_int <= 'h2d28;
    4757: romdata_int <= 'h20b5;
    4758: romdata_int <= 'h2419;
    4759: romdata_int <= 'h2e24;
    4760: romdata_int <= 'h14d9;
    4761: romdata_int <= 'h41e; // Line Descriptor
    4762: romdata_int <= 'h1e00;
    4763: romdata_int <= 'h8d2;
    4764: romdata_int <= 'h2fe;
    4765: romdata_int <= 'h41e; // Line Descriptor
    4766: romdata_int <= 'h2000;
    4767: romdata_int <= 'h24d8;
    4768: romdata_int <= 'h3b32;
    4769: romdata_int <= 'h41e; // Line Descriptor
    4770: romdata_int <= 'h2200;
    4771: romdata_int <= 'h6f3;
    4772: romdata_int <= 'hce2;
    4773: romdata_int <= 'h41e; // Line Descriptor
    4774: romdata_int <= 'h2400;
    4775: romdata_int <= 'h14c6;
    4776: romdata_int <= 'h3838;
    4777: romdata_int <= 'h41e; // Line Descriptor
    4778: romdata_int <= 'h2600;
    4779: romdata_int <= 'h31c;
    4780: romdata_int <= 'h2e3b;
    4781: romdata_int <= 'h41e; // Line Descriptor
    4782: romdata_int <= 'h2800;
    4783: romdata_int <= 'h30cd;
    4784: romdata_int <= 'h3105;
    4785: romdata_int <= 'h41e; // Line Descriptor
    4786: romdata_int <= 'h2a00;
    4787: romdata_int <= 'h2f45;
    4788: romdata_int <= 'h2827;
    4789: romdata_int <= 'h41e; // Line Descriptor
    4790: romdata_int <= 'h2c00;
    4791: romdata_int <= 'hf3d;
    4792: romdata_int <= 'h1156;
    4793: romdata_int <= 'h41e; // Line Descriptor
    4794: romdata_int <= 'h2e00;
    4795: romdata_int <= 'h2a48;
    4796: romdata_int <= 'h2737;
    4797: romdata_int <= 'h41e; // Line Descriptor
    4798: romdata_int <= 'h3000;
    4799: romdata_int <= 'h3a40;
    4800: romdata_int <= 'h14b9;
    4801: romdata_int <= 'h41e; // Line Descriptor
    4802: romdata_int <= 'h3200;
    4803: romdata_int <= 'h3433;
    4804: romdata_int <= 'h1e12;
    4805: romdata_int <= 'h41e; // Line Descriptor
    4806: romdata_int <= 'h3400;
    4807: romdata_int <= 'h291e;
    4808: romdata_int <= 'h227f;
    4809: romdata_int <= 'h41e; // Line Descriptor
    4810: romdata_int <= 'h3600;
    4811: romdata_int <= 'h4a9;
    4812: romdata_int <= 'he23;
    4813: romdata_int <= 'h41e; // Line Descriptor
    4814: romdata_int <= 'h3800;
    4815: romdata_int <= 'h1108;
    4816: romdata_int <= 'h476;
    4817: romdata_int <= 'h41e; // Line Descriptor
    4818: romdata_int <= 'h3a00;
    4819: romdata_int <= 'h206b;
    4820: romdata_int <= 'h187d;
    4821: romdata_int <= 'h41e; // Line Descriptor
    4822: romdata_int <= 'h0;
    4823: romdata_int <= 'h32ea;
    4824: romdata_int <= 'h2850;
    4825: romdata_int <= 'h41e; // Line Descriptor
    4826: romdata_int <= 'h200;
    4827: romdata_int <= 'h1f41;
    4828: romdata_int <= 'h258;
    4829: romdata_int <= 'h41e; // Line Descriptor
    4830: romdata_int <= 'h400;
    4831: romdata_int <= 'h1c5c;
    4832: romdata_int <= 'h2c51;
    4833: romdata_int <= 'h41e; // Line Descriptor
    4834: romdata_int <= 'h600;
    4835: romdata_int <= 'h2ab1;
    4836: romdata_int <= 'h2a43;
    4837: romdata_int <= 'h41e; // Line Descriptor
    4838: romdata_int <= 'h800;
    4839: romdata_int <= 'h1539;
    4840: romdata_int <= 'h6fa;
    4841: romdata_int <= 'h41e; // Line Descriptor
    4842: romdata_int <= 'ha00;
    4843: romdata_int <= 'h283d;
    4844: romdata_int <= 'h384d;
    4845: romdata_int <= 'h41e; // Line Descriptor
    4846: romdata_int <= 'hc00;
    4847: romdata_int <= 'h215c;
    4848: romdata_int <= 'h3145;
    4849: romdata_int <= 'h41e; // Line Descriptor
    4850: romdata_int <= 'he00;
    4851: romdata_int <= 'h1838;
    4852: romdata_int <= 'hd35;
    4853: romdata_int <= 'h41e; // Line Descriptor
    4854: romdata_int <= 'h1000;
    4855: romdata_int <= 'h234e;
    4856: romdata_int <= 'h2486;
    4857: romdata_int <= 'h41e; // Line Descriptor
    4858: romdata_int <= 'h1200;
    4859: romdata_int <= 'h884;
    4860: romdata_int <= 'h100b;
    4861: romdata_int <= 'h41e; // Line Descriptor
    4862: romdata_int <= 'h1400;
    4863: romdata_int <= 'h58;
    4864: romdata_int <= 'h22a9;
    4865: romdata_int <= 'h41e; // Line Descriptor
    4866: romdata_int <= 'h1600;
    4867: romdata_int <= 'h241c;
    4868: romdata_int <= 'h2e73;
    4869: romdata_int <= 'h41e; // Line Descriptor
    4870: romdata_int <= 'h1800;
    4871: romdata_int <= 'h4ba;
    4872: romdata_int <= 'h1abd;
    4873: romdata_int <= 'h41e; // Line Descriptor
    4874: romdata_int <= 'h1a00;
    4875: romdata_int <= 'h1b3d;
    4876: romdata_int <= 'h201e;
    4877: romdata_int <= 'h41e; // Line Descriptor
    4878: romdata_int <= 'h1c00;
    4879: romdata_int <= 'h3688;
    4880: romdata_int <= 'h3a33;
    4881: romdata_int <= 'h41e; // Line Descriptor
    4882: romdata_int <= 'h1e00;
    4883: romdata_int <= 'hc96;
    4884: romdata_int <= 'h1674;
    4885: romdata_int <= 'h41e; // Line Descriptor
    4886: romdata_int <= 'h2000;
    4887: romdata_int <= 'h311;
    4888: romdata_int <= 'h188b;
    4889: romdata_int <= 'h41e; // Line Descriptor
    4890: romdata_int <= 'h2200;
    4891: romdata_int <= 'h2d53;
    4892: romdata_int <= 'hecd;
    4893: romdata_int <= 'h41e; // Line Descriptor
    4894: romdata_int <= 'h2400;
    4895: romdata_int <= 'h38bc;
    4896: romdata_int <= 'ha6e;
    4897: romdata_int <= 'h41e; // Line Descriptor
    4898: romdata_int <= 'h2600;
    4899: romdata_int <= 'h3a72;
    4900: romdata_int <= 'h1433;
    4901: romdata_int <= 'h41e; // Line Descriptor
    4902: romdata_int <= 'h2800;
    4903: romdata_int <= 'h349e;
    4904: romdata_int <= 'h3659;
    4905: romdata_int <= 'h41e; // Line Descriptor
    4906: romdata_int <= 'h2a00;
    4907: romdata_int <= 'h2687;
    4908: romdata_int <= 'h1ede;
    4909: romdata_int <= 'h41e; // Line Descriptor
    4910: romdata_int <= 'h2c00;
    4911: romdata_int <= 'he25;
    4912: romdata_int <= 'h3421;
    4913: romdata_int <= 'h41e; // Line Descriptor
    4914: romdata_int <= 'h2e00;
    4915: romdata_int <= 'h12bb;
    4916: romdata_int <= 'h3266;
    4917: romdata_int <= 'h41e; // Line Descriptor
    4918: romdata_int <= 'h3000;
    4919: romdata_int <= 'h2f1a;
    4920: romdata_int <= 'h118;
    4921: romdata_int <= 'h41e; // Line Descriptor
    4922: romdata_int <= 'h3200;
    4923: romdata_int <= 'hb13;
    4924: romdata_int <= 'h80d;
    4925: romdata_int <= 'h41e; // Line Descriptor
    4926: romdata_int <= 'h3400;
    4927: romdata_int <= 'h10d3;
    4928: romdata_int <= 'h4a8;
    4929: romdata_int <= 'h41e; // Line Descriptor
    4930: romdata_int <= 'h3600;
    4931: romdata_int <= 'h30cd;
    4932: romdata_int <= 'h26aa;
    4933: romdata_int <= 'h41e; // Line Descriptor
    4934: romdata_int <= 'h3800;
    4935: romdata_int <= 'h6f0;
    4936: romdata_int <= 'h1242;
    4937: romdata_int <= 'h41e; // Line Descriptor
    4938: romdata_int <= 'h3a00;
    4939: romdata_int <= 'h163b;
    4940: romdata_int <= 'h1cac;
    4941: romdata_int <= 'h41e; // Line Descriptor
    4942: romdata_int <= 'h0;
    4943: romdata_int <= 'h3030;
    4944: romdata_int <= 'h2676;
    4945: romdata_int <= 'h41e; // Line Descriptor
    4946: romdata_int <= 'h200;
    4947: romdata_int <= 'h2070;
    4948: romdata_int <= 'h1c8c;
    4949: romdata_int <= 'h41e; // Line Descriptor
    4950: romdata_int <= 'h400;
    4951: romdata_int <= 'h10f1;
    4952: romdata_int <= 'he02;
    4953: romdata_int <= 'h41e; // Line Descriptor
    4954: romdata_int <= 'h600;
    4955: romdata_int <= 'hb61;
    4956: romdata_int <= 'h1726;
    4957: romdata_int <= 'h41e; // Line Descriptor
    4958: romdata_int <= 'h800;
    4959: romdata_int <= 'h2a28;
    4960: romdata_int <= 'h6d9;
    4961: romdata_int <= 'h41e; // Line Descriptor
    4962: romdata_int <= 'ha00;
    4963: romdata_int <= 'h28b0;
    4964: romdata_int <= 'h49b;
    4965: romdata_int <= 'h41e; // Line Descriptor
    4966: romdata_int <= 'hc00;
    4967: romdata_int <= 'h262f;
    4968: romdata_int <= 'h3b44;
    4969: romdata_int <= 'h41e; // Line Descriptor
    4970: romdata_int <= 'he00;
    4971: romdata_int <= 'h2506;
    4972: romdata_int <= 'h2ab;
    4973: romdata_int <= 'h41e; // Line Descriptor
    4974: romdata_int <= 'h1000;
    4975: romdata_int <= 'h3293;
    4976: romdata_int <= 'h3156;
    4977: romdata_int <= 'h41e; // Line Descriptor
    4978: romdata_int <= 'h1200;
    4979: romdata_int <= 'h2d3;
    4980: romdata_int <= 'h22b7;
    4981: romdata_int <= 'h41e; // Line Descriptor
    4982: romdata_int <= 'h1400;
    4983: romdata_int <= 'h4de;
    4984: romdata_int <= 'h2aa4;
    4985: romdata_int <= 'h41e; // Line Descriptor
    4986: romdata_int <= 'h1600;
    4987: romdata_int <= 'h1d40;
    4988: romdata_int <= 'h1155;
    4989: romdata_int <= 'h41e; // Line Descriptor
    4990: romdata_int <= 'h1800;
    4991: romdata_int <= 'h118;
    4992: romdata_int <= 'h1f0b;
    4993: romdata_int <= 'h41e; // Line Descriptor
    4994: romdata_int <= 'h1a00;
    4995: romdata_int <= 'hd31;
    4996: romdata_int <= 'h28bb;
    4997: romdata_int <= 'h41e; // Line Descriptor
    4998: romdata_int <= 'h1c00;
    4999: romdata_int <= 'h22eb;
    5000: romdata_int <= 'h3927;
    5001: romdata_int <= 'h41e; // Line Descriptor
    5002: romdata_int <= 'h1e00;
    5003: romdata_int <= 'h372c;
    5004: romdata_int <= 'h3271;
    5005: romdata_int <= 'h41e; // Line Descriptor
    5006: romdata_int <= 'h2000;
    5007: romdata_int <= 'h1438;
    5008: romdata_int <= 'h3480;
    5009: romdata_int <= 'h41e; // Line Descriptor
    5010: romdata_int <= 'h2200;
    5011: romdata_int <= 'h85f;
    5012: romdata_int <= 'h131a;
    5013: romdata_int <= 'h41e; // Line Descriptor
    5014: romdata_int <= 'h2400;
    5015: romdata_int <= 'h34ce;
    5016: romdata_int <= 'h15;
    5017: romdata_int <= 'h41e; // Line Descriptor
    5018: romdata_int <= 'h2600;
    5019: romdata_int <= 'h60c;
    5020: romdata_int <= 'h2eb5;
    5021: romdata_int <= 'h41e; // Line Descriptor
    5022: romdata_int <= 'h2800;
    5023: romdata_int <= 'h1e89;
    5024: romdata_int <= 'h24e9;
    5025: romdata_int <= 'h41e; // Line Descriptor
    5026: romdata_int <= 'h2a00;
    5027: romdata_int <= 'h2c35;
    5028: romdata_int <= 'h18df;
    5029: romdata_int <= 'h41e; // Line Descriptor
    5030: romdata_int <= 'h2c00;
    5031: romdata_int <= 'h132e;
    5032: romdata_int <= 'h2133;
    5033: romdata_int <= 'h41e; // Line Descriptor
    5034: romdata_int <= 'h2e00;
    5035: romdata_int <= 'hec0;
    5036: romdata_int <= 'h1487;
    5037: romdata_int <= 'h41e; // Line Descriptor
    5038: romdata_int <= 'h3000;
    5039: romdata_int <= 'h2e7c;
    5040: romdata_int <= 'h3733;
    5041: romdata_int <= 'h41e; // Line Descriptor
    5042: romdata_int <= 'h3200;
    5043: romdata_int <= 'h38e9;
    5044: romdata_int <= 'h2cb9;
    5045: romdata_int <= 'h41e; // Line Descriptor
    5046: romdata_int <= 'h3400;
    5047: romdata_int <= 'h1928;
    5048: romdata_int <= 'hc97;
    5049: romdata_int <= 'h41e; // Line Descriptor
    5050: romdata_int <= 'h3600;
    5051: romdata_int <= 'h1a1c;
    5052: romdata_int <= 'h8ca;
    5053: romdata_int <= 'h41e; // Line Descriptor
    5054: romdata_int <= 'h3800;
    5055: romdata_int <= 'h3b0c;
    5056: romdata_int <= 'h1ac4;
    5057: romdata_int <= 'h41e; // Line Descriptor
    5058: romdata_int <= 'h3a00;
    5059: romdata_int <= 'h1644;
    5060: romdata_int <= 'ha60;
    5061: romdata_int <= 'h41e; // Line Descriptor
    5062: romdata_int <= 'h0;
    5063: romdata_int <= 'h1764;
    5064: romdata_int <= 'h669;
    5065: romdata_int <= 'h41e; // Line Descriptor
    5066: romdata_int <= 'h200;
    5067: romdata_int <= 'h478;
    5068: romdata_int <= 'ha87;
    5069: romdata_int <= 'h41e; // Line Descriptor
    5070: romdata_int <= 'h400;
    5071: romdata_int <= 'h380a;
    5072: romdata_int <= 'he39;
    5073: romdata_int <= 'h41e; // Line Descriptor
    5074: romdata_int <= 'h600;
    5075: romdata_int <= 'h3a49;
    5076: romdata_int <= 'h3b35;
    5077: romdata_int <= 'h41e; // Line Descriptor
    5078: romdata_int <= 'h800;
    5079: romdata_int <= 'h2640;
    5080: romdata_int <= 'h1107;
    5081: romdata_int <= 'h41e; // Line Descriptor
    5082: romdata_int <= 'ha00;
    5083: romdata_int <= 'h2214;
    5084: romdata_int <= 'h3406;
    5085: romdata_int <= 'h41e; // Line Descriptor
    5086: romdata_int <= 'hc00;
    5087: romdata_int <= 'h311c;
    5088: romdata_int <= 'h302d;
    5089: romdata_int <= 'h41e; // Line Descriptor
    5090: romdata_int <= 'he00;
    5091: romdata_int <= 'h3563;
    5092: romdata_int <= 'h6c;
    5093: romdata_int <= 'h41e; // Line Descriptor
    5094: romdata_int <= 'h1000;
    5095: romdata_int <= 'h18de;
    5096: romdata_int <= 'h133c;
    5097: romdata_int <= 'h41e; // Line Descriptor
    5098: romdata_int <= 'h1200;
    5099: romdata_int <= 'h2869;
    5100: romdata_int <= 'h22f8;
    5101: romdata_int <= 'h41e; // Line Descriptor
    5102: romdata_int <= 'h1400;
    5103: romdata_int <= 'h1106;
    5104: romdata_int <= 'h2bf;
    5105: romdata_int <= 'h41e; // Line Descriptor
    5106: romdata_int <= 'h1600;
    5107: romdata_int <= 'h2cc;
    5108: romdata_int <= 'h2d65;
    5109: romdata_int <= 'h41e; // Line Descriptor
    5110: romdata_int <= 'h1800;
    5111: romdata_int <= 'h1aa1;
    5112: romdata_int <= 'h1930;
    5113: romdata_int <= 'h41e; // Line Descriptor
    5114: romdata_int <= 'h1a00;
    5115: romdata_int <= 'h1413;
    5116: romdata_int <= 'h2b3f;
    5117: romdata_int <= 'h41e; // Line Descriptor
    5118: romdata_int <= 'h1c00;
    5119: romdata_int <= 'h36d0;
    5120: romdata_int <= 'h2935;
    5121: romdata_int <= 'h41e; // Line Descriptor
    5122: romdata_int <= 'h1e00;
    5123: romdata_int <= 'h1264;
    5124: romdata_int <= 'h244b;
    5125: romdata_int <= 'h41e; // Line Descriptor
    5126: romdata_int <= 'h2000;
    5127: romdata_int <= 'h1e06;
    5128: romdata_int <= 'h2650;
    5129: romdata_int <= 'h41e; // Line Descriptor
    5130: romdata_int <= 'h2200;
    5131: romdata_int <= 'hd0b;
    5132: romdata_int <= 'h3633;
    5133: romdata_int <= 'h41e; // Line Descriptor
    5134: romdata_int <= 'h2400;
    5135: romdata_int <= 'h2032;
    5136: romdata_int <= 'h1f32;
    5137: romdata_int <= 'h41e; // Line Descriptor
    5138: romdata_int <= 'h2600;
    5139: romdata_int <= 'h2d0c;
    5140: romdata_int <= 'h92e;
    5141: romdata_int <= 'h41e; // Line Descriptor
    5142: romdata_int <= 'h2800;
    5143: romdata_int <= 'h3245;
    5144: romdata_int <= 'h392a;
    5145: romdata_int <= 'h41e; // Line Descriptor
    5146: romdata_int <= 'h2a00;
    5147: romdata_int <= 'h619;
    5148: romdata_int <= 'hcf4;
    5149: romdata_int <= 'h41e; // Line Descriptor
    5150: romdata_int <= 'h2c00;
    5151: romdata_int <= 'h2ad1;
    5152: romdata_int <= 'h2e7f;
    5153: romdata_int <= 'h41e; // Line Descriptor
    5154: romdata_int <= 'h2e00;
    5155: romdata_int <= 'h857;
    5156: romdata_int <= 'h1d05;
    5157: romdata_int <= 'h41e; // Line Descriptor
    5158: romdata_int <= 'h3000;
    5159: romdata_int <= 'h2e4c;
    5160: romdata_int <= 'h2015;
    5161: romdata_int <= 'h41e; // Line Descriptor
    5162: romdata_int <= 'h3200;
    5163: romdata_int <= 'ha45;
    5164: romdata_int <= 'h1614;
    5165: romdata_int <= 'h41e; // Line Descriptor
    5166: romdata_int <= 'h3400;
    5167: romdata_int <= 'he9c;
    5168: romdata_int <= 'h40c;
    5169: romdata_int <= 'h41e; // Line Descriptor
    5170: romdata_int <= 'h3600;
    5171: romdata_int <= 'h1d21;
    5172: romdata_int <= 'h154b;
    5173: romdata_int <= 'h41e; // Line Descriptor
    5174: romdata_int <= 'h3800;
    5175: romdata_int <= 'ha1;
    5176: romdata_int <= 'h3244;
    5177: romdata_int <= 'h41e; // Line Descriptor
    5178: romdata_int <= 'h3a00;
    5179: romdata_int <= 'h24ea;
    5180: romdata_int <= 'h1a2d;
    5181: romdata_int <= 'h41e; // Line Descriptor
    5182: romdata_int <= 'h0;
    5183: romdata_int <= 'h3a3a;
    5184: romdata_int <= 'hf05;
    5185: romdata_int <= 'h41e; // Line Descriptor
    5186: romdata_int <= 'h200;
    5187: romdata_int <= 'h2a7e;
    5188: romdata_int <= 'h1238;
    5189: romdata_int <= 'h41e; // Line Descriptor
    5190: romdata_int <= 'h400;
    5191: romdata_int <= 'h294f;
    5192: romdata_int <= 'h264e;
    5193: romdata_int <= 'h41e; // Line Descriptor
    5194: romdata_int <= 'h600;
    5195: romdata_int <= 'he7a;
    5196: romdata_int <= 'h254a;
    5197: romdata_int <= 'h41e; // Line Descriptor
    5198: romdata_int <= 'h800;
    5199: romdata_int <= 'h303f;
    5200: romdata_int <= 'h28e6;
    5201: romdata_int <= 'h41e; // Line Descriptor
    5202: romdata_int <= 'ha00;
    5203: romdata_int <= 'h1c8d;
    5204: romdata_int <= 'h3abc;
    5205: romdata_int <= 'h41e; // Line Descriptor
    5206: romdata_int <= 'hc00;
    5207: romdata_int <= 'h1f55;
    5208: romdata_int <= 'h2b04;
    5209: romdata_int <= 'h41e; // Line Descriptor
    5210: romdata_int <= 'he00;
    5211: romdata_int <= 'h38fe;
    5212: romdata_int <= 'h1c83;
    5213: romdata_int <= 'h41e; // Line Descriptor
    5214: romdata_int <= 'h1000;
    5215: romdata_int <= 'h146e;
    5216: romdata_int <= 'h38b6;
    5217: romdata_int <= 'h41e; // Line Descriptor
    5218: romdata_int <= 'h1200;
    5219: romdata_int <= 'h20d3;
    5220: romdata_int <= 'hd42;
    5221: romdata_int <= 'h41e; // Line Descriptor
    5222: romdata_int <= 'h1400;
    5223: romdata_int <= 'h10ec;
    5224: romdata_int <= 'h4cc;
    5225: romdata_int <= 'h41e; // Line Descriptor
    5226: romdata_int <= 'h1600;
    5227: romdata_int <= 'h22b;
    5228: romdata_int <= 'h3704;
    5229: romdata_int <= 'h41e; // Line Descriptor
    5230: romdata_int <= 'h1800;
    5231: romdata_int <= 'h561;
    5232: romdata_int <= 'hb2a;
    5233: romdata_int <= 'h41e; // Line Descriptor
    5234: romdata_int <= 'h1a00;
    5235: romdata_int <= 'h1278;
    5236: romdata_int <= 'h14ed;
    5237: romdata_int <= 'h41e; // Line Descriptor
    5238: romdata_int <= 'h1c00;
    5239: romdata_int <= 'h2531;
    5240: romdata_int <= 'h2d2f;
    5241: romdata_int <= 'h41e; // Line Descriptor
    5242: romdata_int <= 'h1e00;
    5243: romdata_int <= 'h2ece;
    5244: romdata_int <= 'h190c;
    5245: romdata_int <= 'h41e; // Line Descriptor
    5246: romdata_int <= 'h2000;
    5247: romdata_int <= 'h6f;
    5248: romdata_int <= 'h1e60;
    5249: romdata_int <= 'h41e; // Line Descriptor
    5250: romdata_int <= 'h2200;
    5251: romdata_int <= 'h88e;
    5252: romdata_int <= 'h760;
    5253: romdata_int <= 'h41e; // Line Descriptor
    5254: romdata_int <= 'h2400;
    5255: romdata_int <= 'h355f;
    5256: romdata_int <= 'h20d8;
    5257: romdata_int <= 'h41e; // Line Descriptor
    5258: romdata_int <= 'h2600;
    5259: romdata_int <= 'h2325;
    5260: romdata_int <= 'h32fe;
    5261: romdata_int <= 'h41e; // Line Descriptor
    5262: romdata_int <= 'h2800;
    5263: romdata_int <= 'h2642;
    5264: romdata_int <= 'h97;
    5265: romdata_int <= 'h41e; // Line Descriptor
    5266: romdata_int <= 'h2a00;
    5267: romdata_int <= 'h2d32;
    5268: romdata_int <= 'h10e3;
    5269: romdata_int <= 'h41e; // Line Descriptor
    5270: romdata_int <= 'h2c00;
    5271: romdata_int <= 'h1a71;
    5272: romdata_int <= 'h3039;
    5273: romdata_int <= 'h41e; // Line Descriptor
    5274: romdata_int <= 'h2e00;
    5275: romdata_int <= 'hc46;
    5276: romdata_int <= 'h2f2c;
    5277: romdata_int <= 'h41e; // Line Descriptor
    5278: romdata_int <= 'h3000;
    5279: romdata_int <= 'h16e5;
    5280: romdata_int <= 'h1a81;
    5281: romdata_int <= 'h41e; // Line Descriptor
    5282: romdata_int <= 'h3200;
    5283: romdata_int <= 'h3281;
    5284: romdata_int <= 'h1648;
    5285: romdata_int <= 'h41e; // Line Descriptor
    5286: romdata_int <= 'h3400;
    5287: romdata_int <= 'h1887;
    5288: romdata_int <= 'h8d6;
    5289: romdata_int <= 'h41e; // Line Descriptor
    5290: romdata_int <= 'h3600;
    5291: romdata_int <= 'ha7d;
    5292: romdata_int <= 'h353d;
    5293: romdata_int <= 'h41e; // Line Descriptor
    5294: romdata_int <= 'h3800;
    5295: romdata_int <= 'h69c;
    5296: romdata_int <= 'h247;
    5297: romdata_int <= 'h51e; // Line Descriptor
    5298: romdata_int <= 'h3a00;
    5299: romdata_int <= 'h36f4;
    5300: romdata_int <= 'h230b;
    5301: romdata_int <= 'h614; // Line Descriptor
    5302: romdata_int <= 'h0;
    5303: romdata_int <= 'h1f37;
    5304: romdata_int <= 'h108e;
    5305: romdata_int <= 'h4a1;
    5306: romdata_int <= 'h614; // Line Descriptor
    5307: romdata_int <= 'h200;
    5308: romdata_int <= 'h122;
    5309: romdata_int <= 'h18ae;
    5310: romdata_int <= 'h110b;
    5311: romdata_int <= 'h614; // Line Descriptor
    5312: romdata_int <= 'h400;
    5313: romdata_int <= 'h2289;
    5314: romdata_int <= 'he2e;
    5315: romdata_int <= 'h1404;
    5316: romdata_int <= 'h614; // Line Descriptor
    5317: romdata_int <= 'h600;
    5318: romdata_int <= 'h35c;
    5319: romdata_int <= 'h20e1;
    5320: romdata_int <= 'h26ec;
    5321: romdata_int <= 'h614; // Line Descriptor
    5322: romdata_int <= 'h800;
    5323: romdata_int <= 'h183a;
    5324: romdata_int <= 'h22a1;
    5325: romdata_int <= 'h939;
    5326: romdata_int <= 'h614; // Line Descriptor
    5327: romdata_int <= 'ha00;
    5328: romdata_int <= 'he60;
    5329: romdata_int <= 'ha79;
    5330: romdata_int <= 'h6b8;
    5331: romdata_int <= 'h614; // Line Descriptor
    5332: romdata_int <= 'hc00;
    5333: romdata_int <= 'h1cb9;
    5334: romdata_int <= 'h133b;
    5335: romdata_int <= 'h1e7c;
    5336: romdata_int <= 'h614; // Line Descriptor
    5337: romdata_int <= 'he00;
    5338: romdata_int <= 'h1499;
    5339: romdata_int <= 'h53d;
    5340: romdata_int <= 'h1d65;
    5341: romdata_int <= 'h614; // Line Descriptor
    5342: romdata_int <= 'h1000;
    5343: romdata_int <= 'h1079;
    5344: romdata_int <= 'h1a1e;
    5345: romdata_int <= 'h2bc;
    5346: romdata_int <= 'h614; // Line Descriptor
    5347: romdata_int <= 'h1200;
    5348: romdata_int <= 'hc91;
    5349: romdata_int <= 'h80d;
    5350: romdata_int <= 'hf28;
    5351: romdata_int <= 'h614; // Line Descriptor
    5352: romdata_int <= 'h1400;
    5353: romdata_int <= 'h2055;
    5354: romdata_int <= 'h1461;
    5355: romdata_int <= 'h1ad5;
    5356: romdata_int <= 'h614; // Line Descriptor
    5357: romdata_int <= 'h1600;
    5358: romdata_int <= 'h1ae6;
    5359: romdata_int <= 'h2734;
    5360: romdata_int <= 'h16ae;
    5361: romdata_int <= 'h614; // Line Descriptor
    5362: romdata_int <= 'h1800;
    5363: romdata_int <= 'haf3;
    5364: romdata_int <= 'hca4;
    5365: romdata_int <= 'hb2c;
    5366: romdata_int <= 'h614; // Line Descriptor
    5367: romdata_int <= 'h1a00;
    5368: romdata_int <= 'h643;
    5369: romdata_int <= 'h728;
    5370: romdata_int <= 'h12b0;
    5371: romdata_int <= 'h614; // Line Descriptor
    5372: romdata_int <= 'h1c00;
    5373: romdata_int <= 'h12e5;
    5374: romdata_int <= 'h1ec9;
    5375: romdata_int <= 'h186a;
    5376: romdata_int <= 'h614; // Line Descriptor
    5377: romdata_int <= 'h1e00;
    5378: romdata_int <= 'h264e;
    5379: romdata_int <= 'hc4;
    5380: romdata_int <= 'h2350;
    5381: romdata_int <= 'h614; // Line Descriptor
    5382: romdata_int <= 'h2000;
    5383: romdata_int <= 'h852;
    5384: romdata_int <= 'h163b;
    5385: romdata_int <= 'h252b;
    5386: romdata_int <= 'h614; // Line Descriptor
    5387: romdata_int <= 'h2200;
    5388: romdata_int <= 'h44a;
    5389: romdata_int <= 'h277;
    5390: romdata_int <= 'he7;
    5391: romdata_int <= 'h614; // Line Descriptor
    5392: romdata_int <= 'h2400;
    5393: romdata_int <= 'h1753;
    5394: romdata_int <= 'h1d2c;
    5395: romdata_int <= 'h2149;
    5396: romdata_int <= 'h614; // Line Descriptor
    5397: romdata_int <= 'h2600;
    5398: romdata_int <= 'h2488;
    5399: romdata_int <= 'h2527;
    5400: romdata_int <= 'hcbd;
    5401: romdata_int <= 'h414; // Line Descriptor
    5402: romdata_int <= 'h0;
    5403: romdata_int <= 'h2101;
    5404: romdata_int <= 'hd34;
    5405: romdata_int <= 'h414; // Line Descriptor
    5406: romdata_int <= 'h200;
    5407: romdata_int <= 'h84b;
    5408: romdata_int <= 'h20d9;
    5409: romdata_int <= 'h414; // Line Descriptor
    5410: romdata_int <= 'h400;
    5411: romdata_int <= 'h1406;
    5412: romdata_int <= 'h85f;
    5413: romdata_int <= 'h414; // Line Descriptor
    5414: romdata_int <= 'h600;
    5415: romdata_int <= 'hf2d;
    5416: romdata_int <= 'he9f;
    5417: romdata_int <= 'h414; // Line Descriptor
    5418: romdata_int <= 'h800;
    5419: romdata_int <= 'h254f;
    5420: romdata_int <= 'h2625;
    5421: romdata_int <= 'h414; // Line Descriptor
    5422: romdata_int <= 'ha00;
    5423: romdata_int <= 'h138;
    5424: romdata_int <= 'h148f;
    5425: romdata_int <= 'h414; // Line Descriptor
    5426: romdata_int <= 'hc00;
    5427: romdata_int <= 'h675;
    5428: romdata_int <= 'h1641;
    5429: romdata_int <= 'h414; // Line Descriptor
    5430: romdata_int <= 'he00;
    5431: romdata_int <= 'h2633;
    5432: romdata_int <= 'hb11;
    5433: romdata_int <= 'h414; // Line Descriptor
    5434: romdata_int <= 'h1000;
    5435: romdata_int <= 'h234a;
    5436: romdata_int <= 'h1a7d;
    5437: romdata_int <= 'h414; // Line Descriptor
    5438: romdata_int <= 'h1200;
    5439: romdata_int <= 'h104f;
    5440: romdata_int <= 'h505;
    5441: romdata_int <= 'h414; // Line Descriptor
    5442: romdata_int <= 'h1400;
    5443: romdata_int <= 'h348;
    5444: romdata_int <= 'h1e1a;
    5445: romdata_int <= 'h414; // Line Descriptor
    5446: romdata_int <= 'h1600;
    5447: romdata_int <= 'haee;
    5448: romdata_int <= 'h1c66;
    5449: romdata_int <= 'h414; // Line Descriptor
    5450: romdata_int <= 'h1800;
    5451: romdata_int <= 'hd2a;
    5452: romdata_int <= 'h1958;
    5453: romdata_int <= 'h414; // Line Descriptor
    5454: romdata_int <= 'h1a00;
    5455: romdata_int <= 'h1262;
    5456: romdata_int <= 'h12c1;
    5457: romdata_int <= 'h414; // Line Descriptor
    5458: romdata_int <= 'h1c00;
    5459: romdata_int <= 'h16b2;
    5460: romdata_int <= 'h79;
    5461: romdata_int <= 'h414; // Line Descriptor
    5462: romdata_int <= 'h1e00;
    5463: romdata_int <= 'h18e7;
    5464: romdata_int <= 'h231;
    5465: romdata_int <= 'h414; // Line Descriptor
    5466: romdata_int <= 'h2000;
    5467: romdata_int <= 'h1ea0;
    5468: romdata_int <= 'h6d0;
    5469: romdata_int <= 'h414; // Line Descriptor
    5470: romdata_int <= 'h2200;
    5471: romdata_int <= 'h1a30;
    5472: romdata_int <= 'h229b;
    5473: romdata_int <= 'h414; // Line Descriptor
    5474: romdata_int <= 'h2400;
    5475: romdata_int <= 'h4be;
    5476: romdata_int <= 'h2535;
    5477: romdata_int <= 'h414; // Line Descriptor
    5478: romdata_int <= 'h2600;
    5479: romdata_int <= 'h1cbd;
    5480: romdata_int <= 'h10c5;
    5481: romdata_int <= 'h414; // Line Descriptor
    5482: romdata_int <= 'h0;
    5483: romdata_int <= 'h209f;
    5484: romdata_int <= 'hd32;
    5485: romdata_int <= 'h414; // Line Descriptor
    5486: romdata_int <= 'h200;
    5487: romdata_int <= 'h1a1c;
    5488: romdata_int <= 'h125f;
    5489: romdata_int <= 'h414; // Line Descriptor
    5490: romdata_int <= 'h400;
    5491: romdata_int <= 'h142a;
    5492: romdata_int <= 'h1cc9;
    5493: romdata_int <= 'h414; // Line Descriptor
    5494: romdata_int <= 'h600;
    5495: romdata_int <= 'h519;
    5496: romdata_int <= 'h250;
    5497: romdata_int <= 'h414; // Line Descriptor
    5498: romdata_int <= 'h800;
    5499: romdata_int <= 'hb2c;
    5500: romdata_int <= 'h81a;
    5501: romdata_int <= 'h414; // Line Descriptor
    5502: romdata_int <= 'ha00;
    5503: romdata_int <= 'h1706;
    5504: romdata_int <= 'h721;
    5505: romdata_int <= 'h414; // Line Descriptor
    5506: romdata_int <= 'hc00;
    5507: romdata_int <= 'h1808;
    5508: romdata_int <= 'h1865;
    5509: romdata_int <= 'h414; // Line Descriptor
    5510: romdata_int <= 'he00;
    5511: romdata_int <= 'h1e5d;
    5512: romdata_int <= 'h1e7b;
    5513: romdata_int <= 'h414; // Line Descriptor
    5514: romdata_int <= 'h1000;
    5515: romdata_int <= 'h2218;
    5516: romdata_int <= 'h1640;
    5517: romdata_int <= 'h414; // Line Descriptor
    5518: romdata_int <= 'h1200;
    5519: romdata_int <= 'hc80;
    5520: romdata_int <= 'h14ab;
    5521: romdata_int <= 'h414; // Line Descriptor
    5522: romdata_int <= 'h1400;
    5523: romdata_int <= 'h123e;
    5524: romdata_int <= 'h25;
    5525: romdata_int <= 'h414; // Line Descriptor
    5526: romdata_int <= 'h1600;
    5527: romdata_int <= 'h893;
    5528: romdata_int <= 'h1061;
    5529: romdata_int <= 'h414; // Line Descriptor
    5530: romdata_int <= 'h1800;
    5531: romdata_int <= 'h1146;
    5532: romdata_int <= 'h2690;
    5533: romdata_int <= 'h414; // Line Descriptor
    5534: romdata_int <= 'h1a00;
    5535: romdata_int <= 'h670;
    5536: romdata_int <= 'h20b4;
    5537: romdata_int <= 'h414; // Line Descriptor
    5538: romdata_int <= 'h1c00;
    5539: romdata_int <= 'he2b;
    5540: romdata_int <= 'h1aba;
    5541: romdata_int <= 'h414; // Line Descriptor
    5542: romdata_int <= 'h1e00;
    5543: romdata_int <= 'h1c44;
    5544: romdata_int <= 'h4eb;
    5545: romdata_int <= 'h414; // Line Descriptor
    5546: romdata_int <= 'h2000;
    5547: romdata_int <= 'h24ea;
    5548: romdata_int <= 'ha72;
    5549: romdata_int <= 'h414; // Line Descriptor
    5550: romdata_int <= 'h2200;
    5551: romdata_int <= 'hee;
    5552: romdata_int <= 'h22c3;
    5553: romdata_int <= 'h414; // Line Descriptor
    5554: romdata_int <= 'h2400;
    5555: romdata_int <= 'h265c;
    5556: romdata_int <= 'h24ca;
    5557: romdata_int <= 'h414; // Line Descriptor
    5558: romdata_int <= 'h2600;
    5559: romdata_int <= 'h333;
    5560: romdata_int <= 'heb0;
    5561: romdata_int <= 'h414; // Line Descriptor
    5562: romdata_int <= 'h0;
    5563: romdata_int <= 'h106b;
    5564: romdata_int <= 'hcfd;
    5565: romdata_int <= 'h414; // Line Descriptor
    5566: romdata_int <= 'h200;
    5567: romdata_int <= 'hc41;
    5568: romdata_int <= 'ha07;
    5569: romdata_int <= 'h414; // Line Descriptor
    5570: romdata_int <= 'h400;
    5571: romdata_int <= 'h2673;
    5572: romdata_int <= 'h162b;
    5573: romdata_int <= 'h414; // Line Descriptor
    5574: romdata_int <= 'h600;
    5575: romdata_int <= 'h6ad;
    5576: romdata_int <= 'h235;
    5577: romdata_int <= 'h414; // Line Descriptor
    5578: romdata_int <= 'h800;
    5579: romdata_int <= 'h1d15;
    5580: romdata_int <= 'hf4c;
    5581: romdata_int <= 'h414; // Line Descriptor
    5582: romdata_int <= 'ha00;
    5583: romdata_int <= 'h2323;
    5584: romdata_int <= 'h2610;
    5585: romdata_int <= 'h414; // Line Descriptor
    5586: romdata_int <= 'hc00;
    5587: romdata_int <= 'h323;
    5588: romdata_int <= 'h18f6;
    5589: romdata_int <= 'h414; // Line Descriptor
    5590: romdata_int <= 'he00;
    5591: romdata_int <= 'h213d;
    5592: romdata_int <= 'h20ed;
    5593: romdata_int <= 'h414; // Line Descriptor
    5594: romdata_int <= 'h1000;
    5595: romdata_int <= 'h14c4;
    5596: romdata_int <= 'h2414;
    5597: romdata_int <= 'h414; // Line Descriptor
    5598: romdata_int <= 'h1200;
    5599: romdata_int <= 'h160a;
    5600: romdata_int <= 'h1c9a;
    5601: romdata_int <= 'h414; // Line Descriptor
    5602: romdata_int <= 'h1400;
    5603: romdata_int <= 'he32;
    5604: romdata_int <= 'h10f6;
    5605: romdata_int <= 'h414; // Line Descriptor
    5606: romdata_int <= 'h1600;
    5607: romdata_int <= 'h8b3;
    5608: romdata_int <= 'h1e3d;
    5609: romdata_int <= 'h414; // Line Descriptor
    5610: romdata_int <= 'h1800;
    5611: romdata_int <= 'h55d;
    5612: romdata_int <= 'h128f;
    5613: romdata_int <= 'h414; // Line Descriptor
    5614: romdata_int <= 'h1a00;
    5615: romdata_int <= 'h1850;
    5616: romdata_int <= 'h1a32;
    5617: romdata_int <= 'h414; // Line Descriptor
    5618: romdata_int <= 'h1c00;
    5619: romdata_int <= 'h1a2f;
    5620: romdata_int <= 'h8f8;
    5621: romdata_int <= 'h414; // Line Descriptor
    5622: romdata_int <= 'h1e00;
    5623: romdata_int <= 'h1ee3;
    5624: romdata_int <= 'h14dc;
    5625: romdata_int <= 'h414; // Line Descriptor
    5626: romdata_int <= 'h2000;
    5627: romdata_int <= 'haf6;
    5628: romdata_int <= 'h4f2;
    5629: romdata_int <= 'h414; // Line Descriptor
    5630: romdata_int <= 'h2200;
    5631: romdata_int <= 'h2520;
    5632: romdata_int <= 'h1e;
    5633: romdata_int <= 'h414; // Line Descriptor
    5634: romdata_int <= 'h2400;
    5635: romdata_int <= 'h1345;
    5636: romdata_int <= 'h2278;
    5637: romdata_int <= 'h414; // Line Descriptor
    5638: romdata_int <= 'h2600;
    5639: romdata_int <= 'h3f;
    5640: romdata_int <= 'h6f5;
    5641: romdata_int <= 'h414; // Line Descriptor
    5642: romdata_int <= 'h0;
    5643: romdata_int <= 'h12a8;
    5644: romdata_int <= 'h1697;
    5645: romdata_int <= 'h414; // Line Descriptor
    5646: romdata_int <= 'h200;
    5647: romdata_int <= 'h22b1;
    5648: romdata_int <= 'h8a1;
    5649: romdata_int <= 'h414; // Line Descriptor
    5650: romdata_int <= 'h400;
    5651: romdata_int <= 'h1097;
    5652: romdata_int <= 'h61d;
    5653: romdata_int <= 'h414; // Line Descriptor
    5654: romdata_int <= 'h600;
    5655: romdata_int <= 'h24a2;
    5656: romdata_int <= 'h16;
    5657: romdata_int <= 'h414; // Line Descriptor
    5658: romdata_int <= 'h800;
    5659: romdata_int <= 'hd37;
    5660: romdata_int <= 'h1f4c;
    5661: romdata_int <= 'h414; // Line Descriptor
    5662: romdata_int <= 'ha00;
    5663: romdata_int <= 'h1ef4;
    5664: romdata_int <= 'h1c36;
    5665: romdata_int <= 'h414; // Line Descriptor
    5666: romdata_int <= 'hc00;
    5667: romdata_int <= 'h24a;
    5668: romdata_int <= 'hf56;
    5669: romdata_int <= 'h414; // Line Descriptor
    5670: romdata_int <= 'he00;
    5671: romdata_int <= 'h1add;
    5672: romdata_int <= 'h1860;
    5673: romdata_int <= 'h414; // Line Descriptor
    5674: romdata_int <= 'h1000;
    5675: romdata_int <= 'he69;
    5676: romdata_int <= 'h1252;
    5677: romdata_int <= 'h414; // Line Descriptor
    5678: romdata_int <= 'h1200;
    5679: romdata_int <= 'h2669;
    5680: romdata_int <= 'ha67;
    5681: romdata_int <= 'h414; // Line Descriptor
    5682: romdata_int <= 'h1400;
    5683: romdata_int <= 'h6c8;
    5684: romdata_int <= 'h113f;
    5685: romdata_int <= 'h414; // Line Descriptor
    5686: romdata_int <= 'h1600;
    5687: romdata_int <= 'h150;
    5688: romdata_int <= 'h4b5;
    5689: romdata_int <= 'h414; // Line Descriptor
    5690: romdata_int <= 'h1800;
    5691: romdata_int <= 'h1cb8;
    5692: romdata_int <= 'h2e2;
    5693: romdata_int <= 'h414; // Line Descriptor
    5694: romdata_int <= 'h1a00;
    5695: romdata_int <= 'h83a;
    5696: romdata_int <= 'h1560;
    5697: romdata_int <= 'h414; // Line Descriptor
    5698: romdata_int <= 'h1c00;
    5699: romdata_int <= 'ha62;
    5700: romdata_int <= 'h1ab4;
    5701: romdata_int <= 'h414; // Line Descriptor
    5702: romdata_int <= 'h1e00;
    5703: romdata_int <= 'h16d8;
    5704: romdata_int <= 'hc03;
    5705: romdata_int <= 'h414; // Line Descriptor
    5706: romdata_int <= 'h2000;
    5707: romdata_int <= 'h1494;
    5708: romdata_int <= 'h2059;
    5709: romdata_int <= 'h414; // Line Descriptor
    5710: romdata_int <= 'h2200;
    5711: romdata_int <= 'h18e8;
    5712: romdata_int <= 'h24a0;
    5713: romdata_int <= 'h414; // Line Descriptor
    5714: romdata_int <= 'h2400;
    5715: romdata_int <= 'h458;
    5716: romdata_int <= 'h22ee;
    5717: romdata_int <= 'h414; // Line Descriptor
    5718: romdata_int <= 'h2600;
    5719: romdata_int <= 'h211e;
    5720: romdata_int <= 'h2645;
    5721: romdata_int <= 'h414; // Line Descriptor
    5722: romdata_int <= 'h0;
    5723: romdata_int <= 'h1430;
    5724: romdata_int <= 'h1880;
    5725: romdata_int <= 'h414; // Line Descriptor
    5726: romdata_int <= 'h200;
    5727: romdata_int <= 'h467;
    5728: romdata_int <= 'h2749;
    5729: romdata_int <= 'h414; // Line Descriptor
    5730: romdata_int <= 'h400;
    5731: romdata_int <= 'h22e5;
    5732: romdata_int <= 'h14f3;
    5733: romdata_int <= 'h414; // Line Descriptor
    5734: romdata_int <= 'h600;
    5735: romdata_int <= 'h103d;
    5736: romdata_int <= 'h1b59;
    5737: romdata_int <= 'h414; // Line Descriptor
    5738: romdata_int <= 'h800;
    5739: romdata_int <= 'h26cf;
    5740: romdata_int <= 'h2233;
    5741: romdata_int <= 'h414; // Line Descriptor
    5742: romdata_int <= 'ha00;
    5743: romdata_int <= 'h2091;
    5744: romdata_int <= 'h476;
    5745: romdata_int <= 'h414; // Line Descriptor
    5746: romdata_int <= 'hc00;
    5747: romdata_int <= 'h1e13;
    5748: romdata_int <= 'hc3d;
    5749: romdata_int <= 'h414; // Line Descriptor
    5750: romdata_int <= 'he00;
    5751: romdata_int <= 'h1759;
    5752: romdata_int <= 'h10e3;
    5753: romdata_int <= 'h414; // Line Descriptor
    5754: romdata_int <= 'h1000;
    5755: romdata_int <= 'h24e6;
    5756: romdata_int <= 'h270;
    5757: romdata_int <= 'h414; // Line Descriptor
    5758: romdata_int <= 'h1200;
    5759: romdata_int <= 'hce;
    5760: romdata_int <= 'hd6;
    5761: romdata_int <= 'h414; // Line Descriptor
    5762: romdata_int <= 'h1400;
    5763: romdata_int <= 'hb23;
    5764: romdata_int <= 'h1c17;
    5765: romdata_int <= 'h414; // Line Descriptor
    5766: romdata_int <= 'h1600;
    5767: romdata_int <= 'h1c6b;
    5768: romdata_int <= 'h2515;
    5769: romdata_int <= 'h414; // Line Descriptor
    5770: romdata_int <= 'h1800;
    5771: romdata_int <= 'h1abd;
    5772: romdata_int <= 'h1711;
    5773: romdata_int <= 'h414; // Line Descriptor
    5774: romdata_int <= 'h1a00;
    5775: romdata_int <= 'hf1d;
    5776: romdata_int <= 'h1e4f;
    5777: romdata_int <= 'h414; // Line Descriptor
    5778: romdata_int <= 'h1c00;
    5779: romdata_int <= 'h646;
    5780: romdata_int <= 'ha10;
    5781: romdata_int <= 'h414; // Line Descriptor
    5782: romdata_int <= 'h1e00;
    5783: romdata_int <= 'h34a;
    5784: romdata_int <= 'h703;
    5785: romdata_int <= 'h414; // Line Descriptor
    5786: romdata_int <= 'h2000;
    5787: romdata_int <= 'h133e;
    5788: romdata_int <= 'h12e4;
    5789: romdata_int <= 'h414; // Line Descriptor
    5790: romdata_int <= 'h2200;
    5791: romdata_int <= 'hcf2;
    5792: romdata_int <= 'h202c;
    5793: romdata_int <= 'h414; // Line Descriptor
    5794: romdata_int <= 'h2400;
    5795: romdata_int <= 'h1962;
    5796: romdata_int <= 'h935;
    5797: romdata_int <= 'h414; // Line Descriptor
    5798: romdata_int <= 'h2600;
    5799: romdata_int <= 'h952;
    5800: romdata_int <= 'hf64;
    5801: romdata_int <= 'h414; // Line Descriptor
    5802: romdata_int <= 'h0;
    5803: romdata_int <= 'h253d;
    5804: romdata_int <= 'h1661;
    5805: romdata_int <= 'h414; // Line Descriptor
    5806: romdata_int <= 'h200;
    5807: romdata_int <= 'h229b;
    5808: romdata_int <= 'h15c;
    5809: romdata_int <= 'h414; // Line Descriptor
    5810: romdata_int <= 'h400;
    5811: romdata_int <= 'h1487;
    5812: romdata_int <= 'h561;
    5813: romdata_int <= 'h414; // Line Descriptor
    5814: romdata_int <= 'h600;
    5815: romdata_int <= 'h1a38;
    5816: romdata_int <= 'h8b4;
    5817: romdata_int <= 'h414; // Line Descriptor
    5818: romdata_int <= 'h800;
    5819: romdata_int <= 'h1cb8;
    5820: romdata_int <= 'h2220;
    5821: romdata_int <= 'h414; // Line Descriptor
    5822: romdata_int <= 'ha00;
    5823: romdata_int <= 'h1e43;
    5824: romdata_int <= 'h1405;
    5825: romdata_int <= 'h414; // Line Descriptor
    5826: romdata_int <= 'hc00;
    5827: romdata_int <= 'h12a6;
    5828: romdata_int <= 'h2150;
    5829: romdata_int <= 'h414; // Line Descriptor
    5830: romdata_int <= 'he00;
    5831: romdata_int <= 'ha7d;
    5832: romdata_int <= 'heaa;
    5833: romdata_int <= 'h414; // Line Descriptor
    5834: romdata_int <= 'h1000;
    5835: romdata_int <= 'h47b;
    5836: romdata_int <= 'hcf0;
    5837: romdata_int <= 'h414; // Line Descriptor
    5838: romdata_int <= 'h1200;
    5839: romdata_int <= 'h20d2;
    5840: romdata_int <= 'h1c0a;
    5841: romdata_int <= 'h414; // Line Descriptor
    5842: romdata_int <= 'h1400;
    5843: romdata_int <= 'h110b;
    5844: romdata_int <= 'h2718;
    5845: romdata_int <= 'h414; // Line Descriptor
    5846: romdata_int <= 'h1600;
    5847: romdata_int <= 'hf4b;
    5848: romdata_int <= 'h738;
    5849: romdata_int <= 'h414; // Line Descriptor
    5850: romdata_int <= 'h1800;
    5851: romdata_int <= 'h884;
    5852: romdata_int <= 'h1afd;
    5853: romdata_int <= 'h414; // Line Descriptor
    5854: romdata_int <= 'h1a00;
    5855: romdata_int <= 'h18d2;
    5856: romdata_int <= 'h10fe;
    5857: romdata_int <= 'h414; // Line Descriptor
    5858: romdata_int <= 'h1c00;
    5859: romdata_int <= 'h6ad;
    5860: romdata_int <= 'h12c2;
    5861: romdata_int <= 'h414; // Line Descriptor
    5862: romdata_int <= 'h1e00;
    5863: romdata_int <= 'hd09;
    5864: romdata_int <= 'h2417;
    5865: romdata_int <= 'h414; // Line Descriptor
    5866: romdata_int <= 'h2000;
    5867: romdata_int <= 'hd8;
    5868: romdata_int <= 'h332;
    5869: romdata_int <= 'h414; // Line Descriptor
    5870: romdata_int <= 'h2200;
    5871: romdata_int <= 'h2c6;
    5872: romdata_int <= 'ha38;
    5873: romdata_int <= 'h414; // Line Descriptor
    5874: romdata_int <= 'h2400;
    5875: romdata_int <= 'h271c;
    5876: romdata_int <= 'h1e3b;
    5877: romdata_int <= 'h414; // Line Descriptor
    5878: romdata_int <= 'h2600;
    5879: romdata_int <= 'h1745;
    5880: romdata_int <= 'h1827;
    5881: romdata_int <= 'h414; // Line Descriptor
    5882: romdata_int <= 'h0;
    5883: romdata_int <= 'h1cc4;
    5884: romdata_int <= 'h248a;
    5885: romdata_int <= 'h414; // Line Descriptor
    5886: romdata_int <= 'h200;
    5887: romdata_int <= 'h24a1;
    5888: romdata_int <= 'hf49;
    5889: romdata_int <= 'h414; // Line Descriptor
    5890: romdata_int <= 'h400;
    5891: romdata_int <= 'h1637;
    5892: romdata_int <= 'h2149;
    5893: romdata_int <= 'h414; // Line Descriptor
    5894: romdata_int <= 'h600;
    5895: romdata_int <= 'h2248;
    5896: romdata_int <= 'hd37;
    5897: romdata_int <= 'h414; // Line Descriptor
    5898: romdata_int <= 'h800;
    5899: romdata_int <= 'hc48;
    5900: romdata_int <= 'hac2;
    5901: romdata_int <= 'h414; // Line Descriptor
    5902: romdata_int <= 'ha00;
    5903: romdata_int <= 'hec3;
    5904: romdata_int <= 'h6ca;
    5905: romdata_int <= 'h414; // Line Descriptor
    5906: romdata_int <= 'hc00;
    5907: romdata_int <= 'h2755;
    5908: romdata_int <= 'h1a8f;
    5909: romdata_int <= 'h414; // Line Descriptor
    5910: romdata_int <= 'he00;
    5911: romdata_int <= 'h1a56;
    5912: romdata_int <= 'h1f18;
    5913: romdata_int <= 'h414; // Line Descriptor
    5914: romdata_int <= 'h1000;
    5915: romdata_int <= 'h504;
    5916: romdata_int <= 'h12d5;
    5917: romdata_int <= 'h414; // Line Descriptor
    5918: romdata_int <= 'h1200;
    5919: romdata_int <= 'h897;
    5920: romdata_int <= 'h4ec;
    5921: romdata_int <= 'h414; // Line Descriptor
    5922: romdata_int <= 'h1400;
    5923: romdata_int <= 'hb10;
    5924: romdata_int <= 'h193e;
    5925: romdata_int <= 'h414; // Line Descriptor
    5926: romdata_int <= 'h1600;
    5927: romdata_int <= 'h1412;
    5928: romdata_int <= 'h105b;
    5929: romdata_int <= 'h414; // Line Descriptor
    5930: romdata_int <= 'h1800;
    5931: romdata_int <= 'h1eea;
    5932: romdata_int <= 'h50;
    5933: romdata_int <= 'h414; // Line Descriptor
    5934: romdata_int <= 'h1a00;
    5935: romdata_int <= 'h22;
    5936: romdata_int <= 'h1c67;
    5937: romdata_int <= 'h414; // Line Descriptor
    5938: romdata_int <= 'h1c00;
    5939: romdata_int <= 'h25a;
    5940: romdata_int <= 'h154e;
    5941: romdata_int <= 'h414; // Line Descriptor
    5942: romdata_int <= 'h1e00;
    5943: romdata_int <= 'h1285;
    5944: romdata_int <= 'h2244;
    5945: romdata_int <= 'h414; // Line Descriptor
    5946: romdata_int <= 'h2000;
    5947: romdata_int <= 'h67b;
    5948: romdata_int <= 'h254;
    5949: romdata_int <= 'h414; // Line Descriptor
    5950: romdata_int <= 'h2200;
    5951: romdata_int <= 'h192a;
    5952: romdata_int <= 'h1702;
    5953: romdata_int <= 'h414; // Line Descriptor
    5954: romdata_int <= 'h2400;
    5955: romdata_int <= 'h111e;
    5956: romdata_int <= 'h8d6;
    5957: romdata_int <= 'h514; // Line Descriptor
    5958: romdata_int <= 'h2600;
    5959: romdata_int <= 'h2054;
    5960: romdata_int <= 'h2648;
    5961: romdata_int <= 'h612; // Line Descriptor
    5962: romdata_int <= 'h0;
    5963: romdata_int <= 'h1b37;
    5964: romdata_int <= 'he8e;
    5965: romdata_int <= 'h4a1;
    5966: romdata_int <= 'h612; // Line Descriptor
    5967: romdata_int <= 'h200;
    5968: romdata_int <= 'h122;
    5969: romdata_int <= 'h16ae;
    5970: romdata_int <= 'hf0b;
    5971: romdata_int <= 'h612; // Line Descriptor
    5972: romdata_int <= 'h400;
    5973: romdata_int <= 'h1e89;
    5974: romdata_int <= 'hc2e;
    5975: romdata_int <= 'h1204;
    5976: romdata_int <= 'h612; // Line Descriptor
    5977: romdata_int <= 'h600;
    5978: romdata_int <= 'h35c;
    5979: romdata_int <= 'h1ce1;
    5980: romdata_int <= 'h22ec;
    5981: romdata_int <= 'h612; // Line Descriptor
    5982: romdata_int <= 'h800;
    5983: romdata_int <= 'h163a;
    5984: romdata_int <= 'h20a1;
    5985: romdata_int <= 'h939;
    5986: romdata_int <= 'h612; // Line Descriptor
    5987: romdata_int <= 'ha00;
    5988: romdata_int <= 'hc60;
    5989: romdata_int <= 'h879;
    5990: romdata_int <= 'h6b8;
    5991: romdata_int <= 'h612; // Line Descriptor
    5992: romdata_int <= 'hc00;
    5993: romdata_int <= 'h18b9;
    5994: romdata_int <= 'h113b;
    5995: romdata_int <= 'h1c7c;
    5996: romdata_int <= 'h612; // Line Descriptor
    5997: romdata_int <= 'he00;
    5998: romdata_int <= 'he79;
    5999: romdata_int <= 'h181e;
    6000: romdata_int <= 'h2bc;
    6001: romdata_int <= 'h612; // Line Descriptor
    6002: romdata_int <= 'h1000;
    6003: romdata_int <= 'ha91;
    6004: romdata_int <= 'h40d;
    6005: romdata_int <= 'hd28;
    6006: romdata_int <= 'h612; // Line Descriptor
    6007: romdata_int <= 'h1200;
    6008: romdata_int <= 'h2055;
    6009: romdata_int <= 'h1261;
    6010: romdata_int <= 'h18d5;
    6011: romdata_int <= 'h612; // Line Descriptor
    6012: romdata_int <= 'h1400;
    6013: romdata_int <= 'h1ce6;
    6014: romdata_int <= 'h2334;
    6015: romdata_int <= 'h14ae;
    6016: romdata_int <= 'h612; // Line Descriptor
    6017: romdata_int <= 'h1600;
    6018: romdata_int <= 'h10f3;
    6019: romdata_int <= 'haa4;
    6020: romdata_int <= 'h12c;
    6021: romdata_int <= 'h612; // Line Descriptor
    6022: romdata_int <= 'h1800;
    6023: romdata_int <= 'h643;
    6024: romdata_int <= 'h328;
    6025: romdata_int <= 'h16b0;
    6026: romdata_int <= 'h612; // Line Descriptor
    6027: romdata_int <= 'h1a00;
    6028: romdata_int <= 'h224e;
    6029: romdata_int <= 'hc4;
    6030: romdata_int <= 'h1f50;
    6031: romdata_int <= 'h612; // Line Descriptor
    6032: romdata_int <= 'h1c00;
    6033: romdata_int <= 'h852;
    6034: romdata_int <= 'h143b;
    6035: romdata_int <= 'h212b;
    6036: romdata_int <= 'h612; // Line Descriptor
    6037: romdata_int <= 'h1e00;
    6038: romdata_int <= 'h12d5;
    6039: romdata_int <= 'h1a62;
    6040: romdata_int <= 'h1af2;
    6041: romdata_int <= 'h612; // Line Descriptor
    6042: romdata_int <= 'h2000;
    6043: romdata_int <= 'h44a;
    6044: romdata_int <= 'h677;
    6045: romdata_int <= 'hae7;
    6046: romdata_int <= 'h612; // Line Descriptor
    6047: romdata_int <= 'h2200;
    6048: romdata_int <= 'h1483;
    6049: romdata_int <= 'h1f18;
    6050: romdata_int <= 'h100e;
    6051: romdata_int <= 'h412; // Line Descriptor
    6052: romdata_int <= 'h0;
    6053: romdata_int <= 'h2153;
    6054: romdata_int <= 'hb2c;
    6055: romdata_int <= 'h412; // Line Descriptor
    6056: romdata_int <= 'h200;
    6057: romdata_int <= 'hca6;
    6058: romdata_int <= 'h1cf2;
    6059: romdata_int <= 'h412; // Line Descriptor
    6060: romdata_int <= 'h400;
    6061: romdata_int <= 'h6bd;
    6062: romdata_int <= 'h1a5c;
    6063: romdata_int <= 'h412; // Line Descriptor
    6064: romdata_int <= 'h600;
    6065: romdata_int <= 'h1d01;
    6066: romdata_int <= 'hd34;
    6067: romdata_int <= 'h412; // Line Descriptor
    6068: romdata_int <= 'h800;
    6069: romdata_int <= 'h84b;
    6070: romdata_int <= 'h1ed9;
    6071: romdata_int <= 'h412; // Line Descriptor
    6072: romdata_int <= 'ha00;
    6073: romdata_int <= 'h1206;
    6074: romdata_int <= 'h65f;
    6075: romdata_int <= 'h412; // Line Descriptor
    6076: romdata_int <= 'hc00;
    6077: romdata_int <= 'hf2d;
    6078: romdata_int <= 'h89f;
    6079: romdata_int <= 'h412; // Line Descriptor
    6080: romdata_int <= 'he00;
    6081: romdata_int <= 'h234f;
    6082: romdata_int <= 'h2225;
    6083: romdata_int <= 'h412; // Line Descriptor
    6084: romdata_int <= 'h1000;
    6085: romdata_int <= 'h138;
    6086: romdata_int <= 'h108f;
    6087: romdata_int <= 'h412; // Line Descriptor
    6088: romdata_int <= 'h1200;
    6089: romdata_int <= 'h475;
    6090: romdata_int <= 'h1241;
    6091: romdata_int <= 'h412; // Line Descriptor
    6092: romdata_int <= 'h1400;
    6093: romdata_int <= 'h1e33;
    6094: romdata_int <= 'hf11;
    6095: romdata_int <= 'h412; // Line Descriptor
    6096: romdata_int <= 'h1600;
    6097: romdata_int <= 'h1b4a;
    6098: romdata_int <= 'h167d;
    6099: romdata_int <= 'h412; // Line Descriptor
    6100: romdata_int <= 'h1800;
    6101: romdata_int <= 'h104f;
    6102: romdata_int <= 'h305;
    6103: romdata_int <= 'h412; // Line Descriptor
    6104: romdata_int <= 'h1a00;
    6105: romdata_int <= 'h348;
    6106: romdata_int <= 'h181a;
    6107: romdata_int <= 'h412; // Line Descriptor
    6108: romdata_int <= 'h1c00;
    6109: romdata_int <= 'haee;
    6110: romdata_int <= 'h1466;
    6111: romdata_int <= 'h412; // Line Descriptor
    6112: romdata_int <= 'h1e00;
    6113: romdata_int <= 'h152a;
    6114: romdata_int <= 'h2158;
    6115: romdata_int <= 'h412; // Line Descriptor
    6116: romdata_int <= 'h2000;
    6117: romdata_int <= 'h1662;
    6118: romdata_int <= 'h4c1;
    6119: romdata_int <= 'h412; // Line Descriptor
    6120: romdata_int <= 'h2200;
    6121: romdata_int <= 'h18b2;
    6122: romdata_int <= 'h79;
    6123: romdata_int <= 'h412; // Line Descriptor
    6124: romdata_int <= 'h0;
    6125: romdata_int <= 'hee7;
    6126: romdata_int <= 'h431;
    6127: romdata_int <= 'h412; // Line Descriptor
    6128: romdata_int <= 'h200;
    6129: romdata_int <= 'h20a0;
    6130: romdata_int <= 'hd0;
    6131: romdata_int <= 'h412; // Line Descriptor
    6132: romdata_int <= 'h400;
    6133: romdata_int <= 'h1430;
    6134: romdata_int <= 'h169b;
    6135: romdata_int <= 'h412; // Line Descriptor
    6136: romdata_int <= 'h600;
    6137: romdata_int <= 'h6be;
    6138: romdata_int <= 'h2335;
    6139: romdata_int <= 'h412; // Line Descriptor
    6140: romdata_int <= 'h800;
    6141: romdata_int <= 'h4bd;
    6142: romdata_int <= 'hcc5;
    6143: romdata_int <= 'h412; // Line Descriptor
    6144: romdata_int <= 'ha00;
    6145: romdata_int <= 'h1c9f;
    6146: romdata_int <= 'hf32;
    6147: romdata_int <= 'h412; // Line Descriptor
    6148: romdata_int <= 'hc00;
    6149: romdata_int <= 'h181c;
    6150: romdata_int <= 'h125f;
    6151: romdata_int <= 'h412; // Line Descriptor
    6152: romdata_int <= 'he00;
    6153: romdata_int <= 'h122a;
    6154: romdata_int <= 'h1ac9;
    6155: romdata_int <= 'h412; // Line Descriptor
    6156: romdata_int <= 'h1000;
    6157: romdata_int <= 'h319;
    6158: romdata_int <= 'h250;
    6159: romdata_int <= 'h412; // Line Descriptor
    6160: romdata_int <= 'h1200;
    6161: romdata_int <= 'h1b38;
    6162: romdata_int <= 'h821;
    6163: romdata_int <= 'h412; // Line Descriptor
    6164: romdata_int <= 'h1400;
    6165: romdata_int <= 'hb2c;
    6166: romdata_int <= 'ha1a;
    6167: romdata_int <= 'h412; // Line Descriptor
    6168: romdata_int <= 'h1600;
    6169: romdata_int <= 'h1106;
    6170: romdata_int <= 'h1121;
    6171: romdata_int <= 'h412; // Line Descriptor
    6172: romdata_int <= 'h1800;
    6173: romdata_int <= 'h1608;
    6174: romdata_int <= 'h1c65;
    6175: romdata_int <= 'h412; // Line Descriptor
    6176: romdata_int <= 'h1a00;
    6177: romdata_int <= 'h1e5d;
    6178: romdata_int <= 'h1e7b;
    6179: romdata_int <= 'h412; // Line Descriptor
    6180: romdata_int <= 'h1c00;
    6181: romdata_int <= 'h2218;
    6182: romdata_int <= 'h1840;
    6183: romdata_int <= 'h412; // Line Descriptor
    6184: romdata_int <= 'h1e00;
    6185: romdata_int <= 'h880;
    6186: romdata_int <= 'h14ab;
    6187: romdata_int <= 'h412; // Line Descriptor
    6188: romdata_int <= 'h2000;
    6189: romdata_int <= 'hc3e;
    6190: romdata_int <= 'h625;
    6191: romdata_int <= 'h412; // Line Descriptor
    6192: romdata_int <= 'h2200;
    6193: romdata_int <= 'h7e;
    6194: romdata_int <= 'h213f;
    6195: romdata_int <= 'h412; // Line Descriptor
    6196: romdata_int <= 'h0;
    6197: romdata_int <= 'h1546;
    6198: romdata_int <= 'h2290;
    6199: romdata_int <= 'h412; // Line Descriptor
    6200: romdata_int <= 'h200;
    6201: romdata_int <= 'h102b;
    6202: romdata_int <= 'h16ba;
    6203: romdata_int <= 'h412; // Line Descriptor
    6204: romdata_int <= 'h400;
    6205: romdata_int <= 'he44;
    6206: romdata_int <= 'h2eb;
    6207: romdata_int <= 'h412; // Line Descriptor
    6208: romdata_int <= 'h600;
    6209: romdata_int <= 'h1aea;
    6210: romdata_int <= 'h72;
    6211: romdata_int <= 'h412; // Line Descriptor
    6212: romdata_int <= 'h800;
    6213: romdata_int <= 'h4ee;
    6214: romdata_int <= 'hec3;
    6215: romdata_int <= 'h412; // Line Descriptor
    6216: romdata_int <= 'ha00;
    6217: romdata_int <= 'hb33;
    6218: romdata_int <= 'h20b0;
    6219: romdata_int <= 'h412; // Line Descriptor
    6220: romdata_int <= 'hc00;
    6221: romdata_int <= 'h126b;
    6222: romdata_int <= 'hcfd;
    6223: romdata_int <= 'h412; // Line Descriptor
    6224: romdata_int <= 'he00;
    6225: romdata_int <= 'h841;
    6226: romdata_int <= 'ha07;
    6227: romdata_int <= 'h412; // Line Descriptor
    6228: romdata_int <= 'h1000;
    6229: romdata_int <= 'h2ad;
    6230: romdata_int <= 'h435;
    6231: romdata_int <= 'h412; // Line Descriptor
    6232: romdata_int <= 'h1200;
    6233: romdata_int <= 'h1ead;
    6234: romdata_int <= 'h103c;
    6235: romdata_int <= 'h412; // Line Descriptor
    6236: romdata_int <= 'h1400;
    6237: romdata_int <= 'h123;
    6238: romdata_int <= 'h18f6;
    6239: romdata_int <= 'h412; // Line Descriptor
    6240: romdata_int <= 'h1600;
    6241: romdata_int <= 'h213d;
    6242: romdata_int <= 'h1ced;
    6243: romdata_int <= 'h412; // Line Descriptor
    6244: romdata_int <= 'h1800;
    6245: romdata_int <= 'h18c4;
    6246: romdata_int <= 'h1e14;
    6247: romdata_int <= 'h412; // Line Descriptor
    6248: romdata_int <= 'h1a00;
    6249: romdata_int <= 'h160a;
    6250: romdata_int <= 'h149a;
    6251: romdata_int <= 'h412; // Line Descriptor
    6252: romdata_int <= 'h1c00;
    6253: romdata_int <= 'hc32;
    6254: romdata_int <= 'h8f6;
    6255: romdata_int <= 'h412; // Line Descriptor
    6256: romdata_int <= 'h1e00;
    6257: romdata_int <= 'h6b3;
    6258: romdata_int <= 'h1a3d;
    6259: romdata_int <= 'h412; // Line Descriptor
    6260: romdata_int <= 'h2000;
    6261: romdata_int <= 'h1d5d;
    6262: romdata_int <= 'h128f;
    6263: romdata_int <= 'h412; // Line Descriptor
    6264: romdata_int <= 'h2200;
    6265: romdata_int <= 'h2250;
    6266: romdata_int <= 'h632;
    6267: romdata_int <= 'h412; // Line Descriptor
    6268: romdata_int <= 'h0;
    6269: romdata_int <= 'h122f;
    6270: romdata_int <= 'h16f8;
    6271: romdata_int <= 'h412; // Line Descriptor
    6272: romdata_int <= 'h200;
    6273: romdata_int <= 'h16e3;
    6274: romdata_int <= 'h14dc;
    6275: romdata_int <= 'h412; // Line Descriptor
    6276: romdata_int <= 'h400;
    6277: romdata_int <= 'haf6;
    6278: romdata_int <= 'haf2;
    6279: romdata_int <= 'h412; // Line Descriptor
    6280: romdata_int <= 'h600;
    6281: romdata_int <= 'h1d20;
    6282: romdata_int <= 'h21e;
    6283: romdata_int <= 'h412; // Line Descriptor
    6284: romdata_int <= 'h800;
    6285: romdata_int <= 'h183f;
    6286: romdata_int <= 'h20f5;
    6287: romdata_int <= 'h412; // Line Descriptor
    6288: romdata_int <= 'ha00;
    6289: romdata_int <= 'h20b1;
    6290: romdata_int <= 'h8a1;
    6291: romdata_int <= 'h412; // Line Descriptor
    6292: romdata_int <= 'hc00;
    6293: romdata_int <= 'hc97;
    6294: romdata_int <= 'h61d;
    6295: romdata_int <= 'h412; // Line Descriptor
    6296: romdata_int <= 'he00;
    6297: romdata_int <= 'h63c;
    6298: romdata_int <= 'h4e5;
    6299: romdata_int <= 'h412; // Line Descriptor
    6300: romdata_int <= 'h1000;
    6301: romdata_int <= 'h881;
    6302: romdata_int <= 'h134d;
    6303: romdata_int <= 'h412; // Line Descriptor
    6304: romdata_int <= 'h1200;
    6305: romdata_int <= 'hf37;
    6306: romdata_int <= 'h1d4c;
    6307: romdata_int <= 'h412; // Line Descriptor
    6308: romdata_int <= 'h1400;
    6309: romdata_int <= 'h4f3;
    6310: romdata_int <= 'h1a57;
    6311: romdata_int <= 'h412; // Line Descriptor
    6312: romdata_int <= 'h1600;
    6313: romdata_int <= 'h1ef4;
    6314: romdata_int <= 'h1836;
    6315: romdata_int <= 'h412; // Line Descriptor
    6316: romdata_int <= 'h1800;
    6317: romdata_int <= 'h4a;
    6318: romdata_int <= 'hf56;
    6319: romdata_int <= 'h412; // Line Descriptor
    6320: romdata_int <= 'h1a00;
    6321: romdata_int <= 'h1b29;
    6322: romdata_int <= 'h1edc;
    6323: romdata_int <= 'h412; // Line Descriptor
    6324: romdata_int <= 'h1c00;
    6325: romdata_int <= 'h2269;
    6326: romdata_int <= 'h67;
    6327: romdata_int <= 'h412; // Line Descriptor
    6328: romdata_int <= 'h1e00;
    6329: romdata_int <= 'h2c8;
    6330: romdata_int <= 'hd3f;
    6331: romdata_int <= 'h412; // Line Descriptor
    6332: romdata_int <= 'h2000;
    6333: romdata_int <= 'h1150;
    6334: romdata_int <= 'h10b5;
    6335: romdata_int <= 'h412; // Line Descriptor
    6336: romdata_int <= 'h2200;
    6337: romdata_int <= 'h14b8;
    6338: romdata_int <= 'h22e2;
    6339: romdata_int <= 'h412; // Line Descriptor
    6340: romdata_int <= 'h0;
    6341: romdata_int <= 'h862;
    6342: romdata_int <= 'h8b4;
    6343: romdata_int <= 'h412; // Line Descriptor
    6344: romdata_int <= 'h200;
    6345: romdata_int <= 'he77;
    6346: romdata_int <= 'h8;
    6347: romdata_int <= 'h412; // Line Descriptor
    6348: romdata_int <= 'h400;
    6349: romdata_int <= 'ha58;
    6350: romdata_int <= 'heee;
    6351: romdata_int <= 'h412; // Line Descriptor
    6352: romdata_int <= 'h600;
    6353: romdata_int <= 'hd1e;
    6354: romdata_int <= 'h1445;
    6355: romdata_int <= 'h412; // Line Descriptor
    6356: romdata_int <= 'h800;
    6357: romdata_int <= 'h267;
    6358: romdata_int <= 'h2349;
    6359: romdata_int <= 'h412; // Line Descriptor
    6360: romdata_int <= 'ha00;
    6361: romdata_int <= 'h1d0b;
    6362: romdata_int <= 'hc96;
    6363: romdata_int <= 'h412; // Line Descriptor
    6364: romdata_int <= 'hc00;
    6365: romdata_int <= 'h2251;
    6366: romdata_int <= 'h18ba;
    6367: romdata_int <= 'h412; // Line Descriptor
    6368: romdata_int <= 'he00;
    6369: romdata_int <= 'hed;
    6370: romdata_int <= 'h1226;
    6371: romdata_int <= 'h412; // Line Descriptor
    6372: romdata_int <= 'h1000;
    6373: romdata_int <= 'h20e6;
    6374: romdata_int <= 'h470;
    6375: romdata_int <= 'h412; // Line Descriptor
    6376: romdata_int <= 'h1200;
    6377: romdata_int <= 'h1e74;
    6378: romdata_int <= 'h1c29;
    6379: romdata_int <= 'h412; // Line Descriptor
    6380: romdata_int <= 'h1400;
    6381: romdata_int <= 'h4ce;
    6382: romdata_int <= 'h2d6;
    6383: romdata_int <= 'h412; // Line Descriptor
    6384: romdata_int <= 'h1600;
    6385: romdata_int <= 'h171c;
    6386: romdata_int <= 'h1a33;
    6387: romdata_int <= 'h412; // Line Descriptor
    6388: romdata_int <= 'h1800;
    6389: romdata_int <= 'h1155;
    6390: romdata_int <= 'h16b8;
    6391: romdata_int <= 'h412; // Line Descriptor
    6392: romdata_int <= 'h1a00;
    6393: romdata_int <= 'h1a6b;
    6394: romdata_int <= 'h2115;
    6395: romdata_int <= 'h412; // Line Descriptor
    6396: romdata_int <= 'h1c00;
    6397: romdata_int <= 'h151d;
    6398: romdata_int <= 'h1e4f;
    6399: romdata_int <= 'h412; // Line Descriptor
    6400: romdata_int <= 'h1e00;
    6401: romdata_int <= 'h646;
    6402: romdata_int <= 'ha10;
    6403: romdata_int <= 'h412; // Line Descriptor
    6404: romdata_int <= 'h2000;
    6405: romdata_int <= 'h134a;
    6406: romdata_int <= 'h703;
    6407: romdata_int <= 'h412; // Line Descriptor
    6408: romdata_int <= 'h2200;
    6409: romdata_int <= 'h18fc;
    6410: romdata_int <= 'h1162;
    6411: romdata_int <= 'h412; // Line Descriptor
    6412: romdata_int <= 'h0;
    6413: romdata_int <= 'h6b0;
    6414: romdata_int <= 'h1504;
    6415: romdata_int <= 'h412; // Line Descriptor
    6416: romdata_int <= 'h200;
    6417: romdata_int <= 'h521;
    6418: romdata_int <= 'h1075;
    6419: romdata_int <= 'h412; // Line Descriptor
    6420: romdata_int <= 'h400;
    6421: romdata_int <= 'h1962;
    6422: romdata_int <= 'h735;
    6423: romdata_int <= 'h412; // Line Descriptor
    6424: romdata_int <= 'h600;
    6425: romdata_int <= 'h213d;
    6426: romdata_int <= 'h1661;
    6427: romdata_int <= 'h412; // Line Descriptor
    6428: romdata_int <= 'h800;
    6429: romdata_int <= 'h1e9b;
    6430: romdata_int <= 'h15c;
    6431: romdata_int <= 'h412; // Line Descriptor
    6432: romdata_int <= 'ha00;
    6433: romdata_int <= 'h1c42;
    6434: romdata_int <= 'hc91;
    6435: romdata_int <= 'h412; // Line Descriptor
    6436: romdata_int <= 'hc00;
    6437: romdata_int <= 'h1438;
    6438: romdata_int <= 'h8b4;
    6439: romdata_int <= 'h412; // Line Descriptor
    6440: romdata_int <= 'he00;
    6441: romdata_int <= 'h8df;
    6442: romdata_int <= 'h1f25;
    6443: romdata_int <= 'h412; // Line Descriptor
    6444: romdata_int <= 'h1000;
    6445: romdata_int <= 'he7d;
    6446: romdata_int <= 'heaa;
    6447: romdata_int <= 'h412; // Line Descriptor
    6448: romdata_int <= 'h1200;
    6449: romdata_int <= 'h2289;
    6450: romdata_int <= 'h1aaa;
    6451: romdata_int <= 'h412; // Line Descriptor
    6452: romdata_int <= 'h1400;
    6453: romdata_int <= 'h1042;
    6454: romdata_int <= 'h328;
    6455: romdata_int <= 'h412; // Line Descriptor
    6456: romdata_int <= 'h1600;
    6457: romdata_int <= 'h224;
    6458: romdata_int <= 'h18d9;
    6459: romdata_int <= 'h412; // Line Descriptor
    6460: romdata_int <= 'h1800;
    6461: romdata_int <= 'h16d2;
    6462: romdata_int <= 'h12fe;
    6463: romdata_int <= 'h412; // Line Descriptor
    6464: romdata_int <= 'h1a00;
    6465: romdata_int <= 'hd17;
    6466: romdata_int <= 'had3;
    6467: romdata_int <= 'h412; // Line Descriptor
    6468: romdata_int <= 'h1c00;
    6469: romdata_int <= 'haad;
    6470: romdata_int <= 'h1cc2;
    6471: romdata_int <= 'h412; // Line Descriptor
    6472: romdata_int <= 'h1e00;
    6473: romdata_int <= 'h1309;
    6474: romdata_int <= 'h2217;
    6475: romdata_int <= 'h412; // Line Descriptor
    6476: romdata_int <= 'h2000;
    6477: romdata_int <= 'hd8;
    6478: romdata_int <= 'h532;
    6479: romdata_int <= 'h412; // Line Descriptor
    6480: romdata_int <= 'h2200;
    6481: romdata_int <= 'h1af3;
    6482: romdata_int <= 'h20e2;
    6483: romdata_int <= 'h412; // Line Descriptor
    6484: romdata_int <= 'h0;
    6485: romdata_int <= 'h944;
    6486: romdata_int <= 'h5e;
    6487: romdata_int <= 'h412; // Line Descriptor
    6488: romdata_int <= 'h200;
    6489: romdata_int <= 'h1d1c;
    6490: romdata_int <= 'h203b;
    6491: romdata_int <= 'h412; // Line Descriptor
    6492: romdata_int <= 'h400;
    6493: romdata_int <= 'h1f3d;
    6494: romdata_int <= 'h1356;
    6495: romdata_int <= 'h412; // Line Descriptor
    6496: romdata_int <= 'h600;
    6497: romdata_int <= 'h18c4;
    6498: romdata_int <= 'h1e8a;
    6499: romdata_int <= 'h412; // Line Descriptor
    6500: romdata_int <= 'h800;
    6501: romdata_int <= 'h167b;
    6502: romdata_int <= 'h1960;
    6503: romdata_int <= 'h412; // Line Descriptor
    6504: romdata_int <= 'ha00;
    6505: romdata_int <= 'h3a;
    6506: romdata_int <= 'h1052;
    6507: romdata_int <= 'h412; // Line Descriptor
    6508: romdata_int <= 'hc00;
    6509: romdata_int <= 'hb5f;
    6510: romdata_int <= 'h14e0;
    6511: romdata_int <= 'h412; // Line Descriptor
    6512: romdata_int <= 'he00;
    6513: romdata_int <= 'h2248;
    6514: romdata_int <= 'hb37;
    6515: romdata_int <= 'h412; // Line Descriptor
    6516: romdata_int <= 'h1000;
    6517: romdata_int <= 'he48;
    6518: romdata_int <= 'h8c2;
    6519: romdata_int <= 'h412; // Line Descriptor
    6520: romdata_int <= 'h1200;
    6521: romdata_int <= 'hcc3;
    6522: romdata_int <= 'h6ca;
    6523: romdata_int <= 'h412; // Line Descriptor
    6524: romdata_int <= 'h1400;
    6525: romdata_int <= 'h1b1e;
    6526: romdata_int <= 'he7f;
    6527: romdata_int <= 'h412; // Line Descriptor
    6528: romdata_int <= 'h1600;
    6529: romdata_int <= 'h504;
    6530: romdata_int <= 'h16d5;
    6531: romdata_int <= 'h412; // Line Descriptor
    6532: romdata_int <= 'h1800;
    6533: romdata_int <= 'h6a9;
    6534: romdata_int <= 'h1a23;
    6535: romdata_int <= 'h412; // Line Descriptor
    6536: romdata_int <= 'h1a00;
    6537: romdata_int <= 'h149c;
    6538: romdata_int <= 'hc91;
    6539: romdata_int <= 'h412; // Line Descriptor
    6540: romdata_int <= 'h1c00;
    6541: romdata_int <= 'h12b5;
    6542: romdata_int <= 'h224;
    6543: romdata_int <= 'h412; // Line Descriptor
    6544: romdata_int <= 'h1e00;
    6545: romdata_int <= 'h115a;
    6546: romdata_int <= 'h2220;
    6547: romdata_int <= 'h412; // Line Descriptor
    6548: romdata_int <= 'h2000;
    6549: romdata_int <= 'h2023;
    6550: romdata_int <= 'h1ca3;
    6551: romdata_int <= 'h412; // Line Descriptor
    6552: romdata_int <= 'h2200;
    6553: romdata_int <= 'h2ea;
    6554: romdata_int <= 'h450;
    6555: romdata_int <= 'h412; // Line Descriptor
    6556: romdata_int <= 'h0;
    6557: romdata_int <= 'h341;
    6558: romdata_int <= 'h1858;
    6559: romdata_int <= 'h412; // Line Descriptor
    6560: romdata_int <= 'h200;
    6561: romdata_int <= 'h1285;
    6562: romdata_int <= 'h1a44;
    6563: romdata_int <= 'h412; // Line Descriptor
    6564: romdata_int <= 'h400;
    6565: romdata_int <= 'h67b;
    6566: romdata_int <= 'h454;
    6567: romdata_int <= 'h412; // Line Descriptor
    6568: romdata_int <= 'h600;
    6569: romdata_int <= 'h1737;
    6570: romdata_int <= 'h1c27;
    6571: romdata_int <= 'h412; // Line Descriptor
    6572: romdata_int <= 'h800;
    6573: romdata_int <= 'hf1e;
    6574: romdata_int <= 'hcd6;
    6575: romdata_int <= 'h412; // Line Descriptor
    6576: romdata_int <= 'ha00;
    6577: romdata_int <= 'ha54;
    6578: romdata_int <= 'h2048;
    6579: romdata_int <= 'h412; // Line Descriptor
    6580: romdata_int <= 'hc00;
    6581: romdata_int <= 'h208d;
    6582: romdata_int <= 'h10af;
    6583: romdata_int <= 'h412; // Line Descriptor
    6584: romdata_int <= 'he00;
    6585: romdata_int <= 'hd25;
    6586: romdata_int <= 'h1e92;
    6587: romdata_int <= 'h412; // Line Descriptor
    6588: romdata_int <= 'h1000;
    6589: romdata_int <= 'h915;
    6590: romdata_int <= 'h64b;
    6591: romdata_int <= 'h412; // Line Descriptor
    6592: romdata_int <= 'h1200;
    6593: romdata_int <= 'h1d39;
    6594: romdata_int <= 'h41;
    6595: romdata_int <= 'h412; // Line Descriptor
    6596: romdata_int <= 'h1400;
    6597: romdata_int <= 'h40;
    6598: romdata_int <= 'h14f2;
    6599: romdata_int <= 'h412; // Line Descriptor
    6600: romdata_int <= 'h1600;
    6601: romdata_int <= 'h1ec5;
    6602: romdata_int <= 'h92a;
    6603: romdata_int <= 'h412; // Line Descriptor
    6604: romdata_int <= 'h1800;
    6605: romdata_int <= 'h22c6;
    6606: romdata_int <= 'he4e;
    6607: romdata_int <= 'h412; // Line Descriptor
    6608: romdata_int <= 'h1a00;
    6609: romdata_int <= 'h1b39;
    6610: romdata_int <= 'h2302;
    6611: romdata_int <= 'h412; // Line Descriptor
    6612: romdata_int <= 'h1c00;
    6613: romdata_int <= 'h1855;
    6614: romdata_int <= 'h32c;
    6615: romdata_int <= 'h412; // Line Descriptor
    6616: romdata_int <= 'h1e00;
    6617: romdata_int <= 'h51a;
    6618: romdata_int <= 'ha95;
    6619: romdata_int <= 'h412; // Line Descriptor
    6620: romdata_int <= 'h2000;
    6621: romdata_int <= 'h1411;
    6622: romdata_int <= 'h1261;
    6623: romdata_int <= 'h512; // Line Descriptor
    6624: romdata_int <= 'h2200;
    6625: romdata_int <= 'h10bc;
    6626: romdata_int <= 'h166e;
    6627: romdata_int <= 'h1624; // Line Descriptor
    6628: romdata_int <= 'h3eae;
    6629: romdata_int <= 'h1d0b;
    6630: romdata_int <= 'h2008;
    6631: romdata_int <= 'h36d5;
    6632: romdata_int <= 'h1e86;
    6633: romdata_int <= 'h889;
    6634: romdata_int <= 'h82e;
    6635: romdata_int <= 'h4;
    6636: romdata_int <= 'hf37;
    6637: romdata_int <= 'h2e9a;
    6638: romdata_int <= 'h16b0;
    6639: romdata_int <= 'h3b5c;
    6640: romdata_int <= 'h1624; // Line Descriptor
    6641: romdata_int <= 'h4728;
    6642: romdata_int <= 'h288a;
    6643: romdata_int <= 'he6b;
    6644: romdata_int <= 'h3467;
    6645: romdata_int <= 'h1655;
    6646: romdata_int <= 'h461;
    6647: romdata_int <= 'h26d5;
    6648: romdata_int <= 'h231e;
    6649: romdata_int <= 'h30a5;
    6650: romdata_int <= 'hae0;
    6651: romdata_int <= 'h20e6;
    6652: romdata_int <= 'h534;
    6653: romdata_int <= 'h1624; // Line Descriptor
    6654: romdata_int <= 'h152b;
    6655: romdata_int <= 'h1a64;
    6656: romdata_int <= 'h3090;
    6657: romdata_int <= 'h2336;
    6658: romdata_int <= 'h10d5;
    6659: romdata_int <= 'h2a62;
    6660: romdata_int <= 'h44f2;
    6661: romdata_int <= 'h3eb6;
    6662: romdata_int <= 'h6c9;
    6663: romdata_int <= 'h3354;
    6664: romdata_int <= 'h144a;
    6665: romdata_int <= 'h1077;
    6666: romdata_int <= 'h1624; // Line Descriptor
    6667: romdata_int <= 'h3349;
    6668: romdata_int <= 'h67;
    6669: romdata_int <= 'haa6;
    6670: romdata_int <= 'hcf2;
    6671: romdata_int <= 'h1888;
    6672: romdata_int <= 'h3d27;
    6673: romdata_int <= 'h2bd;
    6674: romdata_int <= 'h2c5c;
    6675: romdata_int <= 'h4648;
    6676: romdata_int <= 'h2b22;
    6677: romdata_int <= 'h4301;
    6678: romdata_int <= 'h4134;
    6679: romdata_int <= 'h424; // Line Descriptor
    6680: romdata_int <= 'h40d9;
    6681: romdata_int <= 'h2655;
    6682: romdata_int <= 'h132b;
    6683: romdata_int <= 'h424; // Line Descriptor
    6684: romdata_int <= 'h25e;
    6685: romdata_int <= 'h252d;
    6686: romdata_int <= 'h2e9f;
    6687: romdata_int <= 'h424; // Line Descriptor
    6688: romdata_int <= 'h3825;
    6689: romdata_int <= 'h2d4d;
    6690: romdata_int <= 'h4552;
    6691: romdata_int <= 'h424; // Line Descriptor
    6692: romdata_int <= 'h42ab;
    6693: romdata_int <= 'h3a75;
    6694: romdata_int <= 'h641;
    6695: romdata_int <= 'h524; // Line Descriptor
    6696: romdata_int <= 'h1911;
    6697: romdata_int <= 'h2561;
    6698: romdata_int <= 'h128a;
    6699: romdata_int <= 'h161e; // Line Descriptor
    6700: romdata_int <= 'h340d;
    6701: romdata_int <= 'h3b28;
    6702: romdata_int <= 'h208a;
    6703: romdata_int <= 'hc6b;
    6704: romdata_int <= 'h2c67;
    6705: romdata_int <= 'h1455;
    6706: romdata_int <= 'h461;
    6707: romdata_int <= 'h1ed5;
    6708: romdata_int <= 'h1b1e;
    6709: romdata_int <= 'h26a5;
    6710: romdata_int <= 'h6e0;
    6711: romdata_int <= 'h18e6;
    6712: romdata_int <= 'h161e; // Line Descriptor
    6713: romdata_int <= 'h112b;
    6714: romdata_int <= 'h1664;
    6715: romdata_int <= 'h2690;
    6716: romdata_int <= 'h1936;
    6717: romdata_int <= 'hcd5;
    6718: romdata_int <= 'h2262;
    6719: romdata_int <= 'h38f2;
    6720: romdata_int <= 'h32b6;
    6721: romdata_int <= 'h2c9;
    6722: romdata_int <= 'h2554;
    6723: romdata_int <= 'hc4a;
    6724: romdata_int <= 'ha77;
    6725: romdata_int <= 'h161e; // Line Descriptor
    6726: romdata_int <= 'h2e70;
    6727: romdata_int <= 'h134f;
    6728: romdata_int <= 'h825;
    6729: romdata_int <= 'h254d;
    6730: romdata_int <= 'hf52;
    6731: romdata_int <= 'h3138;
    6732: romdata_int <= 'h8f;
    6733: romdata_int <= 'h1c0e;
    6734: romdata_int <= 'h12ab;
    6735: romdata_int <= 'h3475;
    6736: romdata_int <= 'h1e41;
    6737: romdata_int <= 'h164c;
    6738: romdata_int <= 'h161e; // Line Descriptor
    6739: romdata_int <= 'he5d;
    6740: romdata_int <= 'h67b;
    6741: romdata_int <= 'h32fd;
    6742: romdata_int <= 'h36eb;
    6743: romdata_int <= 'h2e18;
    6744: romdata_int <= 'h2a40;
    6745: romdata_int <= 'h2122;
    6746: romdata_int <= 'hacf;
    6747: romdata_int <= 'h80;
    6748: romdata_int <= 'h14ab;
    6749: romdata_int <= 'h2c98;
    6750: romdata_int <= 'h28b4;
    6751: romdata_int <= 'h161e; // Line Descriptor
    6752: romdata_int <= 'h28cb;
    6753: romdata_int <= 'h31d;
    6754: romdata_int <= 'h1e32;
    6755: romdata_int <= 'h30f6;
    6756: romdata_int <= 'h26a2;
    6757: romdata_int <= 'h34a4;
    6758: romdata_int <= 'h1ab3;
    6759: romdata_int <= 'h23d;
    6760: romdata_int <= 'h2a72;
    6761: romdata_int <= 'h3b3e;
    6762: romdata_int <= 'h55d;
    6763: romdata_int <= 'h208f;
    6764: romdata_int <= 'h41e; // Line Descriptor
    6765: romdata_int <= 'ha32;
    6766: romdata_int <= 'h18bd;
    6767: romdata_int <= 'h1103;
    6768: romdata_int <= 'h41e; // Line Descriptor
    6769: romdata_int <= 'h4ef;
    6770: romdata_int <= 'h28e3;
    6771: romdata_int <= 'h2edc;
    6772: romdata_int <= 'h41e; // Line Descriptor
    6773: romdata_int <= 'h2af2;
    6774: romdata_int <= 'h1683;
    6775: romdata_int <= 'h3274;
    6776: romdata_int <= 'h41e; // Line Descriptor
    6777: romdata_int <= 'h1556;
    6778: romdata_int <= 'h3b20;
    6779: romdata_int <= 'h1c1e;
    6780: romdata_int <= 'h41e; // Line Descriptor
    6781: romdata_int <= 'h2c78;
    6782: romdata_int <= 'h6fc;
    6783: romdata_int <= 'h3938;
    6784: romdata_int <= 'h41e; // Line Descriptor
    6785: romdata_int <= 'h14b;
    6786: romdata_int <= 'h24a8;
    6787: romdata_int <= 'h3097;
    6788: romdata_int <= 'h41e; // Line Descriptor
    6789: romdata_int <= 'h1ca1;
    6790: romdata_int <= 'h1340;
    6791: romdata_int <= 'he5a;
    6792: romdata_int <= 'h41e; // Line Descriptor
    6793: romdata_int <= 'h1ae5;
    6794: romdata_int <= 'h366b;
    6795: romdata_int <= 'h839;
    6796: romdata_int <= 'h41e; // Line Descriptor
    6797: romdata_int <= 'h389e;
    6798: romdata_int <= 'h1081;
    6799: romdata_int <= 'h374d;
    6800: romdata_int <= 'h51e; // Line Descriptor
    6801: romdata_int <= 'h2351;
    6802: romdata_int <= 'h86f;
    6803: romdata_int <= 'h2313;
    6804: romdata_int <= 'h161b; // Line Descriptor
    6805: romdata_int <= 'hed1;
    6806: romdata_int <= 'h1899;
    6807: romdata_int <= 'h544;
    6808: romdata_int <= 'h2015;
    6809: romdata_int <= 'h30f8;
    6810: romdata_int <= 'h332a;
    6811: romdata_int <= 'h1c17;
    6812: romdata_int <= 'h1841;
    6813: romdata_int <= 'h2a31;
    6814: romdata_int <= 'h1500;
    6815: romdata_int <= 'h121b;
    6816: romdata_int <= 'h20f6;
    6817: romdata_int <= 'h161b; // Line Descriptor
    6818: romdata_int <= 'h34d2;
    6819: romdata_int <= 'h163e;
    6820: romdata_int <= 'h2a76;
    6821: romdata_int <= 'h140f;
    6822: romdata_int <= 'h3503;
    6823: romdata_int <= 'h2ba;
    6824: romdata_int <= 'h26cf;
    6825: romdata_int <= 'h1a60;
    6826: romdata_int <= 'h281f;
    6827: romdata_int <= 'h700;
    6828: romdata_int <= 'h1e41;
    6829: romdata_int <= 'h3128;
    6830: romdata_int <= 'h161b; // Line Descriptor
    6831: romdata_int <= 'h2e93;
    6832: romdata_int <= 'h1e1c;
    6833: romdata_int <= 'h651;
    6834: romdata_int <= 'h2d0c;
    6835: romdata_int <= 'hd4c;
    6836: romdata_int <= 'h2120;
    6837: romdata_int <= 'h2842;
    6838: romdata_int <= 'h645;
    6839: romdata_int <= 'h10e3;
    6840: romdata_int <= 'h1947;
    6841: romdata_int <= 'h2c20;
    6842: romdata_int <= 'h1c47;
    6843: romdata_int <= 'h161b; // Line Descriptor
    6844: romdata_int <= 'h898;
    6845: romdata_int <= 'h28c;
    6846: romdata_int <= 'h2318;
    6847: romdata_int <= 'hcfc;
    6848: romdata_int <= 'hf59;
    6849: romdata_int <= 'h2530;
    6850: romdata_int <= 'h2ec7;
    6851: romdata_int <= 'h10d9;
    6852: romdata_int <= 'ha4;
    6853: romdata_int <= 'h3346;
    6854: romdata_int <= 'h231f;
    6855: romdata_int <= 'h1a53;
    6856: romdata_int <= 'h161b; // Line Descriptor
    6857: romdata_int <= 'h109d;
    6858: romdata_int <= 'h3020;
    6859: romdata_int <= 'h28a1;
    6860: romdata_int <= 'h2746;
    6861: romdata_int <= 'h2b65;
    6862: romdata_int <= 'hc;
    6863: romdata_int <= 'had9;
    6864: romdata_int <= 'h2cb0;
    6865: romdata_int <= 'h1608;
    6866: romdata_int <= 'hb24;
    6867: romdata_int <= 'hced;
    6868: romdata_int <= 'h354b;
    6869: romdata_int <= 'h161b; // Line Descriptor
    6870: romdata_int <= 'h167;
    6871: romdata_int <= 'h1c12;
    6872: romdata_int <= 'h125d;
    6873: romdata_int <= 'h1a52;
    6874: romdata_int <= 'h443;
    6875: romdata_int <= 'h1f59;
    6876: romdata_int <= 'h1647;
    6877: romdata_int <= 'h14be;
    6878: romdata_int <= 'he95;
    6879: romdata_int <= 'h24b2;
    6880: romdata_int <= 'h2e1d;
    6881: romdata_int <= 'h474;
    6882: romdata_int <= 'h41b; // Line Descriptor
    6883: romdata_int <= 'ha3d;
    6884: romdata_int <= 'h232e;
    6885: romdata_int <= 'h835;
    6886: romdata_int <= 'h41b; // Line Descriptor
    6887: romdata_int <= 'h247c;
    6888: romdata_int <= 'h12f2;
    6889: romdata_int <= 'h268a;
    6890: romdata_int <= 'h41b; // Line Descriptor
    6891: romdata_int <= 'h3357;
    6892: romdata_int <= 'h93b;
    6893: romdata_int <= 'h2ac;
    6894: romdata_int <= 'h41b; // Line Descriptor
    6895: romdata_int <= 'h3511;
    6896: romdata_int <= 'h18d6;
    6897: romdata_int <= 'h114c;
    6898: romdata_int <= 'h41b; // Line Descriptor
    6899: romdata_int <= 'h12f4;
    6900: romdata_int <= 'h2aa3;
    6901: romdata_int <= 'h2242;
    6902: romdata_int <= 'h41b; // Line Descriptor
    6903: romdata_int <= 'h1f57;
    6904: romdata_int <= 'h2495;
    6905: romdata_int <= 'h1a8e;
    6906: romdata_int <= 'h41b; // Line Descriptor
    6907: romdata_int <= 'h2141;
    6908: romdata_int <= 'hf11;
    6909: romdata_int <= 'hab7;
    6910: romdata_int <= 'h41b; // Line Descriptor
    6911: romdata_int <= 'h4c6;
    6912: romdata_int <= 'h2c49;
    6913: romdata_int <= 'hd54;
    6914: romdata_int <= 'h41b; // Line Descriptor
    6915: romdata_int <= 'h2f9;
    6916: romdata_int <= 'h314d;
    6917: romdata_int <= 'h6d1;
    6918: romdata_int <= 'h41b; // Line Descriptor
    6919: romdata_int <= 'h28a6;
    6920: romdata_int <= 'h16a4;
    6921: romdata_int <= 'h2f39;
    6922: romdata_int <= 'h41b; // Line Descriptor
    6923: romdata_int <= 'h8bd;
    6924: romdata_int <= 'h330f;
    6925: romdata_int <= 'h275d;
    6926: romdata_int <= 'h51b; // Line Descriptor
    6927: romdata_int <= 'h1433;
    6928: romdata_int <= 'h14a;
    6929: romdata_int <= 'h1c62;
    6930: romdata_int <= 'he19; // Line Descriptor
    6931: romdata_int <= 'h2800;
    6932: romdata_int <= 'h181c;
    6933: romdata_int <= 'h165f;
    6934: romdata_int <= 'h8fe;
    6935: romdata_int <= 'h16a2;
    6936: romdata_int <= 'h182a;
    6937: romdata_int <= 'h28c9;
    6938: romdata_int <= 'h10ce;
    6939: romdata_int <= 'he19; // Line Descriptor
    6940: romdata_int <= 'h2a00;
    6941: romdata_int <= 'h2465;
    6942: romdata_int <= 'h2ee5;
    6943: romdata_int <= 'h2cc0;
    6944: romdata_int <= 'h2e5d;
    6945: romdata_int <= 'h1c7b;
    6946: romdata_int <= 'h6fd;
    6947: romdata_int <= 'h2eb;
    6948: romdata_int <= 'he19; // Line Descriptor
    6949: romdata_int <= 'h2c00;
    6950: romdata_int <= 'h225;
    6951: romdata_int <= 'h2e4;
    6952: romdata_int <= 'h260a;
    6953: romdata_int <= 'h2493;
    6954: romdata_int <= 'h1a61;
    6955: romdata_int <= 'h1e7f;
    6956: romdata_int <= 'he8c;
    6957: romdata_int <= 'he19; // Line Descriptor
    6958: romdata_int <= 'h2e00;
    6959: romdata_int <= 'h470;
    6960: romdata_int <= 'h28b4;
    6961: romdata_int <= 'h48f;
    6962: romdata_int <= 'h30d4;
    6963: romdata_int <= 'h202b;
    6964: romdata_int <= 'h22ba;
    6965: romdata_int <= 'h30b1;
    6966: romdata_int <= 'he19; // Line Descriptor
    6967: romdata_int <= 'h3000;
    6968: romdata_int <= 'h1ecd;
    6969: romdata_int <= 'h650;
    6970: romdata_int <= 'h1a32;
    6971: romdata_int <= 'h22bd;
    6972: romdata_int <= 'h2d03;
    6973: romdata_int <= 'h142f;
    6974: romdata_int <= 'h4f8;
    6975: romdata_int <= 'h419; // Line Descriptor
    6976: romdata_int <= 'h0;
    6977: romdata_int <= 'h2aa1;
    6978: romdata_int <= 'h1315;
    6979: romdata_int <= 'h419; // Line Descriptor
    6980: romdata_int <= 'h200;
    6981: romdata_int <= 'ha72;
    6982: romdata_int <= 'h2002;
    6983: romdata_int <= 'h419; // Line Descriptor
    6984: romdata_int <= 'h400;
    6985: romdata_int <= 'h270b;
    6986: romdata_int <= 'h1808;
    6987: romdata_int <= 'h419; // Line Descriptor
    6988: romdata_int <= 'h600;
    6989: romdata_int <= 'h1c89;
    6990: romdata_int <= 'h102e;
    6991: romdata_int <= 'h419; // Line Descriptor
    6992: romdata_int <= 'h800;
    6993: romdata_int <= 'h9a;
    6994: romdata_int <= 'h2cb0;
    6995: romdata_int <= 'h419; // Line Descriptor
    6996: romdata_int <= 'ha00;
    6997: romdata_int <= 'h30ec;
    6998: romdata_int <= 'h1e0b;
    6999: romdata_int <= 'h419; // Line Descriptor
    7000: romdata_int <= 'hc00;
    7001: romdata_int <= 'h223a;
    7002: romdata_int <= 'h30a1;
    7003: romdata_int <= 'h419; // Line Descriptor
    7004: romdata_int <= 'he00;
    7005: romdata_int <= 'h2938;
    7006: romdata_int <= 'h2259;
    7007: romdata_int <= 'h419; // Line Descriptor
    7008: romdata_int <= 'h1000;
    7009: romdata_int <= 'hcb8;
    7010: romdata_int <= 'ha7b;
    7011: romdata_int <= 'h419; // Line Descriptor
    7012: romdata_int <= 'h1200;
    7013: romdata_int <= 'h10b9;
    7014: romdata_int <= 'h53b;
    7015: romdata_int <= 'h419; // Line Descriptor
    7016: romdata_int <= 'h1400;
    7017: romdata_int <= 'h129b;
    7018: romdata_int <= 'h2512;
    7019: romdata_int <= 'h419; // Line Descriptor
    7020: romdata_int <= 'h1600;
    7021: romdata_int <= 'h1565;
    7022: romdata_int <= 'h2ac7;
    7023: romdata_int <= 'h419; // Line Descriptor
    7024: romdata_int <= 'h1800;
    7025: romdata_int <= 'h679;
    7026: romdata_int <= 'h1c1e;
    7027: romdata_int <= 'h419; // Line Descriptor
    7028: romdata_int <= 'h1a00;
    7029: romdata_int <= 'h1aef;
    7030: romdata_int <= 'he2a;
    7031: romdata_int <= 'h519; // Line Descriptor
    7032: romdata_int <= 'h1c00;
    7033: romdata_int <= 'h1728;
    7034: romdata_int <= 'h8a;
    7035: romdata_int <= 'h1612; // Line Descriptor
    7036: romdata_int <= 'h1699;
    7037: romdata_int <= 'hf3d;
    7038: romdata_int <= 'h165;
    7039: romdata_int <= 'h1cc7;
    7040: romdata_int <= 'hc4c;
    7041: romdata_int <= 'hb0b;
    7042: romdata_int <= 'h879;
    7043: romdata_int <= 'h81e;
    7044: romdata_int <= 'h14bc;
    7045: romdata_int <= 'h1c9d;
    7046: romdata_int <= 'h10ef;
    7047: romdata_int <= 'h1e2a;
    7048: romdata_int <= 'h1612; // Line Descriptor
    7049: romdata_int <= 'h313;
    7050: romdata_int <= 'h1a0b;
    7051: romdata_int <= 'h187a;
    7052: romdata_int <= 'h628;
    7053: romdata_int <= 'h845;
    7054: romdata_int <= 'h18a2;
    7055: romdata_int <= 'h416;
    7056: romdata_int <= 'h1f3e;
    7057: romdata_int <= 'h1a0e;
    7058: romdata_int <= 'h737;
    7059: romdata_int <= 'h234c;
    7060: romdata_int <= 'ha91;
    7061: romdata_int <= 'h1612; // Line Descriptor
    7062: romdata_int <= 'h180b;
    7063: romdata_int <= 'h1d06;
    7064: romdata_int <= 'h2340;
    7065: romdata_int <= 'hac;
    7066: romdata_int <= 'h20ed;
    7067: romdata_int <= 'h155a;
    7068: romdata_int <= 'hf12;
    7069: romdata_int <= 'h63e;
    7070: romdata_int <= 'h367;
    7071: romdata_int <= 'hd26;
    7072: romdata_int <= 'h55f;
    7073: romdata_int <= 'h4df;
    7074: romdata_int <= 'h1612; // Line Descriptor
    7075: romdata_int <= 'h12e7;
    7076: romdata_int <= 'h1672;
    7077: romdata_int <= 'hb08;
    7078: romdata_int <= 'heaf;
    7079: romdata_int <= 'h193a;
    7080: romdata_int <= 'h1cdb;
    7081: romdata_int <= 'h1f4f;
    7082: romdata_int <= 'ha1f;
    7083: romdata_int <= 'hee;
    7084: romdata_int <= 'h1687;
    7085: romdata_int <= 'h14bd;
    7086: romdata_int <= 'h215f;
    7087: romdata_int <= 'h1612; // Line Descriptor
    7088: romdata_int <= 'hee9;
    7089: romdata_int <= 'h2086;
    7090: romdata_int <= 'h14f8;
    7091: romdata_int <= 'ha03;
    7092: romdata_int <= 'h165f;
    7093: romdata_int <= 'h2028;
    7094: romdata_int <= 'h12a6;
    7095: romdata_int <= 'h1c17;
    7096: romdata_int <= 'h12d3;
    7097: romdata_int <= 'h254;
    7098: romdata_int <= 'h2106;
    7099: romdata_int <= 'h758;
    7100: romdata_int <= 'h1612; // Line Descriptor
    7101: romdata_int <= 'hc94;
    7102: romdata_int <= 'h6ab;
    7103: romdata_int <= 'h131d;
    7104: romdata_int <= 'h14cf;
    7105: romdata_int <= 'h26f;
    7106: romdata_int <= 'h747;
    7107: romdata_int <= 'hcf2;
    7108: romdata_int <= 'h10d3;
    7109: romdata_int <= 'h20fb;
    7110: romdata_int <= 'h132c;
    7111: romdata_int <= 'h1962;
    7112: romdata_int <= 'h1b42;
    7113: romdata_int <= 'h1612; // Line Descriptor
    7114: romdata_int <= 'h1132;
    7115: romdata_int <= 'h45a;
    7116: romdata_int <= 'h10a1;
    7117: romdata_int <= 'h12b6;
    7118: romdata_int <= 'h1e45;
    7119: romdata_int <= 'h342;
    7120: romdata_int <= 'hd4;
    7121: romdata_int <= 'he2d;
    7122: romdata_int <= 'h1630;
    7123: romdata_int <= 'he80;
    7124: romdata_int <= 'h1ec4;
    7125: romdata_int <= 'h2242;
    7126: romdata_int <= 'h1612; // Line Descriptor
    7127: romdata_int <= 'h1ceb;
    7128: romdata_int <= 'hc79;
    7129: romdata_int <= 'h1f2c;
    7130: romdata_int <= 'h1a5e;
    7131: romdata_int <= 'h1139;
    7132: romdata_int <= 'h110f;
    7133: romdata_int <= 'h1681;
    7134: romdata_int <= 'h220f;
    7135: romdata_int <= 'h1866;
    7136: romdata_int <= 'ha3e;
    7137: romdata_int <= 'h1ac7;
    7138: romdata_int <= 'h154e;
    7139: romdata_int <= 'h1612; // Line Descriptor
    7140: romdata_int <= 'h77;
    7141: romdata_int <= 'h89d;
    7142: romdata_int <= 'h2e2;
    7143: romdata_int <= 'h53a;
    7144: romdata_int <= 'h2247;
    7145: romdata_int <= 'h22a3;
    7146: romdata_int <= 'h1ad9;
    7147: romdata_int <= 'hc4b;
    7148: romdata_int <= 'h431;
    7149: romdata_int <= 'h863;
    7150: romdata_int <= 'h16;
    7151: romdata_int <= 'h907;
    7152: romdata_int <= 'h412; // Line Descriptor
    7153: romdata_int <= 'h0;
    7154: romdata_int <= 'h278;
    7155: romdata_int <= 'he93;
    7156: romdata_int <= 'h412; // Line Descriptor
    7157: romdata_int <= 'h200;
    7158: romdata_int <= 'h184c;
    7159: romdata_int <= 'h651;
    7160: romdata_int <= 'h412; // Line Descriptor
    7161: romdata_int <= 'h400;
    7162: romdata_int <= 'h8b;
    7163: romdata_int <= 'h22cd;
    7164: romdata_int <= 'h412; // Line Descriptor
    7165: romdata_int <= 'h600;
    7166: romdata_int <= 'h16dc;
    7167: romdata_int <= 'h1a3a;
    7168: romdata_int <= 'h412; // Line Descriptor
    7169: romdata_int <= 'h800;
    7170: romdata_int <= 'h134c;
    7171: romdata_int <= 'h1d50;
    7172: romdata_int <= 'h412; // Line Descriptor
    7173: romdata_int <= 'ha00;
    7174: romdata_int <= 'ha60;
    7175: romdata_int <= 'h214e;
    7176: romdata_int <= 'h412; // Line Descriptor
    7177: romdata_int <= 'hc00;
    7178: romdata_int <= 'hcd2;
    7179: romdata_int <= 'h146b;
    7180: romdata_int <= 'h412; // Line Descriptor
    7181: romdata_int <= 'he00;
    7182: romdata_int <= 'h10ee;
    7183: romdata_int <= 'h435;
    7184: romdata_int <= 'h412; // Line Descriptor
    7185: romdata_int <= 'h1000;
    7186: romdata_int <= 'h93c;
    7187: romdata_int <= 'h1ebd;
    7188: romdata_int <= 'h412; // Line Descriptor
    7189: romdata_int <= 'h1200;
    7190: romdata_int <= 'h1c0e;
    7191: romdata_int <= 'h10f;
    7192: romdata_int <= 'h412; // Line Descriptor
    7193: romdata_int <= 'h1400;
    7194: romdata_int <= 'h2310;
    7195: romdata_int <= 'heb4;
    7196: romdata_int <= 'h412; // Line Descriptor
    7197: romdata_int <= 'h1600;
    7198: romdata_int <= 'h1708;
    7199: romdata_int <= 'h1ada;
    7200: romdata_int <= 'h412; // Line Descriptor
    7201: romdata_int <= 'h1800;
    7202: romdata_int <= 'h10c7;
    7203: romdata_int <= 'haa1;
    7204: romdata_int <= 'h412; // Line Descriptor
    7205: romdata_int <= 'h1a00;
    7206: romdata_int <= 'h148e;
    7207: romdata_int <= 'h6ea;
    7208: romdata_int <= 'h412; // Line Descriptor
    7209: romdata_int <= 'h1c00;
    7210: romdata_int <= 'hd21;
    7211: romdata_int <= 'h1305;
    7212: romdata_int <= 'h412; // Line Descriptor
    7213: romdata_int <= 'h1e00;
    7214: romdata_int <= 'h20da;
    7215: romdata_int <= 'h8bc;
    7216: romdata_int <= 'h412; // Line Descriptor
    7217: romdata_int <= 'h2000;
    7218: romdata_int <= 'h1f1b;
    7219: romdata_int <= 'h4fd;
    7220: romdata_int <= 'h512; // Line Descriptor
    7221: romdata_int <= 'h2200;
    7222: romdata_int <= 'h1910;
    7223: romdata_int <= 'h2e8;
    7224: romdata_int <= 'h180f; // Line Descriptor
    7225: romdata_int <= 'h0;
    7226: romdata_int <= 'h1c8a;
    7227: romdata_int <= 'h106b;
    7228: romdata_int <= 'h667;
    7229: romdata_int <= 'h1655;
    7230: romdata_int <= 'ha61;
    7231: romdata_int <= 'h2d5;
    7232: romdata_int <= 'hf1e;
    7233: romdata_int <= 'hca5;
    7234: romdata_int <= 'h12e0;
    7235: romdata_int <= 'h2e6;
    7236: romdata_int <= 'h134;
    7237: romdata_int <= 'h18ae;
    7238: romdata_int <= 'h180f; // Line Descriptor
    7239: romdata_int <= 'h200;
    7240: romdata_int <= 'h408;
    7241: romdata_int <= 'h265;
    7242: romdata_int <= 'h1ae5;
    7243: romdata_int <= 'hc0;
    7244: romdata_int <= 'h185d;
    7245: romdata_int <= 'h47b;
    7246: romdata_int <= 'h8fd;
    7247: romdata_int <= 'h8eb;
    7248: romdata_int <= 'h1a18;
    7249: romdata_int <= 'h1640;
    7250: romdata_int <= 'h1122;
    7251: romdata_int <= 'h6cf;
    7252: romdata_int <= 'h180f; // Line Descriptor
    7253: romdata_int <= 'h400;
    7254: romdata_int <= 'h811;
    7255: romdata_int <= 'h12e2;
    7256: romdata_int <= 'h1c3d;
    7257: romdata_int <= 'h14b0;
    7258: romdata_int <= 'h1239;
    7259: romdata_int <= 'hd0a;
    7260: romdata_int <= 'h10ff;
    7261: romdata_int <= 'h407;
    7262: romdata_int <= 'hf60;
    7263: romdata_int <= 'h1c0a;
    7264: romdata_int <= 'had0;
    7265: romdata_int <= 'h149c;
    7266: romdata_int <= 'h40f; // Line Descriptor
    7267: romdata_int <= 'h600;
    7268: romdata_int <= 'h1816;
    7269: romdata_int <= 'h8eb;
    7270: romdata_int <= 'h40f; // Line Descriptor
    7271: romdata_int <= 'h800;
    7272: romdata_int <= 'h1b17;
    7273: romdata_int <= 'h48f;
    7274: romdata_int <= 'h40f; // Line Descriptor
    7275: romdata_int <= 'ha00;
    7276: romdata_int <= 'ha7d;
    7277: romdata_int <= 'hd42;
    7278: romdata_int <= 'h40f; // Line Descriptor
    7279: romdata_int <= 'hc00;
    7280: romdata_int <= 'h1301;
    7281: romdata_int <= 'hb47;
    7282: romdata_int <= 'h40f; // Line Descriptor
    7283: romdata_int <= 'he00;
    7284: romdata_int <= 'h610;
    7285: romdata_int <= 'h1866;
    7286: romdata_int <= 'h40f; // Line Descriptor
    7287: romdata_int <= 'h1000;
    7288: romdata_int <= 'h16c8;
    7289: romdata_int <= 'h165f;
    7290: romdata_int <= 'h40f; // Line Descriptor
    7291: romdata_int <= 'h1200;
    7292: romdata_int <= 'he90;
    7293: romdata_int <= 'hea7;
    7294: romdata_int <= 'h40f; // Line Descriptor
    7295: romdata_int <= 'h1400;
    7296: romdata_int <= 'h333;
    7297: romdata_int <= 'h1a42;
    7298: romdata_int <= 'h40f; // Line Descriptor
    7299: romdata_int <= 'h1600;
    7300: romdata_int <= 'hbd;
    7301: romdata_int <= 'h2f;
    7302: romdata_int <= 'h40f; // Line Descriptor
    7303: romdata_int <= 'h1800;
    7304: romdata_int <= 'hce4;
    7305: romdata_int <= 'h149d;
    7306: romdata_int <= 'h40f; // Line Descriptor
    7307: romdata_int <= 'h1a00;
    7308: romdata_int <= 'h1100;
    7309: romdata_int <= 'h1ca4;
    7310: romdata_int <= 'h40f; // Line Descriptor
    7311: romdata_int <= 'h1c00;
    7312: romdata_int <= 'h145a;
    7313: romdata_int <= 'h674;
    7314: romdata_int <= 'h40f; // Line Descriptor
    7315: romdata_int <= 'h0;
    7316: romdata_int <= 'h1a0a;
    7317: romdata_int <= 'h2a9;
    7318: romdata_int <= 'h40f; // Line Descriptor
    7319: romdata_int <= 'h200;
    7320: romdata_int <= 'h6ac;
    7321: romdata_int <= 'h144e;
    7322: romdata_int <= 'h40f; // Line Descriptor
    7323: romdata_int <= 'h400;
    7324: romdata_int <= 'h1866;
    7325: romdata_int <= 'h1c21;
    7326: romdata_int <= 'h40f; // Line Descriptor
    7327: romdata_int <= 'h600;
    7328: romdata_int <= 'h1126;
    7329: romdata_int <= 'h43;
    7330: romdata_int <= 'h40f; // Line Descriptor
    7331: romdata_int <= 'h800;
    7332: romdata_int <= 'hf5b;
    7333: romdata_int <= 'h555;
    7334: romdata_int <= 'h40f; // Line Descriptor
    7335: romdata_int <= 'ha00;
    7336: romdata_int <= 'h148f;
    7337: romdata_int <= 'h18c2;
    7338: romdata_int <= 'h40f; // Line Descriptor
    7339: romdata_int <= 'hc00;
    7340: romdata_int <= 'h417;
    7341: romdata_int <= 'h16b3;
    7342: romdata_int <= 'h40f; // Line Descriptor
    7343: romdata_int <= 'he00;
    7344: romdata_int <= 'h20f;
    7345: romdata_int <= 'hd1e;
    7346: romdata_int <= 'h40f; // Line Descriptor
    7347: romdata_int <= 'h1000;
    7348: romdata_int <= 'h68;
    7349: romdata_int <= 'he20;
    7350: romdata_int <= 'h40f; // Line Descriptor
    7351: romdata_int <= 'h1200;
    7352: romdata_int <= 'h1705;
    7353: romdata_int <= 'ha6d;
    7354: romdata_int <= 'h40f; // Line Descriptor
    7355: romdata_int <= 'h1400;
    7356: romdata_int <= 'h1c09;
    7357: romdata_int <= 'h6c3;
    7358: romdata_int <= 'h40f; // Line Descriptor
    7359: romdata_int <= 'h1600;
    7360: romdata_int <= 'h129d;
    7361: romdata_int <= 'h1025;
    7362: romdata_int <= 'h40f; // Line Descriptor
    7363: romdata_int <= 'h1800;
    7364: romdata_int <= 'ha2a;
    7365: romdata_int <= 'h1a2d;
    7366: romdata_int <= 'h40f; // Line Descriptor
    7367: romdata_int <= 'h1a00;
    7368: romdata_int <= 'hc0f;
    7369: romdata_int <= 'h870;
    7370: romdata_int <= 'h50f; // Line Descriptor
    7371: romdata_int <= 'h1c00;
    7372: romdata_int <= 'h84b;
    7373: romdata_int <= 'h1303;
    7374: romdata_int <= 'h160c; // Line Descriptor
    7375: romdata_int <= 'h600;
    7376: romdata_int <= 'hd0a;
    7377: romdata_int <= 'h1427;
    7378: romdata_int <= 'hf5e;
    7379: romdata_int <= 'ha7b;
    7380: romdata_int <= 'h254;
    7381: romdata_int <= 'hda;
    7382: romdata_int <= 'h8a0;
    7383: romdata_int <= 'hb1e;
    7384: romdata_int <= 'h42e;
    7385: romdata_int <= 'h1638;
    7386: romdata_int <= 'h296;
    7387: romdata_int <= 'h40c; // Line Descriptor
    7388: romdata_int <= 'h800;
    7389: romdata_int <= 'hadf;
    7390: romdata_int <= 'h16b1;
    7391: romdata_int <= 'h40c; // Line Descriptor
    7392: romdata_int <= 'ha00;
    7393: romdata_int <= 'h1702;
    7394: romdata_int <= 'hf4f;
    7395: romdata_int <= 'h40c; // Line Descriptor
    7396: romdata_int <= 'hc00;
    7397: romdata_int <= 'h12db;
    7398: romdata_int <= 'h319;
    7399: romdata_int <= 'h40c; // Line Descriptor
    7400: romdata_int <= 'he00;
    7401: romdata_int <= 'h53f;
    7402: romdata_int <= 'hb1f;
    7403: romdata_int <= 'h40c; // Line Descriptor
    7404: romdata_int <= 'h1000;
    7405: romdata_int <= 'h358;
    7406: romdata_int <= 'h10ab;
    7407: romdata_int <= 'h40c; // Line Descriptor
    7408: romdata_int <= 'h1200;
    7409: romdata_int <= 'h115c;
    7410: romdata_int <= 'hce4;
    7411: romdata_int <= 'h40c; // Line Descriptor
    7412: romdata_int <= 'h1400;
    7413: romdata_int <= 'h1548;
    7414: romdata_int <= 'h459;
    7415: romdata_int <= 'h40c; // Line Descriptor
    7416: romdata_int <= 'h1600;
    7417: romdata_int <= 'heba;
    7418: romdata_int <= 'h52;
    7419: romdata_int <= 'h40c; // Line Descriptor
    7420: romdata_int <= 'h0;
    7421: romdata_int <= 'hc79;
    7422: romdata_int <= 'hefc;
    7423: romdata_int <= 'h40c; // Line Descriptor
    7424: romdata_int <= 'h200;
    7425: romdata_int <= 'h6fa;
    7426: romdata_int <= 'h106e;
    7427: romdata_int <= 'h40c; // Line Descriptor
    7428: romdata_int <= 'h400;
    7429: romdata_int <= 'h125e;
    7430: romdata_int <= 'h8f;
    7431: romdata_int <= 'h40c; // Line Descriptor
    7432: romdata_int <= 'h600;
    7433: romdata_int <= 'hb;
    7434: romdata_int <= 'hb36;
    7435: romdata_int <= 'h40c; // Line Descriptor
    7436: romdata_int <= 'h800;
    7437: romdata_int <= 'ha97;
    7438: romdata_int <= 'h435;
    7439: romdata_int <= 'h40c; // Line Descriptor
    7440: romdata_int <= 'ha00;
    7441: romdata_int <= 'h1493;
    7442: romdata_int <= 'h71f;
    7443: romdata_int <= 'h40c; // Line Descriptor
    7444: romdata_int <= 'hc00;
    7445: romdata_int <= 'h112e;
    7446: romdata_int <= 'h1268;
    7447: romdata_int <= 'h40c; // Line Descriptor
    7448: romdata_int <= 'he00;
    7449: romdata_int <= 'h42d;
    7450: romdata_int <= 'h1533;
    7451: romdata_int <= 'h40c; // Line Descriptor
    7452: romdata_int <= 'h1000;
    7453: romdata_int <= 'he54;
    7454: romdata_int <= 'h2a2;
    7455: romdata_int <= 'h40c; // Line Descriptor
    7456: romdata_int <= 'h1200;
    7457: romdata_int <= 'h8a2;
    7458: romdata_int <= 'h822;
    7459: romdata_int <= 'h40c; // Line Descriptor
    7460: romdata_int <= 'h1400;
    7461: romdata_int <= 'h1652;
    7462: romdata_int <= 'hcba;
    7463: romdata_int <= 'h40c; // Line Descriptor
    7464: romdata_int <= 'h1600;
    7465: romdata_int <= 'h359;
    7466: romdata_int <= 'h169e;
    7467: romdata_int <= 'h40c; // Line Descriptor
    7468: romdata_int <= 'h0;
    7469: romdata_int <= 'h10ce;
    7470: romdata_int <= 'hf00;
    7471: romdata_int <= 'h40c; // Line Descriptor
    7472: romdata_int <= 'h200;
    7473: romdata_int <= 'h12fb;
    7474: romdata_int <= 'h105a;
    7475: romdata_int <= 'h40c; // Line Descriptor
    7476: romdata_int <= 'h400;
    7477: romdata_int <= 'ha3b;
    7478: romdata_int <= 'h1672;
    7479: romdata_int <= 'h40c; // Line Descriptor
    7480: romdata_int <= 'h600;
    7481: romdata_int <= 'h253;
    7482: romdata_int <= 'h745;
    7483: romdata_int <= 'h40c; // Line Descriptor
    7484: romdata_int <= 'h800;
    7485: romdata_int <= 'hec1;
    7486: romdata_int <= 'h318;
    7487: romdata_int <= 'h40c; // Line Descriptor
    7488: romdata_int <= 'ha00;
    7489: romdata_int <= 'hc5c;
    7490: romdata_int <= 'h452;
    7491: romdata_int <= 'h40c; // Line Descriptor
    7492: romdata_int <= 'hc00;
    7493: romdata_int <= 'hd3;
    7494: romdata_int <= 'h140b;
    7495: romdata_int <= 'h40c; // Line Descriptor
    7496: romdata_int <= 'he00;
    7497: romdata_int <= 'h148c;
    7498: romdata_int <= 'hac8;
    7499: romdata_int <= 'h40c; // Line Descriptor
    7500: romdata_int <= 'h1000;
    7501: romdata_int <= 'h46c;
    7502: romdata_int <= 'h129c;
    7503: romdata_int <= 'h40c; // Line Descriptor
    7504: romdata_int <= 'h1200;
    7505: romdata_int <= 'h633;
    7506: romdata_int <= 'hc0e;
    7507: romdata_int <= 'h40c; // Line Descriptor
    7508: romdata_int <= 'h1400;
    7509: romdata_int <= 'h889;
    7510: romdata_int <= 'h903;
    7511: romdata_int <= 'h50c; // Line Descriptor
    7512: romdata_int <= 'h1600;
    7513: romdata_int <= 'h1675;
    7514: romdata_int <= 'hea;
    7515: romdata_int <= 'h40a; // Line Descriptor
    7516: romdata_int <= 'ha00;
    7517: romdata_int <= 'hc59;
    7518: romdata_int <= 'ha9c;
    7519: romdata_int <= 'h40a; // Line Descriptor
    7520: romdata_int <= 'hc00;
    7521: romdata_int <= 'h6f9;
    7522: romdata_int <= 'h812;
    7523: romdata_int <= 'h40a; // Line Descriptor
    7524: romdata_int <= 'he00;
    7525: romdata_int <= 'h415;
    7526: romdata_int <= 'h141;
    7527: romdata_int <= 'h40a; // Line Descriptor
    7528: romdata_int <= 'h1000;
    7529: romdata_int <= 'he48;
    7530: romdata_int <= 'h1285;
    7531: romdata_int <= 'h40a; // Line Descriptor
    7532: romdata_int <= 'h1200;
    7533: romdata_int <= 'h1156;
    7534: romdata_int <= 'h43d;
    7535: romdata_int <= 'h40a; // Line Descriptor
    7536: romdata_int <= 'h0;
    7537: romdata_int <= 'h70a;
    7538: romdata_int <= 'hec2;
    7539: romdata_int <= 'h40a; // Line Descriptor
    7540: romdata_int <= 'h200;
    7541: romdata_int <= 'h17;
    7542: romdata_int <= 'hb0d;
    7543: romdata_int <= 'h40a; // Line Descriptor
    7544: romdata_int <= 'h400;
    7545: romdata_int <= 'haca;
    7546: romdata_int <= 'h917;
    7547: romdata_int <= 'h40a; // Line Descriptor
    7548: romdata_int <= 'h600;
    7549: romdata_int <= 'h132f;
    7550: romdata_int <= 'h61c;
    7551: romdata_int <= 'h40a; // Line Descriptor
    7552: romdata_int <= 'h800;
    7553: romdata_int <= 'h456;
    7554: romdata_int <= 'h1320;
    7555: romdata_int <= 'h40a; // Line Descriptor
    7556: romdata_int <= 'ha00;
    7557: romdata_int <= 'hc25;
    7558: romdata_int <= 'hd3;
    7559: romdata_int <= 'h40a; // Line Descriptor
    7560: romdata_int <= 'hc00;
    7561: romdata_int <= 'h8cb;
    7562: romdata_int <= 'hce4;
    7563: romdata_int <= 'h40a; // Line Descriptor
    7564: romdata_int <= 'he00;
    7565: romdata_int <= 'h25f;
    7566: romdata_int <= 'h10ce;
    7567: romdata_int <= 'h40a; // Line Descriptor
    7568: romdata_int <= 'h1000;
    7569: romdata_int <= 'h1136;
    7570: romdata_int <= 'h562;
    7571: romdata_int <= 'h40a; // Line Descriptor
    7572: romdata_int <= 'h1200;
    7573: romdata_int <= 'he1e;
    7574: romdata_int <= 'h28e;
    7575: romdata_int <= 'h40a; // Line Descriptor
    7576: romdata_int <= 'h0;
    7577: romdata_int <= 'h4e3;
    7578: romdata_int <= 'he77;
    7579: romdata_int <= 'h40a; // Line Descriptor
    7580: romdata_int <= 'h200;
    7581: romdata_int <= 'hb4;
    7582: romdata_int <= 'h148;
    7583: romdata_int <= 'h40a; // Line Descriptor
    7584: romdata_int <= 'h400;
    7585: romdata_int <= 'h221;
    7586: romdata_int <= 'h10e6;
    7587: romdata_int <= 'h40a; // Line Descriptor
    7588: romdata_int <= 'h600;
    7589: romdata_int <= 'ha2e;
    7590: romdata_int <= 'h4ff;
    7591: romdata_int <= 'h40a; // Line Descriptor
    7592: romdata_int <= 'h800;
    7593: romdata_int <= 'h1067;
    7594: romdata_int <= 'h12f7;
    7595: romdata_int <= 'h40a; // Line Descriptor
    7596: romdata_int <= 'ha00;
    7597: romdata_int <= 'h68a;
    7598: romdata_int <= 'h622;
    7599: romdata_int <= 'h40a; // Line Descriptor
    7600: romdata_int <= 'hc00;
    7601: romdata_int <= 'h809;
    7602: romdata_int <= 'hc17;
    7603: romdata_int <= 'h40a; // Line Descriptor
    7604: romdata_int <= 'he00;
    7605: romdata_int <= 'h1305;
    7606: romdata_int <= 'h20c;
    7607: romdata_int <= 'h40a; // Line Descriptor
    7608: romdata_int <= 'h1000;
    7609: romdata_int <= 'he95;
    7610: romdata_int <= 'h915;
    7611: romdata_int <= 'h40a; // Line Descriptor
    7612: romdata_int <= 'h1200;
    7613: romdata_int <= 'hcd3;
    7614: romdata_int <= 'hab9;
    7615: romdata_int <= 'h40a; // Line Descriptor
    7616: romdata_int <= 'h0;
    7617: romdata_int <= 'h448;
    7618: romdata_int <= 'h89e;
    7619: romdata_int <= 'h40a; // Line Descriptor
    7620: romdata_int <= 'h200;
    7621: romdata_int <= 'hf14;
    7622: romdata_int <= 'h2bc;
    7623: romdata_int <= 'h40a; // Line Descriptor
    7624: romdata_int <= 'h400;
    7625: romdata_int <= 'h30e;
    7626: romdata_int <= 'ha1;
    7627: romdata_int <= 'h40a; // Line Descriptor
    7628: romdata_int <= 'h600;
    7629: romdata_int <= 'h748;
    7630: romdata_int <= 'h4ad;
    7631: romdata_int <= 'h40a; // Line Descriptor
    7632: romdata_int <= 'h800;
    7633: romdata_int <= 'h1010;
    7634: romdata_int <= 'h126d;
    7635: romdata_int <= 'h40a; // Line Descriptor
    7636: romdata_int <= 'ha00;
    7637: romdata_int <= 'h933;
    7638: romdata_int <= 'h618;
    7639: romdata_int <= 'h40a; // Line Descriptor
    7640: romdata_int <= 'hc00;
    7641: romdata_int <= 'h15a;
    7642: romdata_int <= 'ha5e;
    7643: romdata_int <= 'h40a; // Line Descriptor
    7644: romdata_int <= 'he00;
    7645: romdata_int <= 'h12cc;
    7646: romdata_int <= 'hcae;
    7647: romdata_int <= 'h40a; // Line Descriptor
    7648: romdata_int <= 'h1000;
    7649: romdata_int <= 'hc38;
    7650: romdata_int <= 'he8e;
    7651: romdata_int <= 'h50a; // Line Descriptor
    7652: romdata_int <= 'h1200;
    7653: romdata_int <= 'hb62;
    7654: romdata_int <= 'h1074;
    7655: romdata_int <= 'h1808; // Line Descriptor
    7656: romdata_int <= 'h600;
    7657: romdata_int <= 'h32d;
    7658: romdata_int <= 'h63e;
    7659: romdata_int <= 'h2b9;
    7660: romdata_int <= 'h871;
    7661: romdata_int <= 'he45;
    7662: romdata_int <= 'h859;
    7663: romdata_int <= 'hc9e;
    7664: romdata_int <= 'ha29;
    7665: romdata_int <= 'h939;
    7666: romdata_int <= 'h11b;
    7667: romdata_int <= 'hcd4;
    7668: romdata_int <= 'hb5e;
    7669: romdata_int <= 'h408; // Line Descriptor
    7670: romdata_int <= 'h800;
    7671: romdata_int <= 'hf31;
    7672: romdata_int <= 'hcf0;
    7673: romdata_int <= 'h408; // Line Descriptor
    7674: romdata_int <= 'ha00;
    7675: romdata_int <= 'hc33;
    7676: romdata_int <= 'h99;
    7677: romdata_int <= 'h408; // Line Descriptor
    7678: romdata_int <= 'hc00;
    7679: romdata_int <= 'h508;
    7680: romdata_int <= 'h469;
    7681: romdata_int <= 'h408; // Line Descriptor
    7682: romdata_int <= 'he00;
    7683: romdata_int <= 'h81a;
    7684: romdata_int <= 'ha47;
    7685: romdata_int <= 'h408; // Line Descriptor
    7686: romdata_int <= 'h0;
    7687: romdata_int <= 'hf29;
    7688: romdata_int <= 'h108;
    7689: romdata_int <= 'h408; // Line Descriptor
    7690: romdata_int <= 'h200;
    7691: romdata_int <= 'hd1d;
    7692: romdata_int <= 'h925;
    7693: romdata_int <= 'h408; // Line Descriptor
    7694: romdata_int <= 'h400;
    7695: romdata_int <= 'h244;
    7696: romdata_int <= 'h666;
    7697: romdata_int <= 'h408; // Line Descriptor
    7698: romdata_int <= 'h600;
    7699: romdata_int <= 'h9e;
    7700: romdata_int <= 'he11;
    7701: romdata_int <= 'h408; // Line Descriptor
    7702: romdata_int <= 'h800;
    7703: romdata_int <= 'had4;
    7704: romdata_int <= 'h51a;
    7705: romdata_int <= 'h408; // Line Descriptor
    7706: romdata_int <= 'ha00;
    7707: romdata_int <= 'h878;
    7708: romdata_int <= 'hc14;
    7709: romdata_int <= 'h408; // Line Descriptor
    7710: romdata_int <= 'hc00;
    7711: romdata_int <= 'h40e;
    7712: romdata_int <= 'hb2d;
    7713: romdata_int <= 'h408; // Line Descriptor
    7714: romdata_int <= 'he00;
    7715: romdata_int <= 'h718;
    7716: romdata_int <= 'h20a;
    7717: romdata_int <= 'h408; // Line Descriptor
    7718: romdata_int <= 'h0;
    7719: romdata_int <= 'ha9b;
    7720: romdata_int <= 'hac5;
    7721: romdata_int <= 'h408; // Line Descriptor
    7722: romdata_int <= 'h200;
    7723: romdata_int <= 'he60;
    7724: romdata_int <= 'h215;
    7725: romdata_int <= 'h408; // Line Descriptor
    7726: romdata_int <= 'h400;
    7727: romdata_int <= 'hd4;
    7728: romdata_int <= 'h8a;
    7729: romdata_int <= 'h408; // Line Descriptor
    7730: romdata_int <= 'h600;
    7731: romdata_int <= 'h4ef;
    7732: romdata_int <= 'hf61;
    7733: romdata_int <= 'h408; // Line Descriptor
    7734: romdata_int <= 'h800;
    7735: romdata_int <= 'h842;
    7736: romdata_int <= 'h4b5;
    7737: romdata_int <= 'h408; // Line Descriptor
    7738: romdata_int <= 'ha00;
    7739: romdata_int <= 'h60b;
    7740: romdata_int <= 'hc79;
    7741: romdata_int <= 'h408; // Line Descriptor
    7742: romdata_int <= 'hc00;
    7743: romdata_int <= 'h23e;
    7744: romdata_int <= 'h916;
    7745: romdata_int <= 'h408; // Line Descriptor
    7746: romdata_int <= 'he00;
    7747: romdata_int <= 'hd22;
    7748: romdata_int <= 'h6c5;
    7749: romdata_int <= 'h408; // Line Descriptor
    7750: romdata_int <= 'h0;
    7751: romdata_int <= 'h536;
    7752: romdata_int <= 'h20;
    7753: romdata_int <= 'h408; // Line Descriptor
    7754: romdata_int <= 'h200;
    7755: romdata_int <= 'ha8b;
    7756: romdata_int <= 'ha9d;
    7757: romdata_int <= 'h408; // Line Descriptor
    7758: romdata_int <= 'h400;
    7759: romdata_int <= 'h29d;
    7760: romdata_int <= 'h4cf;
    7761: romdata_int <= 'h408; // Line Descriptor
    7762: romdata_int <= 'h600;
    7763: romdata_int <= 'hcb8;
    7764: romdata_int <= 'h299;
    7765: romdata_int <= 'h408; // Line Descriptor
    7766: romdata_int <= 'h800;
    7767: romdata_int <= 'hf39;
    7768: romdata_int <= 'h87a;
    7769: romdata_int <= 'h408; // Line Descriptor
    7770: romdata_int <= 'ha00;
    7771: romdata_int <= 'h122;
    7772: romdata_int <= 'h74e;
    7773: romdata_int <= 'h408; // Line Descriptor
    7774: romdata_int <= 'hc00;
    7775: romdata_int <= 'h636;
    7776: romdata_int <= 'hc9f;
    7777: romdata_int <= 'h408; // Line Descriptor
    7778: romdata_int <= 'he00;
    7779: romdata_int <= 'h81c;
    7780: romdata_int <= 'he3e;
    7781: romdata_int <= 'h408; // Line Descriptor
    7782: romdata_int <= 'h0;
    7783: romdata_int <= 'haeb;
    7784: romdata_int <= 'h328;
    7785: romdata_int <= 'h408; // Line Descriptor
    7786: romdata_int <= 'h200;
    7787: romdata_int <= 'h207;
    7788: romdata_int <= 'h63c;
    7789: romdata_int <= 'h408; // Line Descriptor
    7790: romdata_int <= 'h400;
    7791: romdata_int <= 'hc68;
    7792: romdata_int <= 'h483;
    7793: romdata_int <= 'h408; // Line Descriptor
    7794: romdata_int <= 'h600;
    7795: romdata_int <= 'he99;
    7796: romdata_int <= 'hcf8;
    7797: romdata_int <= 'h408; // Line Descriptor
    7798: romdata_int <= 'h800;
    7799: romdata_int <= 'h4d9;
    7800: romdata_int <= 'h808;
    7801: romdata_int <= 'h408; // Line Descriptor
    7802: romdata_int <= 'ha00;
    7803: romdata_int <= 'h12b;
    7804: romdata_int <= 'he76;
    7805: romdata_int <= 'h408; // Line Descriptor
    7806: romdata_int <= 'hc00;
    7807: romdata_int <= 'h614;
    7808: romdata_int <= 'ha50;
    7809: romdata_int <= 'h508; // Line Descriptor
    7810: romdata_int <= 'he00;
    7811: romdata_int <= 'h94a;
    7812: romdata_int <= 'hd5;
    7813: romdata_int <= 'h605; // Line Descriptor
    7814: romdata_int <= 'h0;
    7815: romdata_int <= 'h737;
    7816: romdata_int <= 'h48e;
    7817: romdata_int <= 'ha1;
    7818: romdata_int <= 'h605; // Line Descriptor
    7819: romdata_int <= 'h200;
    7820: romdata_int <= 'h122;
    7821: romdata_int <= 'h6ae;
    7822: romdata_int <= 'h50b;
    7823: romdata_int <= 'h605; // Line Descriptor
    7824: romdata_int <= 'h400;
    7825: romdata_int <= 'h35c;
    7826: romdata_int <= 'h8e1;
    7827: romdata_int <= 'h8ec;
    7828: romdata_int <= 'h605; // Line Descriptor
    7829: romdata_int <= 'h600;
    7830: romdata_int <= 'h83a;
    7831: romdata_int <= 'h2a1;
    7832: romdata_int <= 'h339;
    7833: romdata_int <= 'h605; // Line Descriptor
    7834: romdata_int <= 'h800;
    7835: romdata_int <= 'h460;
    7836: romdata_int <= 'h79;
    7837: romdata_int <= 'h6b8;
    7838: romdata_int <= 'h405; // Line Descriptor
    7839: romdata_int <= 'h0;
    7840: romdata_int <= 'h2b9;
    7841: romdata_int <= 'h73b;
    7842: romdata_int <= 'h405; // Line Descriptor
    7843: romdata_int <= 'h200;
    7844: romdata_int <= 'h49b;
    7845: romdata_int <= 'h912;
    7846: romdata_int <= 'h405; // Line Descriptor
    7847: romdata_int <= 'h400;
    7848: romdata_int <= 'h679;
    7849: romdata_int <= 'h21e;
    7850: romdata_int <= 'h405; // Line Descriptor
    7851: romdata_int <= 'h600;
    7852: romdata_int <= 'hef;
    7853: romdata_int <= 'h2a;
    7854: romdata_int <= 'h405; // Line Descriptor
    7855: romdata_int <= 'h800;
    7856: romdata_int <= 'h928;
    7857: romdata_int <= 'h48a;
    7858: romdata_int <= 'h405; // Line Descriptor
    7859: romdata_int <= 'h0;
    7860: romdata_int <= 'h455;
    7861: romdata_int <= 'h661;
    7862: romdata_int <= 'h405; // Line Descriptor
    7863: romdata_int <= 'h200;
    7864: romdata_int <= 'h6a5;
    7865: romdata_int <= 'h8e0;
    7866: romdata_int <= 'h405; // Line Descriptor
    7867: romdata_int <= 'h400;
    7868: romdata_int <= 'h8ae;
    7869: romdata_int <= 'h311;
    7870: romdata_int <= 'h405; // Line Descriptor
    7871: romdata_int <= 'h600;
    7872: romdata_int <= 'h12c;
    7873: romdata_int <= 'ha7;
    7874: romdata_int <= 'h405; // Line Descriptor
    7875: romdata_int <= 'h800;
    7876: romdata_int <= 'h32b;
    7877: romdata_int <= 'h464;
    7878: romdata_int <= 'h405; // Line Descriptor
    7879: romdata_int <= 'h0;
    7880: romdata_int <= 'h2c9;
    7881: romdata_int <= 'h354;
    7882: romdata_int <= 'h405; // Line Descriptor
    7883: romdata_int <= 'h200;
    7884: romdata_int <= 'he7;
    7885: romdata_int <= 'h413;
    7886: romdata_int <= 'h405; // Line Descriptor
    7887: romdata_int <= 'h400;
    7888: romdata_int <= 'h483;
    7889: romdata_int <= 'h718;
    7890: romdata_int <= 'h405; // Line Descriptor
    7891: romdata_int <= 'h600;
    7892: romdata_int <= 'h722;
    7893: romdata_int <= 'h87c;
    7894: romdata_int <= 'h405; // Line Descriptor
    7895: romdata_int <= 'h800;
    7896: romdata_int <= 'h855;
    7897: romdata_int <= 'h12b;
    7898: romdata_int <= 'h405; // Line Descriptor
    7899: romdata_int <= 'h0;
    7900: romdata_int <= 'h8a1;
    7901: romdata_int <= 'h4d;
    7902: romdata_int <= 'h405; // Line Descriptor
    7903: romdata_int <= 'h200;
    7904: romdata_int <= 'h449;
    7905: romdata_int <= 'h21e;
    7906: romdata_int <= 'h405; // Line Descriptor
    7907: romdata_int <= 'h400;
    7908: romdata_int <= 'h708;
    7909: romdata_int <= 'h428;
    7910: romdata_int <= 'h405; // Line Descriptor
    7911: romdata_int <= 'h600;
    7912: romdata_int <= 'hc0;
    7913: romdata_int <= 'h63f;
    7914: romdata_int <= 'h405; // Line Descriptor
    7915: romdata_int <= 'h800;
    7916: romdata_int <= 'h322;
    7917: romdata_int <= 'h8cf;
    7918: romdata_int <= 'h405; // Line Descriptor
    7919: romdata_int <= 'h0;
    7920: romdata_int <= 'h6db;
    7921: romdata_int <= 'h558;
    7922: romdata_int <= 'h405; // Line Descriptor
    7923: romdata_int <= 'h200;
    7924: romdata_int <= 'hcb;
    7925: romdata_int <= 'h71d;
    7926: romdata_int <= 'h405; // Line Descriptor
    7927: romdata_int <= 'h400;
    7928: romdata_int <= 'h2fc;
    7929: romdata_int <= 'h938;
    7930: romdata_int <= 'h405; // Line Descriptor
    7931: romdata_int <= 'h600;
    7932: romdata_int <= 'h86c;
    7933: romdata_int <= 'hee;
    7934: romdata_int <= 'h405; // Line Descriptor
    7935: romdata_int <= 'h800;
    7936: romdata_int <= 'h526;
    7937: romdata_int <= 'h2f9;
    7938: romdata_int <= 'h405; // Line Descriptor
    7939: romdata_int <= 'h0;
    7940: romdata_int <= 'h665;
    7941: romdata_int <= 'h7e;
    7942: romdata_int <= 'h405; // Line Descriptor
    7943: romdata_int <= 'h200;
    7944: romdata_int <= 'h254;
    7945: romdata_int <= 'h954;
    7946: romdata_int <= 'h405; // Line Descriptor
    7947: romdata_int <= 'h400;
    7948: romdata_int <= 'h838;
    7949: romdata_int <= 'h6b3;
    7950: romdata_int <= 'h405; // Line Descriptor
    7951: romdata_int <= 'h600;
    7952: romdata_int <= 'h44e;
    7953: romdata_int <= 'h473;
    7954: romdata_int <= 'h405; // Line Descriptor
    7955: romdata_int <= 'h800;
    7956: romdata_int <= 'he7;
    7957: romdata_int <= 'h26f;
    7958: romdata_int <= 'h405; // Line Descriptor
    7959: romdata_int <= 'h0;
    7960: romdata_int <= 'h27e;
    7961: romdata_int <= 'hc8;
    7962: romdata_int <= 'h405; // Line Descriptor
    7963: romdata_int <= 'h200;
    7964: romdata_int <= 'h492;
    7965: romdata_int <= 'h711;
    7966: romdata_int <= 'h405; // Line Descriptor
    7967: romdata_int <= 'h400;
    7968: romdata_int <= 'h709;
    7969: romdata_int <= 'h841;
    7970: romdata_int <= 'h405; // Line Descriptor
    7971: romdata_int <= 'h600;
    7972: romdata_int <= 'h12f;
    7973: romdata_int <= 'h265;
    7974: romdata_int <= 'h505; // Line Descriptor
    7975: romdata_int <= 'h800;
    7976: romdata_int <= 'h8dc;
    default: romdata_int <= 'h4ea;
  endcase
endmodule
