library ieee;
use ieee.std_logic_1164.all;
use work.fp24_type_pkg.all;

package fp24_init1_pkg is

constant mem_init1:	bit_array_1024x48:=(
(0)=>    "000000000000000000000000010000000000000000000000",
(1)=>    "001011011001010000000000001111101111111111111110",
(2)=>    "001011111001010000000000001111101111111111111110",
(3)=>    "001100010010111000000000001111101111111111111110",
(4)=>    "001100011001001100000000001111101111111111111100",
(5)=>    "001100011111011100000000001111101111111111111100",
(6)=>    "001100110010111000000000001111101111111111111010",
(7)=>    "001100110110000000000000001111101111111111111000",
(8)=>    "001100111001001010000000001111101111111111110110",
(9)=>    "001100111100010010000000001111101111111111110010",
(10)=>    "001100111111011100000000001111101111111111110000",
(11)=>    "001101010001010010000000001111101111111111101100",
(12)=>    "001101010010110111000000001111101111111111101000",
(13)=>    "001101010100011011000000001111101111111111100100",
(14)=>    "001101010110000000000000001111101111111111100000",
(15)=>    "001101010111100100000000001111101111111111011100",
(16)=>    "001101011001001001000000001111101111111111011000",
(17)=>    "001101011010101101000000001111101111111111010010",
(18)=>    "001101011100010010000000001111101111111111001110",
(19)=>    "001101011101110110000000001111101111111111001000",
(20)=>    "001101011111011011000000001111101111111111000010",
(21)=>    "001101110000011111100000001111101111111110111010",
(22)=>    "001101110001010010000000001111101111111110110100",
(23)=>    "001101110010000100000000001111101111111110101110",
(24)=>    "001101110010110110100000001111101111111110100110",
(25)=>    "001101110011101000100000001111101111111110011110",
(26)=>    "001101110100011011000000001111101111111110010110",
(27)=>    "001101110101001101000000001111101111111110001110",
(28)=>    "001101110101111111100000001111101111111110000110",
(29)=>    "001101110110110001100000001111101111111101111110",
(30)=>    "001101110111100011100000001111101111111101110100",
(31)=>    "001101111000010110000000001111101111111101101010",
(32)=>    "001101111001001000000000001111101111111101100010",
(33)=>    "001101111001111010100000001111101111111101011000",
(34)=>    "001101111010101100100000001111101111111101001100",
(35)=>    "001101111011011110100000001111101111111101000010",
(36)=>    "001101111100010001000000001111101111111100111000",
(37)=>    "001101111101000011000000001111101111111100101100",
(38)=>    "001101111101110101100000001111101111111100100000",
(39)=>    "001101111110100111100000001111101111111100010100",
(40)=>    "001101111111011001100000001111101111111100001000",
(41)=>    "001110010000000110000000001111101111111011111100",
(42)=>    "001110010000011111000000001111101111111011110000",
(43)=>    "001110010000111000000000001111101111111011100010",
(44)=>    "001110010001010001010000001111101111111011010100",
(45)=>    "001110010001101010010000001111101111111011000110",
(46)=>    "001110010010000011010000001111101111111010111000",
(47)=>    "001110010010011100010000001111101111111010101010",
(48)=>    "001110010010110101100000001111101111111010011100",
(49)=>    "001110010011001110100000001111101111111010001100",
(50)=>    "001110010011100111100000001111101111111001111110",
(51)=>    "001110010100000000100000001111101111111001101110",
(52)=>    "001110010100011001110000001111101111111001011110",
(53)=>    "001110010100110010110000001111101111111001001110",
(54)=>    "001110010101001011110000001111101111111000111110",
(55)=>    "001110010101100100110000001111101111111000101100",
(56)=>    "001110010101111101110000001111101111111000011100",
(57)=>    "001110010110010110110000001111101111111000001010",
(58)=>    "001110010110110000000000001111101111110111111000",
(59)=>    "001110010111001001000000001111101111110111100110",
(60)=>    "001110010111100010000000001111101111110111010100",
(61)=>    "001110010111111011000000001111101111110111000010",
(62)=>    "001110011000010100000000001111101111110110101110",
(63)=>    "001110011000101101000000001111101111110110011100",
(64)=>    "001110011001000110000000001111101111110110001000",
(65)=>    "001110011001011111000000001111101111110101110100",
(66)=>    "001110011001111000000000001111101111110101100000",
(67)=>    "001110011010010001000000001111101111110101001100",
(68)=>    "001110011010101010000000001111101111110100110110",
(69)=>    "001110011011000011000000001111101111110100100010",
(70)=>    "001110011011011100000000001111101111110100001100",
(71)=>    "001110011011110101000000001111101111110011110110",
(72)=>    "001110011100001110000000001111101111110011100000",
(73)=>    "001110011100100111000000001111101111110011001010",
(74)=>    "001110011101000000000000001111101111110010110100",
(75)=>    "001110011101011001000000001111101111110010011100",
(76)=>    "001110011101110010000000001111101111110010000110",
(77)=>    "001110011110001010110000001111101111110001101110",
(78)=>    "001110011110100011110000001111101111110001010110",
(79)=>    "001110011110111100110000001111101111110000111110",
(80)=>    "001110011111010101110000001111101111110000100110",
(81)=>    "001110011111101110110000001111101111110000001100",
(82)=>    "001110110000000011110000001111101111101111110100",
(83)=>    "001110110000010000010000001111101111101111011010",
(84)=>    "001110110000011100110000001111101111101111000000",
(85)=>    "001110110000101001001000001111101111101110100110",
(86)=>    "001110110000110101101000001111101111101110001100",
(87)=>    "001110110001000010001000001111101111101101110010",
(88)=>    "001110110001001110100000001111101111101101010110",
(89)=>    "001110110001011011000000001111101111101100111100",
(90)=>    "001110110001100111100000001111101111101100100000",
(91)=>    "001110110001110011111000001111101111101100000100",
(92)=>    "001110110010000000011000001111101111101011101000",
(93)=>    "001110110010001100110000001111101111101011001100",
(94)=>    "001110110010011001010000001111101111101010101110",
(95)=>    "001110110010100101101000001111101111101010010010",
(96)=>    "001110110010110010001000001111101111101001110100",
(97)=>    "001110110010111110100000001111101111101001010110",
(98)=>    "001110110011001010111000001111101111101000111000",
(99)=>    "001110110011010111011000001111101111101000011010",
(100)=>    "001110110011100011110000001111101111100111111100",
(101)=>    "001110110011110000010000001111101111100111011110",
(102)=>    "001110110011111100101000001111101111100110111110",
(103)=>    "001110110100001001000000001111101111100110011110",
(104)=>    "001110110100010101011000001111101111100101111110",
(105)=>    "001110110100100001111000001111101111100101011110",
(106)=>    "001110110100101110010000001111101111100100111110",
(107)=>    "001110110100111010101000001111101111100100011110",
(108)=>    "001110110101000111000000001111101111100011111100",
(109)=>    "001110110101010011011000001111101111100011011100",
(110)=>    "001110110101011111111000001111101111100010111010",
(111)=>    "001110110101101100010000001111101111100010011000",
(112)=>    "001110110101111000101000001111101111100001110110",
(113)=>    "001110110110000101000000001111101111100001010010",
(114)=>    "001110110110010001011000001111101111100000110000",
(115)=>    "001110110110011101110000001111101111100000001100",
(116)=>    "001110110110101010001000001111101111011111101010",
(117)=>    "001110110110110110100000001111101111011111000110",
(118)=>    "001110110111000010110000001111101111011110100010",
(119)=>    "001110110111001111001000001111101111011101111110",
(120)=>    "001110110111011011100000001111101111011101011000",
(121)=>    "001110110111100111111000001111101111011100110100",
(122)=>    "001110110111110100010000001111101111011100001110",
(123)=>    "001110111000000000101000001111101111011011101000",
(124)=>    "001110111000001100111000001111101111011011000010",
(125)=>    "001110111000011001010000001111101111011010011100",
(126)=>    "001110111000100101101000001111101111011001110110",
(127)=>    "001110111000110001111000001111101111011001010000",
(128)=>    "001110111000111110010000001111101111011000101000",
(129)=>    "001110111001001010101000001111101111011000000010",
(130)=>    "001110111001010110111000001111101111010111011010",
(131)=>    "001110111001100011010000001111101111010110110010",
(132)=>    "001110111001101111100000001111101111010110001010",
(133)=>    "001110111001111011111000001111101111010101100000",
(134)=>    "001110111010001000001000001111101111010100111000",
(135)=>    "001110111010010100011000001111101111010100001110",
(136)=>    "001110111010100000110000001111101111010011100110",
(137)=>    "001110111010101101000000001111101111010010111100",
(138)=>    "001110111010111001010000001111101111010010010010",
(139)=>    "001110111011000101101000001111101111010001100110",
(140)=>    "001110111011010001111000001111101111010000111100",
(141)=>    "001110111011011110001000001111101111010000010010",
(142)=>    "001110111011101010011000001111101111001111100110",
(143)=>    "001110111011110110101000001111101111001110111010",
(144)=>    "001110111100000011000000001111101111001110001110",
(145)=>    "001110111100001111010000001111101111001101100010",
(146)=>    "001110111100011011100000001111101111001100110110",
(147)=>    "001110111100100111110000001111101111001100001000",
(148)=>    "001110111100110100000000001111101111001011011100",
(149)=>    "001110111101000000010000001111101111001010101110",
(150)=>    "001110111101001100011000001111101111001010000000",
(151)=>    "001110111101011000101000001111101111001001010010",
(152)=>    "001110111101100100111000001111101111001000100100",
(153)=>    "001110111101110001001000001111101111000111110110",
(154)=>    "001110111101111101011000001111101111000111000110",
(155)=>    "001110111110001001100000001111101111000110011000",
(156)=>    "001110111110010101110000001111101111000101101000",
(157)=>    "001110111110100010000000001111101111000100111000",
(158)=>    "001110111110101110001000001111101111000100001000",
(159)=>    "001110111110111010011000001111101111000011011000",
(160)=>    "001110111111000110100000001111101111000010100110",
(161)=>    "001110111111010010110000001111101111000001110110",
(162)=>    "001110111111011110111000001111101111000001000100",
(163)=>    "001110111111101011001000001111101111000000010100",
(164)=>    "001110111111110111010000001111101110111111100010",
(165)=>    "001111010000000001110000001111101110111110101110",
(166)=>    "001111010000000111110100001111101110111101111100",
(167)=>    "001111010000001101111000001111101110111101001010",
(168)=>    "001111010000010011111100001111101110111100010110",
(169)=>    "001111010000011010000100001111101110111011100100",
(170)=>    "001111010000100000001000001111101110111010110000",
(171)=>    "001111010000100110001100001111101110111001111100",
(172)=>    "001111010000101100010000001111101110111001001000",
(173)=>    "001111010000110010010100001111101110111000010010",
(174)=>    "001111010000111000011000001111101110110111011110",
(175)=>    "001111010000111110011100001111101110110110101000",
(176)=>    "001111010001000100100000001111101110110101110100",
(177)=>    "001111010001001010100100001111101110110100111110",
(178)=>    "001111010001010000100100001111101110110100001000",
(179)=>    "001111010001010110101000001111101110110011010000",
(180)=>    "001111010001011100101100001111101110110010011010",
(181)=>    "001111010001100010110000001111101110110001100100",
(182)=>    "001111010001101000110000001111101110110000101100",
(183)=>    "001111010001101110110100001111101110101111110100",
(184)=>    "001111010001110100111000001111101110101110111100",
(185)=>    "001111010001111010111000001111101110101110000100",
(186)=>    "001111010010000000111100001111101110101101001100",
(187)=>    "001111010010000110111100001111101110101100010100",
(188)=>    "001111010010001100111100001111101110101011011010",
(189)=>    "001111010010010011000000001111101110101010100000",
(190)=>    "001111010010011001000000001111101110101001101000",
(191)=>    "001111010010011111000000001111101110101000101110",
(192)=>    "001111010010100101000100001111101110100111110100",
(193)=>    "001111010010101011000100001111101110100110111000",
(194)=>    "001111010010110001000100001111101110100101111110",
(195)=>    "001111010010110111000100001111101110100101000010",
(196)=>    "001111010010111101000100001111101110100100001000",
(197)=>    "001111010011000011000100001111101110100011001100",
(198)=>    "001111010011001001000100001111101110100010010000",
(199)=>    "001111010011001111000100001111101110100001010100",
(200)=>    "001111010011010101000100001111101110100000010110",
(201)=>    "001111010011011011000100001111101110011111011010",
(202)=>    "001111010011100001000000001111101110011110011100",
(203)=>    "001111010011100111000000001111101110011101100000",
(204)=>    "001111010011101101000000001111101110011100100010",
(205)=>    "001111010011110010111100001111101110011011100100",
(206)=>    "001111010011111000111100001111101110011010100110",
(207)=>    "001111010011111110111000001111101110011001100110",
(208)=>    "001111010100000100111000001111101110011000101000",
(209)=>    "001111010100001010110100001111101110010111101000",
(210)=>    "001111010100010000110100001111101110010110101000",
(211)=>    "001111010100010110110000001111101110010101101010",
(212)=>    "001111010100011100101100001111101110010100101000",
(213)=>    "001111010100100010101100001111101110010011101000",
(214)=>    "001111010100101000101000001111101110010010101000",
(215)=>    "001111010100101110100100001111101110010001100110",
(216)=>    "001111010100110100100000001111101110010000100110",
(217)=>    "001111010100111010011100001111101110001111100100",
(218)=>    "001111010101000000011000001111101110001110100010",
(219)=>    "001111010101000110010100001111101110001101100000",
(220)=>    "001111010101001100010000001111101110001100011110",
(221)=>    "001111010101010010001100001111101110001011011010",
(222)=>    "001111010101011000001000001111101110001010011000",
(223)=>    "001111010101011110000000001111101110001001010100",
(224)=>    "001111010101100011111100001111101110001000010010",
(225)=>    "001111010101101001111000001111101110000111001110",
(226)=>    "001111010101101111110000001111101110000110001010",
(227)=>    "001111010101110101101100001111101110000101000100",
(228)=>    "001111010101111011100100001111101110000100000000",
(229)=>    "001111010110000001100000001111101110000010111010",
(230)=>    "001111010110000111011000001111101110000001110110",
(231)=>    "001111010110001101010000001111101110000000110000",
(232)=>    "001111010110010011001000001111101101111111101010",
(233)=>    "001111010110011001000100001111101101111110100100",
(234)=>    "001111010110011110111100001111101101111101011110",
(235)=>    "001111010110100100110100001111101101111100010110",
(236)=>    "001111010110101010101100001111101101111011010000",
(237)=>    "001111010110110000100100001111101101111010001000",
(238)=>    "001111010110110110011100001111101101111001000000",
(239)=>    "001111010110111100010100001111101101110111111000",
(240)=>    "001111010111000010001100001111101101110110110000",
(241)=>    "001111010111001000000000001111101101110101101000",
(242)=>    "001111010111001101111000001111101101110100011110",
(243)=>    "001111010111010011110000001111101101110011010110",
(244)=>    "001111010111011001100100001111101101110010001100",
(245)=>    "001111010111011111011100001111101101110001000010",
(246)=>    "001111010111100101010000001111101101101111111000",
(247)=>    "001111010111101011001000001111101101101110101110",
(248)=>    "001111010111110000111100001111101101101101100100",
(249)=>    "001111010111110110110000001111101101101100011010",
(250)=>    "001111010111111100101000001111101101101011001110",
(251)=>    "001111011000000010011100001111101101101010000010",
(252)=>    "001111011000001000010000001111101101101000111000",
(253)=>    "001111011000001110000100001111101101100111101100",
(254)=>    "001111011000010011111000001111101101100110100000",
(255)=>    "001111011000011001101100001111101101100101010010",
(256)=>    "001111011000011111100000001111101101100100000110",
(257)=>    "001111011000100101010100001111101101100010111000",
(258)=>    "001111011000101011001000001111101101100001101100",
(259)=>    "001111011000110000111000001111101101100000011110",
(260)=>    "001111011000110110101100001111101101011111010000",
(261)=>    "001111011000111100100000001111101101011110000010",
(262)=>    "001111011001000010010000001111101101011100110010",
(263)=>    "001111011001001000000100001111101101011011100100",
(264)=>    "001111011001001101110100001111101101011010010110",
(265)=>    "001111011001010011101000001111101101011001000110",
(266)=>    "001111011001011001011000001111101101010111110110",
(267)=>    "001111011001011111001000001111101101010110100110",
(268)=>    "001111011001100100111000001111101101010101010110",
(269)=>    "001111011001101010101000001111101101010100000110",
(270)=>    "001111011001110000011000001111101101010010110100",
(271)=>    "001111011001110110001000001111101101010001100100",
(272)=>    "001111011001111011111000001111101101010000010010",
(273)=>    "001111011010000001101000001111101101001111000000",
(274)=>    "001111011010000111011000001111101101001101101110",
(275)=>    "001111011010001101001000001111101101001100011100",
(276)=>    "001111011010010010111000001111101101001011001010",
(277)=>    "001111011010011000100100001111101101001001111000",
(278)=>    "001111011010011110010100001111101101001000100100",
(279)=>    "001111011010100100000000001111101101000111010010",
(280)=>    "001111011010101001110000001111101101000101111110",
(281)=>    "001111011010101111011100001111101101000100101010",
(282)=>    "001111011010110101001000001111101101000011010110",
(283)=>    "001111011010111010111000001111101101000010000010",
(284)=>    "001111011011000000100100001111101101000000101100",
(285)=>    "001111011011000110010000001111101100111111011000",
(286)=>    "001111011011001011111100001111101100111110000010",
(287)=>    "001111011011010001101000001111101100111100101100",
(288)=>    "001111011011010111010100001111101100111011010110",
(289)=>    "001111011011011101000000001111101100111010000000",
(290)=>    "001111011011100010101000001111101100111000101010",
(291)=>    "001111011011101000010100001111101100110111010100",
(292)=>    "001111011011101110000000001111101100110101111100",
(293)=>    "001111011011110011101000001111101100110100100110",
(294)=>    "001111011011111001010100001111101100110011001110",
(295)=>    "001111011011111110111100001111101100110001110110",
(296)=>    "001111011100000100101000001111101100110000011110",
(297)=>    "001111011100001010010000001111101100101111000110",
(298)=>    "001111011100001111111000001111101100101101101110",
(299)=>    "001111011100010101100000001111101100101100010100",
(300)=>    "001111011100011011001000001111101100101010111100",
(301)=>    "001111011100100000110100001111101100101001100010",
(302)=>    "001111011100100110011000001111101100101000001000",
(303)=>    "001111011100101100000000001111101100100110101110",
(304)=>    "001111011100110001101000001111101100100101010100",
(305)=>    "001111011100110111010000001111101100100011111010",
(306)=>    "001111011100111100111000001111101100100010011110",
(307)=>    "001111011101000010011100001111101100100001000100",
(308)=>    "001111011101001000000100001111101100011111101000",
(309)=>    "001111011101001101101000001111101100011110001100",
(310)=>    "001111011101010011010000001111101100011100110000",
(311)=>    "001111011101011000110100001111101100011011010100",
(312)=>    "001111011101011110011000001111101100011001111000",
(313)=>    "001111011101100100000000001111101100011000011010",
(314)=>    "001111011101101001100100001111101100010110111110",
(315)=>    "001111011101101111001000001111101100010101100000",
(316)=>    "001111011101110100101100001111101100010100000100",
(317)=>    "001111011101111010010000001111101100010010100110",
(318)=>    "001111011101111111110000001111101100010001001000",
(319)=>    "001111011110000101010100001111101100001111101000",
(320)=>    "001111011110001010111000001111101100001110001010",
(321)=>    "001111011110010000011100001111101100001100101100",
(322)=>    "001111011110010101111100001111101100001011001100",
(323)=>    "001111011110011011100000001111101100001001101100",
(324)=>    "001111011110100001000000001111101100001000001100",
(325)=>    "001111011110100110100000001111101100000110101100",
(326)=>    "001111011110101100000100001111101100000101001100",
(327)=>    "001111011110110001100100001111101100000011101100",
(328)=>    "001111011110110111000100001111101100000010001100",
(329)=>    "001111011110111100100100001111101100000000101010",
(330)=>    "001111011111000010000100001111101011111111001000",
(331)=>    "001111011111000111100100001111101011111101101000",
(332)=>    "001111011111001101000100001111101011111100000110",
(333)=>    "001111011111010010100000001111101011111010100100",
(334)=>    "001111011111011000000000001111101011111001000000",
(335)=>    "001111011111011101100000001111101011110111011110",
(336)=>    "001111011111100010111100001111101011110101111100",
(337)=>    "001111011111101000011100001111101011110100011000",
(338)=>    "001111011111101101111000001111101011110010110100",
(339)=>    "001111011111110011010100001111101011110001010000",
(340)=>    "001111011111111000110000001111101011101111101100",
(341)=>    "001111011111111110001100001111101011101110001000",
(342)=>    "001111110000000001110110001111101011101100100100",
(343)=>    "001111110000000100100010001111101011101010111110",
(344)=>    "001111110000000111010000001111101011101001011010",
(345)=>    "001111110000001001111110001111101011100111110100",
(346)=>    "001111110000001100101100001111101011100110001110",
(347)=>    "001111110000001111011010001111101011100100101000",
(348)=>    "001111110000010010000110001111101011100011000010",
(349)=>    "001111110000010100110100001111101011100001011100",
(350)=>    "001111110000010111100000001111101011011111110110",
(351)=>    "001111110000011010001100001111101011011110001110",
(352)=>    "001111110000011100111010001111101011011100101000",
(353)=>    "001111110000011111100110001111101011011011000000",
(354)=>    "001111110000100010010010001111101011011001011000",
(355)=>    "001111110000100100111110001111101011010111110000",
(356)=>    "001111110000100111101010001111101011010110001000",
(357)=>    "001111110000101010010110001111101011010100100000",
(358)=>    "001111110000101101000010001111101011010010110110",
(359)=>    "001111110000101111101100001111101011010001001110",
(360)=>    "001111110000110010011000001111101011001111100100",
(361)=>    "001111110000110101000100001111101011001101111010",
(362)=>    "001111110000110111101110001111101011001100010000",
(363)=>    "001111110000111010011000001111101011001010100110",
(364)=>    "001111110000111101000100001111101011001000111100",
(365)=>    "001111110000111111101110001111101011000111010010",
(366)=>    "001111110001000010011000001111101011000101100110",
(367)=>    "001111110001000101000010001111101011000011111100",
(368)=>    "001111110001000111101100001111101011000010010000",
(369)=>    "001111110001001010010110001111101011000000100100",
(370)=>    "001111110001001101000000001111101010111110111000",
(371)=>    "001111110001001111101010001111101010111101001100",
(372)=>    "001111110001010010010010001111101010111011100000",
(373)=>    "001111110001010100111100001111101010111001110010",
(374)=>    "001111110001010111100100001111101010111000000110",
(375)=>    "001111110001011010001110001111101010110110011000",
(376)=>    "001111110001011100110110001111101010110100101010",
(377)=>    "001111110001011111011110001111101010110010111110",
(378)=>    "001111110001100010000110001111101010110001001110",
(379)=>    "001111110001100100101110001111101010101111100000",
(380)=>    "001111110001100111010110001111101010101101110010",
(381)=>    "001111110001101001111110001111101010101100000100",
(382)=>    "001111110001101100100110001111101010101010010100",
(383)=>    "001111110001101111001110001111101010101000100100",
(384)=>    "001111110001110001110100001111101010100110110110",
(385)=>    "001111110001110100011100001111101010100101000110",
(386)=>    "001111110001110111000010001111101010100011010110",
(387)=>    "001111110001111001101010001111101010100001100110",
(388)=>    "001111110001111100010000001111101010011111110100",
(389)=>    "001111110001111110110110001111101010011110000100",
(390)=>    "001111110010000001011100001111101010011100010010",
(391)=>    "001111110010000100000010001111101010011010100010",
(392)=>    "001111110010000110101000001111101010011000110000",
(393)=>    "001111110010001001001110001111101010010110111110",
(394)=>    "001111110010001011110100001111101010010101001100",
(395)=>    "001111110010001110011010001111101010010011011010",
(396)=>    "001111110010010000111110001111101010010001100110",
(397)=>    "001111110010010011100100001111101010001111110100",
(398)=>    "001111110010010110001000001111101010001110000000",
(399)=>    "001111110010011000101100001111101010001100001110",
(400)=>    "001111110010011011010010001111101010001010011010",
(401)=>    "001111110010011101110110001111101010001000100110",
(402)=>    "001111110010100000011010001111101010000110110010",
(403)=>    "001111110010100010111110001111101010000100111110",
(404)=>    "001111110010100101100010001111101010000011001000",
(405)=>    "001111110010101000000110001111101010000001010100",
(406)=>    "001111110010101010101000001111101001111111011110",
(407)=>    "001111110010101101001100001111101001111101101000",
(408)=>    "001111110010101111101110001111101001111011110100",
(409)=>    "001111110010110010010010001111101001111001111110",
(410)=>    "001111110010110100110100001111101001111000001000",
(411)=>    "001111110010110111010110001111101001110110010000",
(412)=>    "001111110010111001111010001111101001110100011010",
(413)=>    "001111110010111100011100001111101001110010100100",
(414)=>    "001111110010111110111110001111101001110000101100",
(415)=>    "001111110011000001011110001111101001101110110100",
(416)=>    "001111110011000100000000001111101001101100111110",
(417)=>    "001111110011000110100010001111101001101011000110",
(418)=>    "001111110011001001000100001111101001101001001100",
(419)=>    "001111110011001011100100001111101001100111010100",
(420)=>    "001111110011001110000110001111101001100101011100",
(421)=>    "001111110011010000100110001111101001100011100100",
(422)=>    "001111110011010011000110001111101001100001101010",
(423)=>    "001111110011010101100110001111101001011111110000",
(424)=>    "001111110011011000000110001111101001011101110110",
(425)=>    "001111110011011010100110001111101001011011111110",
(426)=>    "001111110011011101000110001111101001011010000010",
(427)=>    "001111110011011111100110001111101001011000001000",
(428)=>    "001111110011100010000110001111101001010110001110",
(429)=>    "001111110011100100100100001111101001010100010100",
(430)=>    "001111110011100111000100001111101001010010011000",
(431)=>    "001111110011101001100010001111101001010000011100",
(432)=>    "001111110011101100000000001111101001001110100010",
(433)=>    "001111110011101110100000001111101001001100100110",
(434)=>    "001111110011110000111110001111101001001010101010",
(435)=>    "001111110011110011011100001111101001001000101100",
(436)=>    "001111110011110101111010001111101001000110110000",
(437)=>    "001111110011111000010110001111101001000100110100",
(438)=>    "001111110011111010110100001111101001000010110110",
(439)=>    "001111110011111101010010001111101001000000111010",
(440)=>    "001111110011111111101110001111101000111110111100",
(441)=>    "001111110100000010001100001111101000111100111110",
(442)=>    "001111110100000100101000001111101000111011000000",
(443)=>    "001111110100000111000100001111101000111001000010",
(444)=>    "001111110100001001100000001111101000110111000100",
(445)=>    "001111110100001011111110001111101000110101000100",
(446)=>    "001111110100001110011000001111101000110011000110",
(447)=>    "001111110100010000110100001111101000110001000110",
(448)=>    "001111110100010011010000001111101000101111001000",
(449)=>    "001111110100010101101100001111101000101101001000",
(450)=>    "001111110100011000000110001111101000101011001000",
(451)=>    "001111110100011010100010001111101000101001001000",
(452)=>    "001111110100011100111100001111101000100111000110",
(453)=>    "001111110100011111010110001111101000100101000110",
(454)=>    "001111110100100001110010001111101000100011000110",
(455)=>    "001111110100100100001100001111101000100001000100",
(456)=>    "001111110100100110100110001111101000011111000100",
(457)=>    "001111110100101001000000001111101000011101000010",
(458)=>    "001111110100101011011000001111101000011011000000",
(459)=>    "001111110100101101110010001111101000011000111110",
(460)=>    "001111110100110000001100001111101000010110111100",
(461)=>    "001111110100110010100100001111101000010100111000",
(462)=>    "001111110100110100111100001111101000010010110110",
(463)=>    "001111110100110111010110001111101000010000110100",
(464)=>    "001111110100111001101110001111101000001110110000",
(465)=>    "001111110100111100000110001111101000001100101100",
(466)=>    "001111110100111110011110001111101000001010101000",
(467)=>    "001111110101000000110110001111101000001000100100",
(468)=>    "001111110101000011001110001111101000000110100000",
(469)=>    "001111110101000101100100001111101000000100011100",
(470)=>    "001111110101000111111100001111101000000010011000",
(471)=>    "001111110101001010010010001111101000000000010010",
(472)=>    "001111110101001100101010001111100111111110001110",
(473)=>    "001111110101001111000000001111100111111100001000",
(474)=>    "001111110101010001010110001111100111111010000010",
(475)=>    "001111110101010011101100001111100111110111111110",
(476)=>    "001111110101010110000010001111100111110101111000",
(477)=>    "001111110101011000011000001111100111110011110000",
(478)=>    "001111110101011010101110001111100111110001101010",
(479)=>    "001111110101011101000010001111100111101111100100",
(480)=>    "001111110101011111011000001111100111101101011100",
(481)=>    "001111110101100001101100001111100111101011010110",
(482)=>    "001111110101100100000010001111100111101001001110",
(483)=>    "001111110101100110010110001111100111100111000110",
(484)=>    "001111110101101000101010001111100111100101000000",
(485)=>    "001111110101101010111110001111100111100010110110",
(486)=>    "001111110101101101010010001111100111100000101110",
(487)=>    "001111110101101111100110001111100111011110100110",
(488)=>    "001111110101110001111000001111100111011100011110",
(489)=>    "001111110101110100001100001111100111011010010100",
(490)=>    "001111110101110110011110001111100111011000001100",
(491)=>    "001111110101111000110010001111100111010110000010",
(492)=>    "001111110101111011000100001111100111010011111000",
(493)=>    "001111110101111101010110001111100111010001101110",
(494)=>    "001111110101111111101000001111100111001111100100",
(495)=>    "001111110110000001111010001111100111001101011010",
(496)=>    "001111110110000100001100001111100111001011010000",
(497)=>    "001111110110000110011110001111100111001001000100",
(498)=>    "001111110110001000110000001111100111000110111010",
(499)=>    "001111110110001011000000001111100111000100101110",
(500)=>    "001111110110001101010010001111100111000010100100",
(501)=>    "001111110110001111100010001111100111000000011000",
(502)=>    "001111110110010001110010001111100110111110001100",
(503)=>    "001111110110010100000010001111100110111100000000",
(504)=>    "001111110110010110010010001111100110111001110100",
(505)=>    "001111110110011000100010001111100110110111100110",
(506)=>    "001111110110011010110010001111100110110101011010",
(507)=>    "001111110110011101000010001111100110110011001110",
(508)=>    "001111110110011111010000001111100110110001000000",
(509)=>    "001111110110100001100000001111100110101110110010",
(510)=>    "001111110110100011101110001111100110101100100100",
(511)=>    "001111110110100101111100001111100110101010010110",
(512)=>    "001111110110101000001010001111100110101000001000",
(513)=>    "001111110110101010011000001111100110100101111010",
(514)=>    "001111110110101100100110001111100110100011101100",
(515)=>    "001111110110101110110100001111100110100001011110",
(516)=>    "001111110110110001000010001111100110011111001110",
(517)=>    "001111110110110011010000001111100110011101000000",
(518)=>    "001111110110110101011100001111100110011010110000",
(519)=>    "001111110110110111101000001111100110011000100000",
(520)=>    "001111110110111001110110001111100110010110010000",
(521)=>    "001111110110111100000010001111100110010100000000",
(522)=>    "001111110110111110001110001111100110010001110000",
(523)=>    "001111110111000000011010001111100110001111100000",
(524)=>    "001111110111000010100110001111100110001101010000",
(525)=>    "001111110111000100110000001111100110001010111110",
(526)=>    "001111110111000110111100001111100110001000101110",
(527)=>    "001111110111001001000110001111100110000110011100",
(528)=>    "001111110111001011010010001111100110000100001010",
(529)=>    "001111110111001101011100001111100110000001111000",
(530)=>    "001111110111001111100110001111100101111111100110",
(531)=>    "001111110111010001110000001111100101111101010100",
(532)=>    "001111110111010011111010001111100101111011000010",
(533)=>    "001111110111010110000100001111100101111000110000",
(534)=>    "001111110111011000001110001111100101110110011100",
(535)=>    "001111110111011010010110001111100101110100001010",
(536)=>    "001111110111011100100000001111100101110001110110",
(537)=>    "001111110111011110101000001111100101101111100100",
(538)=>    "001111110111100000110000001111100101101101010000",
(539)=>    "001111110111100010111000001111100101101010111100",
(540)=>    "001111110111100101000010001111100101101000101000",
(541)=>    "001111110111100111001000001111100101100110010100",
(542)=>    "001111110111101001010000001111100101100100000000",
(543)=>    "001111110111101011011000001111100101100001101010",
(544)=>    "001111110111101101011110001111100101011111010110",
(545)=>    "001111110111101111100110001111100101011101000000",
(546)=>    "001111110111110001101100001111100101011010101100",
(547)=>    "001111110111110011110010001111100101011000010110",
(548)=>    "001111110111110101111010001111100101010110000000",
(549)=>    "001111110111111000000000001111100101010011101010",
(550)=>    "001111110111111010000100001111100101010001010100",
(551)=>    "001111110111111100001010001111100101001110111110",
(552)=>    "001111110111111110010000001111100101001100101000",
(553)=>    "001111111000000000010100001111100101001010010000",
(554)=>    "001111111000000010011010001111100101000111111010",
(555)=>    "001111111000000100011110001111100101000101100010",
(556)=>    "001111111000000110100010001111100101000011001100",
(557)=>    "001111111000001000100110001111100101000000110100",
(558)=>    "001111111000001010101010001111100100111110011100",
(559)=>    "001111111000001100101110001111100100111100000100",
(560)=>    "001111111000001110110010001111100100111001101100",
(561)=>    "001111111000010000110110001111100100110111010100",
(562)=>    "001111111000010010111000001111100100110100111010",
(563)=>    "001111111000010100111010001111100100110010100010",
(564)=>    "001111111000010110111110001111100100110000001010",
(565)=>    "001111111000011001000000001111100100101101110000",
(566)=>    "001111111000011011000010001111100100101011010110",
(567)=>    "001111111000011101000100001111100100101000111110",
(568)=>    "001111111000011111000110001111100100100110100100",
(569)=>    "001111111000100001000110001111100100100100001010",
(570)=>    "001111111000100011001000001111100100100001110000",
(571)=>    "001111111000100101001000001111100100011111010100",
(572)=>    "001111111000100111001000001111100100011100111010",
(573)=>    "001111111000101001001010001111100100011010100000",
(574)=>    "001111111000101011001010001111100100011000000100",
(575)=>    "001111111000101101001010001111100100010101101010",
(576)=>    "001111111000101111001010001111100100010011001110",
(577)=>    "001111111000110001001000001111100100010000110010",
(578)=>    "001111111000110011001000001111100100001110010110",
(579)=>    "001111111000110101000110001111100100001011111100",
(580)=>    "001111111000110111000110001111100100001001011110",
(581)=>    "001111111000111001000100001111100100000111000010",
(582)=>    "001111111000111011000010001111100100000100100110",
(583)=>    "001111111000111101000000001111100100000010001010",
(584)=>    "001111111000111110111110001111100011111111101100",
(585)=>    "001111111001000000111100001111100011111101010000",
(586)=>    "001111111001000010111000001111100011111010110010",
(587)=>    "001111111001000100110110001111100011111000010100",
(588)=>    "001111111001000110110010001111100011110101111000",
(589)=>    "001111111001001000101110001111100011110011011010",
(590)=>    "001111111001001010101100001111100011110000111100",
(591)=>    "001111111001001100101000001111100011101110011110",
(592)=>    "001111111001001110100100001111100011101011111110",
(593)=>    "001111111001010000011110001111100011101001100000",
(594)=>    "001111111001010010011010001111100011100111000010",
(595)=>    "001111111001010100010110001111100011100100100010",
(596)=>    "001111111001010110010000001111100011100010000100",
(597)=>    "001111111001011000001010001111100011011111100100",
(598)=>    "001111111001011010000100001111100011011101000100",
(599)=>    "001111111001011100000000001111100011011010100100",
(600)=>    "001111111001011101111000001111100011011000000100",
(601)=>    "001111111001011111110010001111100011010101100100",
(602)=>    "001111111001100001101100001111100011010011000100",
(603)=>    "001111111001100011100110001111100011010000100100",
(604)=>    "001111111001100101011110001111100011001110000100",
(605)=>    "001111111001100111010110001111100011001011100010",
(606)=>    "001111111001101001001110001111100011001001000010",
(607)=>    "001111111001101011001000001111100011000110100000",
(608)=>    "001111111001101101000000001111100011000011111110",
(609)=>    "001111111001101110110110001111100011000001011100",
(610)=>    "001111111001110000101110001111100010111110111100",
(611)=>    "001111111001110010100110001111100010111100011010",
(612)=>    "001111111001110100011100001111100010111001111000",
(613)=>    "001111111001110110010010001111100010110111010100",
(614)=>    "001111111001111000001010001111100010110100110010",
(615)=>    "001111111001111010000000001111100010110010010000",
(616)=>    "001111111001111011110110001111100010101111101100",
(617)=>    "001111111001111101101010001111100010101101001010",
(618)=>    "001111111001111111100000001111100010101010100110",
(619)=>    "001111111010000001010110001111100010101000000100",
(620)=>    "001111111010000011001010001111100010100101100000",
(621)=>    "001111111010000101000000001111100010100010111100",
(622)=>    "001111111010000110110100001111100010100000011000",
(623)=>    "001111111010001000101000001111100010011101110100",
(624)=>    "001111111010001010011100001111100010011011010000",
(625)=>    "001111111010001100010000001111100010011000101010",
(626)=>    "001111111010001110000010001111100010010110000110",
(627)=>    "001111111010001111110110001111100010010011100010",
(628)=>    "001111111010010001101000001111100010010000111100",
(629)=>    "001111111010010011011100001111100010001110011000",
(630)=>    "001111111010010101001110001111100010001011110010",
(631)=>    "001111111010010111000000001111100010001001001100",
(632)=>    "001111111010011000110010001111100010000110100110",
(633)=>    "001111111010011010100100001111100010000100000000",
(634)=>    "001111111010011100010100001111100010000001011010",
(635)=>    "001111111010011110000110001111100001111110110100",
(636)=>    "001111111010011111110110001111100001111100001110",
(637)=>    "001111111010100001101000001111100001111001101000",
(638)=>    "001111111010100011011000001111100001110111000000",
(639)=>    "001111111010100101001000001111100001110100011010",
(640)=>    "001111111010100110111000001111100001110001110010",
(641)=>    "001111111010101000100110001111100001101111001100",
(642)=>    "001111111010101010010110001111100001101100100100",
(643)=>    "001111111010101100000110001111100001101001111100",
(644)=>    "001111111010101101110100001111100001100111010100",
(645)=>    "001111111010101111100010001111100001100100101100",
(646)=>    "001111111010110001010000001111100001100010000100",
(647)=>    "001111111010110011000000001111100001011111011100",
(648)=>    "001111111010110100101100001111100001011100110100",
(649)=>    "001111111010110110011010001111100001011010001100",
(650)=>    "001111111010111000001000001111100001010111100010",
(651)=>    "001111111010111001110100001111100001010100111010",
(652)=>    "001111111010111011100010001111100001010010010000",
(653)=>    "001111111010111101001110001111100001001111101000",
(654)=>    "001111111010111110111010001111100001001100111110",
(655)=>    "001111111011000000100110001111100001001010010100",
(656)=>    "001111111011000010010010001111100001000111101010",
(657)=>    "001111111011000011111110001111100001000101000000",
(658)=>    "001111111011000101101000001111100001000010010110",
(659)=>    "001111111011000111010100001111100000111111101100",
(660)=>    "001111111011001000111110001111100000111101000010",
(661)=>    "001111111011001010101000001111100000111010010110",
(662)=>    "001111111011001100010010001111100000110111101100",
(663)=>    "001111111011001101111100001111100000110101000010",
(664)=>    "001111111011001111100110001111100000110010010110",
(665)=>    "001111111011010001010000001111100000101111101010",
(666)=>    "001111111011010010111000001111100000101101000000",
(667)=>    "001111111011010100100010001111100000101010010100",
(668)=>    "001111111011010110001010001111100000100111101000",
(669)=>    "001111111011010111110010001111100000100100111100",
(670)=>    "001111111011011001011010001111100000100010010000",
(671)=>    "001111111011011011000010001111100000011111100100",
(672)=>    "001111111011011100101010001111100000011100111000",
(673)=>    "001111111011011110010000001111100000011010001010",
(674)=>    "001111111011011111111000001111100000010111011110",
(675)=>    "001111111011100001011110001111100000010100110010",
(676)=>    "001111111011100011000100001111100000010010000100",
(677)=>    "001111111011100100101010001111100000001111011000",
(678)=>    "001111111011100110010000001111100000001100101010",
(679)=>    "001111111011100111110110001111100000001001111100",
(680)=>    "001111111011101001011100001111100000000111001110",
(681)=>    "001111111011101011000000001111100000000100100000",
(682)=>    "001111111011101100100110001111100000000001110100",
(683)=>    "001111111011101110001010001111001111111110001000",
(684)=>    "001111111011101111101110001111001111111000101100",
(685)=>    "001111111011110001010010001111001111110011010000",
(686)=>    "001111111011110010110110001111001111101101110100",
(687)=>    "001111111011110100011010001111001111101000011000",
(688)=>    "001111111011110101111110001111001111100010111000",
(689)=>    "001111111011110111100000001111001111011101011100",
(690)=>    "001111111011111001000010001111001111010111111100",
(691)=>    "001111111011111010100110001111001111010010011100",
(692)=>    "001111111011111100001000001111001111001101000000",
(693)=>    "001111111011111101101010001111001111000111100000",
(694)=>    "001111111011111111001010001111001111000010000000",
(695)=>    "001111111100000000101100001111001110111100100000",
(696)=>    "001111111100000010001110001111001110110111000000",
(697)=>    "001111111100000011101110001111001110110001100000",
(698)=>    "001111111100000101001110001111001110101100000000",
(699)=>    "001111111100000110101110001111001110100110011100",
(700)=>    "001111111100001000001110001111001110100000111100",
(701)=>    "001111111100001001101110001111001110011011011100",
(702)=>    "001111111100001011001110001111001110010101111000",
(703)=>    "001111111100001100101110001111001110010000011000",
(704)=>    "001111111100001110001100001111001110001010110100",
(705)=>    "001111111100001111101010001111001110000101010000",
(706)=>    "001111111100010001001010001111001101111111101100",
(707)=>    "001111111100010010101000001111001101111010001100",
(708)=>    "001111111100010100000110001111001101110100101000",
(709)=>    "001111111100010101100010001111001101101111000100",
(710)=>    "001111111100010111000000001111001101101001100000",
(711)=>    "001111111100011000011100001111001101100011111100",
(712)=>    "001111111100011001111010001111001101011110010100",
(713)=>    "001111111100011011010110001111001101011000110000",
(714)=>    "001111111100011100110010001111001101010011001100",
(715)=>    "001111111100011110001110001111001101001101100100",
(716)=>    "001111111100011111101010001111001101001000000000",
(717)=>    "001111111100100001000110001111001101000010011000",
(718)=>    "001111111100100010100000001111001100111100110100",
(719)=>    "001111111100100011111100001111001100110111001100",
(720)=>    "001111111100100101010110001111001100110001100100",
(721)=>    "001111111100100110110000001111001100101011111100",
(722)=>    "001111111100101000001010001111001100100110010100",
(723)=>    "001111111100101001100100001111001100100000110000",
(724)=>    "001111111100101010111110001111001100011011000100",
(725)=>    "001111111100101100010110001111001100010101011100",
(726)=>    "001111111100101101110000001111001100001111110100",
(727)=>    "001111111100101111001000001111001100001010001100",
(728)=>    "001111111100110000100000001111001100000100100100",
(729)=>    "001111111100110001111000001111001011111110111000",
(730)=>    "001111111100110011010000001111001011111001010000",
(731)=>    "001111111100110100101000001111001011110011100100",
(732)=>    "001111111100110101111110001111001011101101111100",
(733)=>    "001111111100110111010110001111001011101000010000",
(734)=>    "001111111100111000101100001111001011100010100100",
(735)=>    "001111111100111010000010001111001011011100111100",
(736)=>    "001111111100111011011000001111001011010111010000",
(737)=>    "001111111100111100101110001111001011010001100100",
(738)=>    "001111111100111110000100001111001011001011111000",
(739)=>    "001111111100111111011010001111001011000110001100",
(740)=>    "001111111101000000101110001111001011000000100000",
(741)=>    "001111111101000010000100001111001010111010110100",
(742)=>    "001111111101000011011000001111001010110101000100",
(743)=>    "001111111101000100101100001111001010101111011000",
(744)=>    "001111111101000110000000001111001010101001101100",
(745)=>    "001111111101000111010100001111001010100011111100",
(746)=>    "001111111101001000100110001111001010011110010000",
(747)=>    "001111111101001001111010001111001010011000100000",
(748)=>    "001111111101001011001100001111001010010010110100",
(749)=>    "001111111101001100011110001111001010001101000100",
(750)=>    "001111111101001101110000001111001010000111010100",
(751)=>    "001111111101001111000010001111001010000001100100",
(752)=>    "001111111101010000010100001111001001111011110100",
(753)=>    "001111111101010001100110001111001001110110000100",
(754)=>    "001111111101010010110110001111001001110000010100",
(755)=>    "001111111101010100001000001111001001101010100100",
(756)=>    "001111111101010101011000001111001001100100110100",
(757)=>    "001111111101010110101000001111001001011111000100",
(758)=>    "001111111101010111111000001111001001011001010100",
(759)=>    "001111111101011001001000001111001001010011100100",
(760)=>    "001111111101011010011000001111001001001101110000",
(761)=>    "001111111101011011100110001111001001001000000000",
(762)=>    "001111111101011100110100001111001001000010001100",
(763)=>    "001111111101011110000100001111001000111100011100",
(764)=>    "001111111101011111010010001111001000110110101000",
(765)=>    "001111111101100000100000001111001000110000110100",
(766)=>    "001111111101100001101110001111001000101011000100",
(767)=>    "001111111101100010111010001111001000100101010000",
(768)=>    "001111111101100100001000001111001000011111011100",
(769)=>    "001111111101100101010100001111001000011001101000",
(770)=>    "001111111101100110100010001111001000010011110100",
(771)=>    "001111111101100111101110001111001000001110000000",
(772)=>    "001111111101101000111010001111001000001000001100",
(773)=>    "001111111101101010000100001111001000000010011000",
(774)=>    "001111111101101011010000001111000111111100100100",
(775)=>    "001111111101101100011100001111000111110110101100",
(776)=>    "001111111101101101100110001111000111110000111000",
(777)=>    "001111111101101110110000001111000111101011000100",
(778)=>    "001111111101101111111010001111000111100101001100",
(779)=>    "001111111101110001000100001111000111011111011000",
(780)=>    "001111111101110010001110001111000111011001100000",
(781)=>    "001111111101110011011000001111000111010011101100",
(782)=>    "001111111101110100100000001111000111001101110100",
(783)=>    "001111111101110101101010001111000111000111111100",
(784)=>    "001111111101110110110010001111000111000010001000",
(785)=>    "001111111101110111111010001111000110111100010000",
(786)=>    "001111111101111001000010001111000110110110011000",
(787)=>    "001111111101111010001010001111000110110000100000",
(788)=>    "001111111101111011010010001111000110101010101000",
(789)=>    "001111111101111100011000001111000110100100110000",
(790)=>    "001111111101111101100000001111000110011110111000",
(791)=>    "001111111101111110100110001111000110011001000000",
(792)=>    "001111111101111111101100001111000110010011000100",
(793)=>    "001111111110000000110010001111000110001101001100",
(794)=>    "001111111110000001111000001111000110000111010100",
(795)=>    "001111111110000010111100001111000110000001011100",
(796)=>    "001111111110000100000010001111000101111011100000",
(797)=>    "001111111110000101000110001111000101110101101000",
(798)=>    "001111111110000110001100001111000101101111101100",
(799)=>    "001111111110000111010000001111000101101001110100",
(800)=>    "001111111110001000010100001111000101100011111000",
(801)=>    "001111111110001001010110001111000101011101111100",
(802)=>    "001111111110001010011010001111000101011000000100",
(803)=>    "001111111110001011011100001111000101010010001000",
(804)=>    "001111111110001100100000001111000101001100001100",
(805)=>    "001111111110001101100010001111000101000110010000",
(806)=>    "001111111110001110100100001111000101000000010100",
(807)=>    "001111111110001111100110001111000100111010011000",
(808)=>    "001111111110010000101000001111000100110100011100",
(809)=>    "001111111110010001101000001111000100101110100000",
(810)=>    "001111111110010010101010001111000100101000100100",
(811)=>    "001111111110010011101010001111000100100010101000",
(812)=>    "001111111110010100101010001111000100011100101000",
(813)=>    "001111111110010101101100001111000100010110101100",
(814)=>    "001111111110010110101010001111000100010000110000",
(815)=>    "001111111110010111101010001111000100001010110000",
(816)=>    "001111111110011000101010001111000100000100110100",
(817)=>    "001111111110011001101000001111000011111110110100",
(818)=>    "001111111110011010101000001111000011111000111000",
(819)=>    "001111111110011011100110001111000011110010111000",
(820)=>    "001111111110011100100100001111000011101100111100",
(821)=>    "001111111110011101100010001111000011100110111100",
(822)=>    "001111111110011110011110001111000011100000111100",
(823)=>    "001111111110011111011100001111000011011011000000",
(824)=>    "001111111110100000011000001111000011010101000000",
(825)=>    "001111111110100001010110001111000011001111000000",
(826)=>    "001111111110100010010010001111000011001001000000",
(827)=>    "001111111110100011001110001111000011000011000000",
(828)=>    "001111111110100100001010001111000010111101000000",
(829)=>    "001111111110100101000100001111000010110111000000",
(830)=>    "001111111110100110000000001111000010110001000000",
(831)=>    "001111111110100110111010001111000010101011000000",
(832)=>    "001111111110100111110110001111000010100101000000",
(833)=>    "001111111110101000110000001111000010011110111100",
(834)=>    "001111111110101001101010001111000010011000111100",
(835)=>    "001111111110101010100010001111000010010010111100",
(836)=>    "001111111110101011011100001111000010001100111000",
(837)=>    "001111111110101100010110001111000010000110111000",
(838)=>    "001111111110101101001110001111000010000000111000",
(839)=>    "001111111110101110000110001111000001111010110100",
(840)=>    "001111111110101110111110001111000001110100110100",
(841)=>    "001111111110101111110110001111000001101110110000",
(842)=>    "001111111110110000101110001111000001101000101100",
(843)=>    "001111111110110001100110001111000001100010101100",
(844)=>    "001111111110110010011100001111000001011100101000",
(845)=>    "001111111110110011010010001111000001010110100100",
(846)=>    "001111111110110100001010001111000001010000100000",
(847)=>    "001111111110110101000000001111000001001010100000",
(848)=>    "001111111110110101110110001111000001000100011100",
(849)=>    "001111111110110110101010001111000000111110011000",
(850)=>    "001111111110110111100000001111000000111000010100",
(851)=>    "001111111110111000010100001111000000110010010000",
(852)=>    "001111111110111001001010001111000000101100001100",
(853)=>    "001111111110111001111110001111000000100110001000",
(854)=>    "001111111110111010110010001111000000100000000100",
(855)=>    "001111111110111011100110001111000000011010000000",
(856)=>    "001111111110111100011000001111000000010011111000",
(857)=>    "001111111110111101001100001111000000001101110100",
(858)=>    "001111111110111101111110001111000000000111110000",
(859)=>    "001111111110111110110000001111000000000001101100",
(860)=>    "001111111110111111100100001110101111110111001000",
(861)=>    "001111111111000000010110001110101111101011000000",
(862)=>    "001111111111000001000110001110101111011110110000",
(863)=>    "001111111111000001111000001110101111010010101000",
(864)=>    "001111111111000010101000001110101111000110011000",
(865)=>    "001111111111000011011010001110101110111010010000",
(866)=>    "001111111111000100001010001110101110101110000000",
(867)=>    "001111111111000100111010001110101110100001111000",
(868)=>    "001111111111000101101010001110101110010101101000",
(869)=>    "001111111111000110011010001110101110001001011000",
(870)=>    "001111111111000111001000001110101101111101010000",
(871)=>    "001111111111000111111000001110101101110001000000",
(872)=>    "001111111111001000100110001110101101100100110000",
(873)=>    "001111111111001001010100001110101101011000100000",
(874)=>    "001111111111001010000010001110101101001100010000",
(875)=>    "001111111111001010110000001110101101000000001000",
(876)=>    "001111111111001011011110001110101100110011111000",
(877)=>    "001111111111001100001010001110101100100111101000",
(878)=>    "001111111111001100111000001110101100011011011000",
(879)=>    "001111111111001101100100001110101100001111001000",
(880)=>    "001111111111001110010000001110101100000010111000",
(881)=>    "001111111111001110111100001110101011110110100000",
(882)=>    "001111111111001111101000001110101011101010010000",
(883)=>    "001111111111010000010100001110101011011110000000",
(884)=>    "001111111111010000111110001110101011010001110000",
(885)=>    "001111111111010001101000001110101011000101100000",
(886)=>    "001111111111010010010100001110101010111001001000",
(887)=>    "001111111111010010111110001110101010101100111000",
(888)=>    "001111111111010011101000001110101010100000101000",
(889)=>    "001111111111010100010000001110101010010100010000",
(890)=>    "001111111111010100111010001110101010001000000000",
(891)=>    "001111111111010101100010001110101001111011110000",
(892)=>    "001111111111010110001100001110101001101111011000",
(893)=>    "001111111111010110110100001110101001100011001000",
(894)=>    "001111111111010111011100001110101001010110110000",
(895)=>    "001111111111011000000100001110101001001010100000",
(896)=>    "001111111111011000101010001110101000111110001000",
(897)=>    "001111111111011001010010001110101000110001110000",
(898)=>    "001111111111011001111000001110101000100101100000",
(899)=>    "001111111111011010011110001110101000011001001000",
(900)=>    "001111111111011011000100001110101000001100110000",
(901)=>    "001111111111011011101010001110101000000000100000",
(902)=>    "001111111111011100010000001110100111110100001000",
(903)=>    "001111111111011100110110001110100111100111110000",
(904)=>    "001111111111011101011010001110100111011011011000",
(905)=>    "001111111111011110000000001110100111001111000000",
(906)=>    "001111111111011110100100001110100111000010101000",
(907)=>    "001111111111011111001000001110100110110110011000",
(908)=>    "001111111111011111101100001110100110101010000000",
(909)=>    "001111111111100000001110001110100110011101101000",
(910)=>    "001111111111100000110010001110100110010001010000",
(911)=>    "001111111111100001010100001110100110000100111000",
(912)=>    "001111111111100001111000001110100101111000100000",
(913)=>    "001111111111100010011010001110100101101100001000",
(914)=>    "001111111111100010111100001110100101011111110000",
(915)=>    "001111111111100011011110001110100101010011010000",
(916)=>    "001111111111100011111110001110100101000110111000",
(917)=>    "001111111111100100100000001110100100111010100000",
(918)=>    "001111111111100101000000001110100100101110001000",
(919)=>    "001111111111100101100000001110100100100001110000",
(920)=>    "001111111111100110000000001110100100010101010000",
(921)=>    "001111111111100110100000001110100100001000111000",
(922)=>    "001111111111100111000000001110100011111100100000",
(923)=>    "001111111111100111100000001110100011110000001000",
(924)=>    "001111111111100111111110001110100011100011101000",
(925)=>    "001111111111101000011100001110100011010111010000",
(926)=>    "001111111111101000111010001110100011001010110000",
(927)=>    "001111111111101001011000001110100010111110011000",
(928)=>    "001111111111101001110110001110100010110010000000",
(929)=>    "001111111111101010010100001110100010100101100000",
(930)=>    "001111111111101010110000001110100010011001001000",
(931)=>    "001111111111101011001110001110100010001100101000",
(932)=>    "001111111111101011101010001110100010000000010000",
(933)=>    "001111111111101100000110001110100001110011110000",
(934)=>    "001111111111101100100010001110100001100111011000",
(935)=>    "001111111111101100111110001110100001011010111000",
(936)=>    "001111111111101101011000001110100001001110011000",
(937)=>    "001111111111101101110100001110100001000010000000",
(938)=>    "001111111111101110001110001110100000110101100000",
(939)=>    "001111111111101110101000001110100000101001000000",
(940)=>    "001111111111101111000010001110100000011100101000",
(941)=>    "001111111111101111011100001110100000010000001000",
(942)=>    "001111111111101111110110001110100000000011101000",
(943)=>    "001111111111110000001110001110001111101110100000",
(944)=>    "001111111111110000101000001110001111010101100000",
(945)=>    "001111111111110001000000001110001110111100100000",
(946)=>    "001111111111110001011000001110001110100011100000",
(947)=>    "001111111111110001110000001110001110001010100000",
(948)=>    "001111111111110010001000001110001101110001110000",
(949)=>    "001111111111110010011110001110001101011000110000",
(950)=>    "001111111111110010110110001110001100111111110000",
(951)=>    "001111111111110011001100001110001100100110110000",
(952)=>    "001111111111110011100010001110001100001101110000",
(953)=>    "001111111111110011111000001110001011110100110000",
(954)=>    "001111111111110100001110001110001011011011110000",
(955)=>    "001111111111110100100100001110001011000010110000",
(956)=>    "001111111111110100111000001110001010101001110000",
(957)=>    "001111111111110101001110001110001010010000110000",
(958)=>    "001111111111110101100010001110001001110111110000",
(959)=>    "001111111111110101110110001110001001011110110000",
(960)=>    "001111111111110110001010001110001001000101110000",
(961)=>    "001111111111110110011110001110001000101100110000",
(962)=>    "001111111111110110110000001110001000010011110000",
(963)=>    "001111111111110111000100001110000111111010110000",
(964)=>    "001111111111110111010110001110000111100001110000",
(965)=>    "001111111111110111101000001110000111001000110000",
(966)=>    "001111111111110111111010001110000110101111110000",
(967)=>    "001111111111111000001100001110000110010110100000",
(968)=>    "001111111111111000011110001110000101111101100000",
(969)=>    "001111111111111000101110001110000101100100100000",
(970)=>    "001111111111111001000000001110000101001011100000",
(971)=>    "001111111111111001010000001110000100110010100000",
(972)=>    "001111111111111001100000001110000100011001100000",
(973)=>    "001111111111111001110000001110000100000000010000",
(974)=>    "001111111111111010000000001110000011100111010000",
(975)=>    "001111111111111010001110001110000011001110010000",
(976)=>    "001111111111111010011110001110000010110101010000",
(977)=>    "001111111111111010101100001110000010011100000000",
(978)=>    "001111111111111010111010001110000010000011000000",
(979)=>    "001111111111111011001000001110000001101010000000",
(980)=>    "001111111111111011010110001110000001010001000000",
(981)=>    "001111111111111011100100001110000000110111110000",
(982)=>    "001111111111111011110010001110000000011110110000",
(983)=>    "001111111111111011111110001110000000000101110000",
(984)=>    "001111111111111100001010001101101111011001000000",
(985)=>    "001111111111111100010110001101101110100111000000",
(986)=>    "001111111111111100100010001101101101110101000000",
(987)=>    "001111111111111100101110001101101101000010100000",
(988)=>    "001111111111111100111010001101101100010000100000",
(989)=>    "001111111111111101000100001101101011011110000000",
(990)=>    "001111111111111101001110001101101010101100000000",
(991)=>    "001111111111111101011010001101101001111010000000",
(992)=>    "001111111111111101100100001101101001000111100000",
(993)=>    "001111111111111101101100001101101000010101100000",
(994)=>    "001111111111111101110110001101100111100011000000",
(995)=>    "001111111111111110000000001101100110110001000000",
(996)=>    "001111111111111110001000001101100101111111000000",
(997)=>    "001111111111111110010000001101100101001100100000",
(998)=>    "001111111111111110011000001101100100011010100000",
(999)=>    "001111111111111110100000001101100011101000000000",
(1000)=>    "001111111111111110101000001101100010110110000000",
(1001)=>    "001111111111111110110000001101100010000011100000",
(1002)=>    "001111111111111110110110001101100001010001100000",
(1003)=>    "001111111111111110111100001101100000011111000000",
(1004)=>    "001111111111111111000100001101001111011010000000",
(1005)=>    "001111111111111111001010001101001101110101000000",
(1006)=>    "001111111111111111010000001101001100010001000000",
(1007)=>    "001111111111111111010100001101001010101100000000",
(1008)=>    "001111111111111111011010001101001001001000000000",
(1009)=>    "001111111111111111011110001101000111100011000000",
(1010)=>    "001111111111111111100010001101000101111111000000",
(1011)=>    "001111111111111111100110001101000100011010000000",
(1012)=>    "001111111111111111101010001101000010110110000000",
(1013)=>    "001111111111111111101110001101000001010001000000",
(1014)=>    "001111111111111111110010001100101111011010000000",
(1015)=>    "001111111111111111110100001100101100010000000000",
(1016)=>    "001111111111111111111000001100101001001000000000",
(1017)=>    "001111111111111111111010001100100101111110000000",
(1018)=>    "001111111111111111111100001100100010110110000000",
(1019)=>    "001111111111111111111110001100001111011000000000",
(1020)=>    "001111111111111111111110001100001001001000000000",
(1021)=>    "001111111111111111111110001100000010110100000000",
(1022)=>    "001111111111111111111110001011101001001000000000",
(1023)=>    "010000010000000000000000001011001001000000000000"

);
end package;
