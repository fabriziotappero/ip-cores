library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library work;
use work.USB_TMC_IP_Defs.all;
use work.USB_TMC_cmp.all;



entity USB_TMC is
  port(
       i_nReset,
       i_SYSCLK : std_logic;
  
  
  
  
  );  
end USB_TMC;



architecture FSM of USB_TMC is



begin





end FSM;