-- obj_code_pkg -- Object code in VHDL constant table for BRAM initialization.
-- Generated automatically with script 'build_rom.py'.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.l80pkg.all;

package obj_code_pkg is

constant obj_code : obj_code_t(0 to 372) := (
    X"c3", X"60", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c3", X"12", X"01", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c3", X"1e", X"01", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"fb", X"c9", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c3", X"2a", X"01", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"31", X"da", X"01", X"21", X"74", X"01", X"22", X"75", 
    X"01", X"21", X"7a", X"01", X"22", X"77", X"01", X"3e", 
    X"00", X"32", X"79", X"01", X"3e", X"00", X"d3", X"86", 
    X"3e", X"0b", X"d3", X"88", X"fb", X"21", X"02", X"01", 
    X"cd", X"66", X"01", X"3e", X"01", X"32", X"73", X"01", 
    X"3e", X"01", X"d3", X"86", X"3a", X"73", X"01", X"fe", 
    X"04", X"ca", X"9c", X"00", X"fe", X"01", X"c2", X"fb", 
    X"00", X"c3", X"8c", X"00", X"3e", X"00", X"d3", X"86", 
    X"3e", X"01", X"32", X"73", X"01", X"3e", X"02", X"d3", 
    X"86", X"3a", X"73", X"01", X"fe", X"02", X"ca", X"b9", 
    X"00", X"fe", X"01", X"c2", X"fb", X"00", X"c3", X"a9", 
    X"00", X"af", X"d3", X"86", X"3e", X"01", X"32", X"73", 
    X"01", X"3e", X"03", X"d3", X"86", X"3a", X"73", X"01", 
    X"fe", X"05", X"ca", X"d5", X"00", X"fe", X"01", X"c2", 
    X"fb", X"00", X"c3", X"c5", X"00", X"af", X"d3", X"86", 
    X"3a", X"79", X"01", X"fe", X"0f", X"c2", X"d8", X"00", 
    X"21", X"7a", X"01", X"11", X"02", X"01", X"1a", X"fe", 
    X"24", X"ca", X"f5", X"00", X"be", X"c2", X"fb", X"00", 
    X"23", X"13", X"c3", X"e6", X"00", X"3e", X"80", X"d3", 
    X"86", X"f3", X"76", X"3e", X"40", X"d3", X"86", X"c3", 
    X"f9", X"00", X"0a", X"0d", X"0a", X"48", X"65", X"6c", 
    X"6c", X"6f", X"20", X"57", X"6f", X"72", X"6c", X"64", 
    X"21", X"24", X"f5", X"3a", X"73", X"01", X"07", X"07", 
    X"32", X"73", X"01", X"f1", X"fb", X"c9", X"f5", X"3a", 
    X"73", X"01", X"c6", X"01", X"32", X"73", X"01", X"f1", 
    X"fb", X"c9", X"e5", X"f5", X"db", X"81", X"e6", X"20", 
    X"ca", X"48", X"01", X"3e", X"20", X"d3", X"81", X"db", 
    X"80", X"2a", X"77", X"01", X"77", X"23", X"22", X"77", 
    X"01", X"3a", X"79", X"01", X"3c", X"32", X"79", X"01", 
    X"db", X"81", X"e6", X"10", X"ca", X"62", X"01", X"3e", 
    X"10", X"d3", X"81", X"2a", X"75", X"01", X"7e", X"fe", 
    X"24", X"ca", X"62", X"01", X"23", X"22", X"75", X"01", 
    X"d3", X"80", X"f1", X"e1", X"fb", X"c9", X"7e", X"23", 
    X"22", X"75", X"01", X"fe", X"24", X"ca", X"72", X"01", 
    X"d3", X"80", X"c9", X"00", X"24" 
);

end package obj_code_pkg;
