-- obj_code_pkg -- Object code in VHDL constant table for BRAM initialization.
-- Generated automatically with script 'build_rom.py'.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.l80pkg.all;

package obj_code_pkg is

constant obj_code : obj_code_t(0 to 235) := (
    X"c3", X"60", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c9", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"c3", X"a7", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", 
    X"31", X"50", X"01", X"21", X"eb", X"00", X"22", X"ec", 
    X"00", X"21", X"f0", X"00", X"22", X"ee", X"00", X"3e", 
    X"14", X"d3", X"83", X"3e", X"58", X"d3", X"82", X"3e", 
    X"00", X"d3", X"86", X"3e", X"08", X"d3", X"88", X"fb", 
    X"21", X"96", X"00", X"cd", X"de", X"00", X"db", X"84", 
    X"4f", X"07", X"07", X"81", X"d3", X"86", X"c3", X"86", 
    X"00", X"f3", X"76", X"c3", X"93", X"00", X"0a", X"0d", 
    X"0a", X"48", X"65", X"6c", X"6c", X"6f", X"20", X"57", 
    X"6f", X"72", X"6c", X"64", X"21", X"24", X"00", X"e5", 
    X"f5", X"db", X"81", X"e6", X"20", X"ca", X"c0", X"00", 
    X"3e", X"20", X"d3", X"81", X"db", X"80", X"d3", X"86", 
    X"2a", X"ee", X"00", X"77", X"23", X"22", X"ee", X"00", 
    X"db", X"81", X"e6", X"10", X"ca", X"da", X"00", X"3e", 
    X"10", X"d3", X"81", X"2a", X"ec", X"00", X"7e", X"fe", 
    X"24", X"ca", X"da", X"00", X"23", X"22", X"ec", X"00", 
    X"d3", X"80", X"f1", X"e1", X"fb", X"c9", X"7e", X"23", 
    X"22", X"ec", X"00", X"fe", X"24", X"ca", X"ea", X"00", 
    X"d3", X"80", X"c9", X"24" 
);

end package obj_code_pkg;
