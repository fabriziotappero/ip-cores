`timescale 1 ns/1 ps
package ahb_wb_pkg;
import global::*;
	`include "../avm_svtb/ahb_wb_stim_gen.svh"
	`include "../avm_svtb/ahb_wb_driver.svh"
	`include "../avm_svtb/ahb_wb_responder.svh"
	`include "../avm_svtb/ahb_wb_monitor.svh"
	`include "../avm_svtb/ahb_wb_scoreboard.svh"
	`include "../avm_svtb/ahb_wb_coverage.svh"
	`include "../avm_svtb/ahb_wb_env.svh"
endpackage
	
