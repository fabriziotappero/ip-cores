-------------------------------------------------------------------------------
--
-- The stack unit.
--
-- $Id: t400_stack-c.vhd 179 2009-04-01 19:48:38Z arniml $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_stack_rtl_c0 of t400_stack is

  for rtl
  end for;

end t400_stack_rtl_c0;
