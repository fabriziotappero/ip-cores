-- Rom file for twiddle factors 
-- ../../../rtl/vhdl/WISHBONE_FFT/rom3.vhd contains 64 points of 16 width 
--  for a 1024 point fft.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;


ENTITY rom3 IS
         GENERIC(
        data_width : integer :=16;
        address_width : integer :=6
    );
    PORT(
        clk :in std_logic;
        address :in std_logic_vector (5      downto 0);
        datar : OUT std_logic_vector (data_width-1 DOWNTO 0) ;
        datai : OUT std_logic_vector (data_width-1 DOWNTO 0)
    );
end rom3;
ARCHITECTURE behavior OF rom3 IS

 BEGIN

process (address,clk)
begin
    	if(rising_edge(clk)) then 
 case address is
        when "000000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "000001" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "000010" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "000011" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "000100" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "000101" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "000110" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "000111" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "001000" => datar <= "0000000000000000";datai <= "1000000000000001"; --256
        when "001001" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "001010" => datar <= "1100111100000101";datai <= "1000100110111111"; --320
        when "001011" => datar <= "1011100011100100";datai <= "1001010110010011"; --352
        when "001100" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "001101" => datar <= "1001010110010011";datai <= "1011100011100100"; --416
        when "001110" => datar <= "1000100110111111";datai <= "1100111100000101"; --448
        when "001111" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "010000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "010001" => datar <= "0111111101100001";datai <= "1111001101110100"; --16
        when "010010" => datar <= "0111110110001001";datai <= "1110011100000111"; --32
        when "010011" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "010100" => datar <= "0111011001000001";datai <= "1100111100000101"; --64
        when "010101" => datar <= "0111000011100010";datai <= "1100001110101010"; --80
        when "010110" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "010111" => datar <= "0110001011110001";datai <= "1010111011001101"; --112
        when "011000" => datar <= "0101101010000010";datai <= "1010010101111110"; --128
        when "011001" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "011010" => datar <= "0100011100011100";datai <= "1001010110010011"; --160
        when "011011" => datar <= "0011110001010110";datai <= "1000111100011110"; --176
        when "011100" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "011101" => datar <= "0010010100101000";datai <= "1000010110000100"; --208
        when "011110" => datar <= "0001100011111001";datai <= "1000001001110111"; --224
        when "011111" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "100000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when "100001" => datar <= "0111101001111100";datai <= "1101101011011000"; --48
        when "100010" => datar <= "0110101001101101";datai <= "1011100011100100"; --96
        when "100011" => datar <= "0101000100110011";datai <= "1001110100001111"; --144
        when "100100" => datar <= "0011000011111011";datai <= "1000100110111111"; --192
        when "100101" => datar <= "0000110010001100";datai <= "1000000010011111"; --240
        when "100110" => datar <= "1110011100000111";datai <= "1000001001110111"; --288
        when "100111" => datar <= "1100001110101010";datai <= "1000111100011110"; --336
        when "101000" => datar <= "1010010101111110";datai <= "1010010101111110"; --384
        when "101001" => datar <= "1000111100011110";datai <= "1100001110101010"; --432
        when "101010" => datar <= "1000001001110111";datai <= "1110011100000111"; --480
        when "101011" => datar <= "1000000010011111";datai <= "0000110010001100"; --528
        when "101100" => datar <= "1000100110111111";datai <= "0011000011111011"; --576
        when "101101" => datar <= "1001110100001111";datai <= "0101000100110011"; --624
        when "101110" => datar <= "1011100011100100";datai <= "0110101001101101"; --672
        when "101111" => datar <= "1101101011011000";datai <= "0111101001111100"; --720
           when "110000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "110111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111000" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111001" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111010" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111011" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111100" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111101" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111110" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
           when "111111" => datar <= "0111111111111111";datai <= "0000000000000000"; --0
        when others => for i in data_width-1 downto 0 loop
            datar(i)<='0';datai(i)<='0';end loop;
    end case;

    end if;

end process;
END behavior;
