/* verilator lint_off UNUSED */
/* verilator lint_off CASEX */
/* verilator lint_off PINNOCONNECT */
/* verilator lint_off PINMISSING */
/* verilator lint_off UNOPTFLAT */

module uart_16750 ( CLK, RST, BAUDCE, CS, WR, RD, A, DIN, DOUT, DDIS, INT, 
        OUT1N, OUT2N, RCLK, BAUDOUTN, RTSN, DTRN, CTSN, DSRN, DCDN, RIN, SIN, 
        SOUT );
  input [2:0] A;
  input [7:0] DIN;
  output [7:0] DOUT;
  input CLK, RST, BAUDCE, CS, WR, RD, RCLK, CTSN, DSRN, DCDN, RIN, SIN;
  output DDIS, INT, OUT1N, OUT2N, BAUDOUTN, RTSN, DTRN, SOUT;
  wire   N48, iWriteFE, iReadFE, iSINr, iCTSNs, iDSRNs, iDCDNs, iRINs,
         iBaudtick2x, iCTSn, iDSRn, iDCDn, iRIn, iTHRInterrupt, iCharTimeout,
         iIIR_6, iLSR_THRERE, N66, iRXFIFOEmpty, iRXFIFOWrite, N94, N95,
         iFCR_5, iPERE, iFERE, iBIRE, iLSR_FIFOERR, iRXFIFOClear, N130, N131,
         N132, N133, N134, N135, N146, iTXFIFOEmpty, iTXRunning, iRTS, N154,
         N155, N156, N157, iCTSnFE, iDSRnFE, iRInFE, iDCDnFE, iBaudtick16x,
         iRCLK, iTXFIFORead, iTXFIFO64Full, \iTXFIFOUsage[4] , N169,
         iRXFIFO64Full, iTXStart, iTXFinished, iSOUT, iSIN, iRXPE, iRXFE,
         iRXBI, N181, N182, N183, State_snps_wire, N190, N191, N197, N198,
         N199, N200, N201, N202, \U3/U1/Z_0 , n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n371, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n424, n425, n426, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n440,
         n441, n442, n443, n444, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, \UART_ED_WRITE/n1 , \UART_ED_WRITE/iDd , \UART_ED_READ/n1 ,
         \UART_ED_READ/iDd , \UART_IS_SIN/n1 , \UART_IS_SIN/iD[0] ,
         \UART_IS_CTS/n1 , \UART_IS_CTS/iD[0] , \UART_IS_DSR/n1 ,
         \UART_IS_DSR/iD[0] , \UART_IS_DCD/n1 , \UART_IS_DCD/iD[0] ,
         \UART_IS_RI/n1 , \UART_IS_RI/iD[0] , \UART_IF_CTS/n8 ,
         \UART_IF_CTS/n7 , \UART_IF_CTS/n6 , \UART_IF_CTS/n5 ,
         \UART_IF_CTS/n4 , \UART_IF_CTS/n2 , \UART_IF_CTS/n1 ,
         \UART_IF_CTS/n18 , \UART_IF_CTS/n17 , \UART_IF_CTS/n16 ,
         \UART_IF_CTS/iCount[0] , \UART_IF_CTS/iCount[1] , \UART_IF_DSR/n11 ,
         \UART_IF_DSR/n10 , \UART_IF_DSR/n9 , \UART_IF_DSR/n8 ,
         \UART_IF_DSR/n7 , \UART_IF_DSR/n6 , \UART_IF_DSR/n5 ,
         \UART_IF_DSR/n4 , \UART_IF_DSR/n2 , \UART_IF_DSR/n1 ,
         \UART_IF_DSR/iCount[0] , \UART_IF_DSR/iCount[1] , \UART_IF_DCD/n11 ,
         \UART_IF_DCD/n10 , \UART_IF_DCD/n9 , \UART_IF_DCD/n7 ,
         \UART_IF_DCD/n6 , \UART_IF_DCD/n5 , \UART_IF_DCD/n4 ,
         \UART_IF_DCD/n2 , \UART_IF_DCD/n1 , \UART_IF_DCD/iCount[0] ,
         \UART_IF_DCD/iCount[1] , \UART_IF_RI/n11 , \UART_IF_RI/n10 ,
         \UART_IF_RI/n9 , \UART_IF_RI/n7 , \UART_IF_RI/n6 , \UART_IF_RI/n5 ,
         \UART_IF_RI/n4 , \UART_IF_RI/n3 , \UART_IF_RI/n2 , \UART_IF_RI/n1 ,
         \UART_IF_RI/iCount[0] , \UART_IF_RI/iCount[1] , \UART_IIC/n9 ,
         \UART_IIC/n8 , \UART_IIC/n7 , \UART_IIC/n6 , \UART_IIC/n5 ,
         \UART_IIC/n4 , \UART_IIC/n3 , \UART_IIC/n2 , \UART_IIC/n1 ,
         \UART_IIC/N22 , \UART_IIC/N21 , \UART_IIC/N20 , \UART_IIC/N19 ,
         \UART_IIC/IIR[0] , \UART_IIC_THRE_ED/n1 , \UART_IIC_THRE_ED/iDd ,
         \UART_PEDET/n1 , \UART_PEDET/iDd , \UART_FEDET/n1 , \UART_FEDET/iDd ,
         \UART_BIDET/n1 , \UART_BIDET/iDd , \UART_ED_CTS/n1 ,
         \UART_ED_CTS/iDd , \UART_ED_DSR/n1 , \UART_ED_DSR/iDd ,
         \UART_ED_RI/n1 , \UART_ED_RI/iDd , \UART_ED_DCD/n1 ,
         \UART_ED_DCD/iDd , \UART_BG16/n72 , \UART_BG16/n71 , \UART_BG16/n70 ,
         \UART_BG16/n69 , \UART_BG16/n68 , \UART_BG16/n67 , \UART_BG16/n66 ,
         \UART_BG16/n65 , \UART_BG16/n64 , \UART_BG16/n63 , \UART_BG16/n62 ,
         \UART_BG16/n61 , \UART_BG16/n60 , \UART_BG16/n59 , \UART_BG16/n58 ,
         \UART_BG16/n57 , \UART_BG16/n56 , \UART_BG16/n39 , \UART_BG16/n38 ,
         \UART_BG16/n37 , \UART_BG16/n35 , \UART_BG16/n33 , \UART_BG16/n32 ,
         \UART_BG16/n31 , \UART_BG16/n30 , \UART_BG16/n29 , \UART_BG16/n28 ,
         \UART_BG16/n27 , \UART_BG16/n26 , \UART_BG16/n25 , \UART_BG16/n24 ,
         \UART_BG16/n23 , \UART_BG16/n22 , \UART_BG16/n21 , \UART_BG16/n20 ,
         \UART_BG16/n19 , \UART_BG16/n18 , \UART_BG16/n17 , \UART_BG16/n16 ,
         \UART_BG16/n15 , \UART_BG16/n14 , \UART_BG16/n13 , \UART_BG16/n12 ,
         \UART_BG16/n11 , \UART_BG16/n10 , \UART_BG16/n9 , \UART_BG16/n8 ,
         \UART_BG16/n7 , \UART_BG16/n6 , \UART_BG16/n5 , \UART_BG16/n4 ,
         \UART_BG16/n2 , \UART_BG16/n1 , \UART_BG16/n55 , \UART_BG16/n54 ,
         \UART_BG16/n53 , \UART_BG16/n52 , \UART_BG16/n51 , \UART_BG16/n50 ,
         \UART_BG16/n49 , \UART_BG16/n48 , \UART_BG16/n47 , \UART_BG16/n46 ,
         \UART_BG16/n45 , \UART_BG16/n44 , \UART_BG16/n43 , \UART_BG16/n42 ,
         \UART_BG16/n41 , \UART_BG16/n40 , \UART_BG16/N40 , \UART_BG16/N22 ,
         \UART_BG16/N21 , \UART_BG16/N20 , \UART_BG16/N19 , \UART_BG16/N18 ,
         \UART_BG16/N17 , \UART_BG16/N16 , \UART_BG16/N15 , \UART_BG16/N14 ,
         \UART_BG16/N13 , \UART_BG16/N12 , \UART_BG16/N11 , \UART_BG16/N10 ,
         \UART_BG16/N9 , \UART_BG16/N8 , \UART_BG16/iCounter[0] ,
         \UART_BG16/iCounter[1] , \UART_BG16/iCounter[2] ,
         \UART_BG16/iCounter[3] , \UART_BG16/iCounter[4] ,
         \UART_BG16/iCounter[5] , \UART_BG16/iCounter[6] ,
         \UART_BG16/iCounter[7] , \UART_BG16/iCounter[8] ,
         \UART_BG16/iCounter[9] , \UART_BG16/iCounter[10] ,
         \UART_BG16/iCounter[11] , \UART_BG16/iCounter[12] ,
         \UART_BG16/iCounter[13] , \UART_BG16/iCounter[14] ,
         \UART_BG16/iCounter[15] , \UART_BG2/n2 , \UART_BG2/n1 , \UART_BG2/n6 ,
         \UART_BG2/n4 , \UART_BG2/n3 , \UART_BG2/N14 , \UART_BG2/iCounter[0] ,
         \UART_BG2/iCounter[1] , \UART_BG2/iCounter[2] , \UART_RCLK/n1 ,
         \UART_RCLK/iDd , \UART_TXFF/n373 , \UART_TXFF/n372 , \UART_TXFF/n371 ,
         \UART_TXFF/n370 , \UART_TXFF/n369 , \UART_TXFF/n368 ,
         \UART_TXFF/n367 , \UART_TXFF/n366 , \UART_TXFF/n365 ,
         \UART_TXFF/n364 , \UART_TXFF/n363 , \UART_TXFF/n362 ,
         \UART_TXFF/n361 , \UART_TXFF/n360 , \UART_TXFF/n359 ,
         \UART_TXFF/n358 , \UART_TXFF/n356 , \UART_TXFF/n355 ,
         \UART_TXFF/n354 , \UART_TXFF/n350 , \UART_TXFF/n349 ,
         \UART_TXFF/n348 , \UART_TXFF/n347 , \UART_TXFF/n346 ,
         \UART_TXFF/n345 , \UART_TXFF/n344 , \UART_TXFF/n343 ,
         \UART_TXFF/n342 , \UART_TXFF/n341 , \UART_TXFF/n340 ,
         \UART_TXFF/n339 , \UART_TXFF/n338 , \UART_TXFF/n337 ,
         \UART_TXFF/n336 , \UART_TXFF/n335 , \UART_TXFF/n334 ,
         \UART_TXFF/n333 , \UART_TXFF/n332 , \UART_TXFF/n331 ,
         \UART_TXFF/n330 , \UART_TXFF/n329 , \UART_TXFF/n328 ,
         \UART_TXFF/n327 , \UART_TXFF/n326 , \UART_TXFF/n325 ,
         \UART_TXFF/n324 , \UART_TXFF/n323 , \UART_TXFF/n322 ,
         \UART_TXFF/n321 , \UART_TXFF/n320 , \UART_TXFF/n319 ,
         \UART_TXFF/n318 , \UART_TXFF/n317 , \UART_TXFF/n316 ,
         \UART_TXFF/n315 , \UART_TXFF/n314 , \UART_TXFF/n313 ,
         \UART_TXFF/n312 , \UART_TXFF/n311 , \UART_TXFF/n310 ,
         \UART_TXFF/n309 , \UART_TXFF/n308 , \UART_TXFF/n307 ,
         \UART_TXFF/n306 , \UART_TXFF/n305 , \UART_TXFF/n304 ,
         \UART_TXFF/n303 , \UART_TXFF/n302 , \UART_TXFF/n301 ,
         \UART_TXFF/n300 , \UART_TXFF/n299 , \UART_TXFF/n298 ,
         \UART_TXFF/n297 , \UART_TXFF/n296 , \UART_TXFF/n295 ,
         \UART_TXFF/n294 , \UART_TXFF/n293 , \UART_TXFF/n292 ,
         \UART_TXFF/n291 , \UART_TXFF/n290 , \UART_TXFF/n289 ,
         \UART_TXFF/n288 , \UART_TXFF/n287 , \UART_TXFF/n286 ,
         \UART_TXFF/n285 , \UART_TXFF/n284 , \UART_TXFF/n283 ,
         \UART_TXFF/n282 , \UART_TXFF/n281 , \UART_TXFF/n280 ,
         \UART_TXFF/n279 , \UART_TXFF/n278 , \UART_TXFF/n277 ,
         \UART_TXFF/n276 , \UART_TXFF/n275 , \UART_TXFF/n274 ,
         \UART_TXFF/n273 , \UART_TXFF/n272 , \UART_TXFF/n271 ,
         \UART_TXFF/n270 , \UART_TXFF/n269 , \UART_TXFF/n268 ,
         \UART_TXFF/n267 , \UART_TXFF/n266 , \UART_TXFF/n265 ,
         \UART_TXFF/n264 , \UART_TXFF/n263 , \UART_TXFF/n262 ,
         \UART_TXFF/n261 , \UART_TXFF/n260 , \UART_TXFF/n259 ,
         \UART_TXFF/n258 , \UART_TXFF/n257 , \UART_TXFF/n256 ,
         \UART_TXFF/n255 , \UART_TXFF/n254 , \UART_TXFF/n253 ,
         \UART_TXFF/n252 , \UART_TXFF/n251 , \UART_TXFF/n250 ,
         \UART_TXFF/n249 , \UART_TXFF/n248 , \UART_TXFF/n247 ,
         \UART_TXFF/n246 , \UART_TXFF/n245 , \UART_TXFF/n244 ,
         \UART_TXFF/n243 , \UART_TXFF/n242 , \UART_TXFF/n240 ,
         \UART_TXFF/n239 , \UART_TXFF/n238 , \UART_TXFF/n237 ,
         \UART_TXFF/n236 , \UART_TXFF/n235 , \UART_TXFF/n234 ,
         \UART_TXFF/n233 , \UART_TXFF/n232 , \UART_TXFF/n231 ,
         \UART_TXFF/n230 , \UART_TXFF/n229 , \UART_TXFF/n228 ,
         \UART_TXFF/n227 , \UART_TXFF/n226 , \UART_TXFF/n225 ,
         \UART_TXFF/n224 , \UART_TXFF/n223 , \UART_TXFF/n222 ,
         \UART_TXFF/n221 , \UART_TXFF/n220 , \UART_TXFF/n219 ,
         \UART_TXFF/n218 , \UART_TXFF/n217 , \UART_TXFF/n216 ,
         \UART_TXFF/n215 , \UART_TXFF/n214 , \UART_TXFF/n213 ,
         \UART_TXFF/n212 , \UART_TXFF/n211 , \UART_TXFF/n210 ,
         \UART_TXFF/n209 , \UART_TXFF/n208 , \UART_TXFF/n207 ,
         \UART_TXFF/n206 , \UART_TXFF/n205 , \UART_TXFF/n204 ,
         \UART_TXFF/n203 , \UART_TXFF/n202 , \UART_TXFF/n201 ,
         \UART_TXFF/n200 , \UART_TXFF/n199 , \UART_TXFF/n198 ,
         \UART_TXFF/n197 , \UART_TXFF/n196 , \UART_TXFF/n195 ,
         \UART_TXFF/n194 , \UART_TXFF/n193 , \UART_TXFF/n192 ,
         \UART_TXFF/n191 , \UART_TXFF/n190 , \UART_TXFF/n189 ,
         \UART_TXFF/n188 , \UART_TXFF/n187 , \UART_TXFF/n186 ,
         \UART_TXFF/n185 , \UART_TXFF/n184 , \UART_TXFF/n183 ,
         \UART_TXFF/n182 , \UART_TXFF/n181 , \UART_TXFF/n180 ,
         \UART_TXFF/n179 , \UART_TXFF/n178 , \UART_TXFF/n177 ,
         \UART_TXFF/n176 , \UART_TXFF/n175 , \UART_TXFF/n174 ,
         \UART_TXFF/n173 , \UART_TXFF/n172 , \UART_TXFF/n171 ,
         \UART_TXFF/n170 , \UART_TXFF/n169 , \UART_TXFF/n168 ,
         \UART_TXFF/n167 , \UART_TXFF/n166 , \UART_TXFF/n165 ,
         \UART_TXFF/n164 , \UART_TXFF/n163 , \UART_TXFF/n162 ,
         \UART_TXFF/n161 , \UART_TXFF/n160 , \UART_TXFF/n159 ,
         \UART_TXFF/n158 , \UART_TXFF/n157 , \UART_TXFF/n156 ,
         \UART_TXFF/n155 , \UART_TXFF/n154 , \UART_TXFF/n153 ,
         \UART_TXFF/n152 , \UART_TXFF/n151 , \UART_TXFF/n150 ,
         \UART_TXFF/n149 , \UART_TXFF/n148 , \UART_TXFF/n147 ,
         \UART_TXFF/n146 , \UART_TXFF/n145 , \UART_TXFF/n144 ,
         \UART_TXFF/n143 , \UART_TXFF/n142 , \UART_TXFF/n141 ,
         \UART_TXFF/n140 , \UART_TXFF/n139 , \UART_TXFF/n138 ,
         \UART_TXFF/n137 , \UART_TXFF/n136 , \UART_TXFF/n135 ,
         \UART_TXFF/n134 , \UART_TXFF/n133 , \UART_TXFF/n132 ,
         \UART_TXFF/n131 , \UART_TXFF/n130 , \UART_TXFF/n129 ,
         \UART_TXFF/n128 , \UART_TXFF/n127 , \UART_TXFF/n126 ,
         \UART_TXFF/n125 , \UART_TXFF/n124 , \UART_TXFF/n123 ,
         \UART_TXFF/n122 , \UART_TXFF/n121 , \UART_TXFF/n120 ,
         \UART_TXFF/n119 , \UART_TXFF/n118 , \UART_TXFF/n117 ,
         \UART_TXFF/n116 , \UART_TXFF/n115 , \UART_TXFF/n114 ,
         \UART_TXFF/n113 , \UART_TXFF/n112 , \UART_TXFF/n111 ,
         \UART_TXFF/n110 , \UART_TXFF/n109 , \UART_TXFF/n108 ,
         \UART_TXFF/n107 , \UART_TXFF/n106 , \UART_TXFF/n105 ,
         \UART_TXFF/n104 , \UART_TXFF/n103 , \UART_TXFF/n102 ,
         \UART_TXFF/n101 , \UART_TXFF/n100 , \UART_TXFF/n99 , \UART_TXFF/n98 ,
         \UART_TXFF/n97 , \UART_TXFF/n96 , \UART_TXFF/n95 , \UART_TXFF/n94 ,
         \UART_TXFF/n93 , \UART_TXFF/n92 , \UART_TXFF/n91 , \UART_TXFF/n90 ,
         \UART_TXFF/n89 , \UART_TXFF/n88 , \UART_TXFF/n87 , \UART_TXFF/n86 ,
         \UART_TXFF/n85 , \UART_TXFF/n84 , \UART_TXFF/n83 , \UART_TXFF/n82 ,
         \UART_TXFF/n81 , \UART_TXFF/n80 , \UART_TXFF/n79 , \UART_TXFF/n78 ,
         \UART_TXFF/n77 , \UART_TXFF/n76 , \UART_TXFF/n75 , \UART_TXFF/n74 ,
         \UART_TXFF/n73 , \UART_TXFF/n72 , \UART_TXFF/n71 , \UART_TXFF/n70 ,
         \UART_TXFF/n69 , \UART_TXFF/n68 , \UART_TXFF/n67 , \UART_TXFF/n66 ,
         \UART_TXFF/n65 , \UART_TXFF/n64 , \UART_TXFF/n63 , \UART_TXFF/n62 ,
         \UART_TXFF/n61 , \UART_TXFF/n60 , \UART_TXFF/n59 , \UART_TXFF/n58 ,
         \UART_TXFF/n57 , \UART_TXFF/n56 , \UART_TXFF/n55 , \UART_TXFF/n54 ,
         \UART_TXFF/n53 , \UART_TXFF/n52 , \UART_TXFF/n51 , \UART_TXFF/n50 ,
         \UART_TXFF/n49 , \UART_TXFF/n48 , \UART_TXFF/n47 , \UART_TXFF/n46 ,
         \UART_TXFF/n45 , \UART_TXFF/n44 , \UART_TXFF/n43 , \UART_TXFF/n42 ,
         \UART_TXFF/n41 , \UART_TXFF/n40 , \UART_TXFF/n39 , \UART_TXFF/n38 ,
         \UART_TXFF/n37 , \UART_TXFF/n36 , \UART_TXFF/n35 , \UART_TXFF/n34 ,
         \UART_TXFF/n32 , \UART_TXFF/n31 , \UART_TXFF/n30 , \UART_TXFF/n29 ,
         \UART_TXFF/n28 , \UART_TXFF/n27 , \UART_TXFF/n26 , \UART_TXFF/n25 ,
         \UART_TXFF/n24 , \UART_TXFF/n23 , \UART_TXFF/n22 , \UART_TXFF/n21 ,
         \UART_TXFF/n20 , \UART_TXFF/n19 , \UART_TXFF/n18 , \UART_TXFF/n17 ,
         \UART_TXFF/n16 , \UART_TXFF/n15 , \UART_TXFF/n14 , \UART_TXFF/n13 ,
         \UART_TXFF/n12 , \UART_TXFF/n11 , \UART_TXFF/n10 , \UART_TXFF/n9 ,
         \UART_TXFF/n8 , \UART_TXFF/n7 , \UART_TXFF/n6 , \UART_TXFF/n5 ,
         \UART_TXFF/n4 , \UART_TXFF/n3 , \UART_TXFF/n2 , \UART_TXFF/n1 ,
         \UART_TXFF/n1817 , \UART_TXFF/n1816 , \UART_TXFF/n1815 ,
         \UART_TXFF/n1814 , \UART_TXFF/n1813 , \UART_TXFF/n1812 ,
         \UART_TXFF/n1811 , \UART_TXFF/n1810 , \UART_TXFF/n1809 ,
         \UART_TXFF/n1808 , \UART_TXFF/n1807 , \UART_TXFF/n1806 ,
         \UART_TXFF/n1805 , \UART_TXFF/n1804 , \UART_TXFF/n1803 ,
         \UART_TXFF/n1802 , \UART_TXFF/n1801 , \UART_TXFF/n1800 ,
         \UART_TXFF/n1799 , \UART_TXFF/n1798 , \UART_TXFF/n1797 ,
         \UART_TXFF/n1796 , \UART_TXFF/n1795 , \UART_TXFF/n1794 ,
         \UART_TXFF/n1793 , \UART_TXFF/n1792 , \UART_TXFF/n1791 ,
         \UART_TXFF/n1790 , \UART_TXFF/n1789 , \UART_TXFF/n1788 ,
         \UART_TXFF/n1787 , \UART_TXFF/n1786 , \UART_TXFF/n1785 ,
         \UART_TXFF/n1784 , \UART_TXFF/n1783 , \UART_TXFF/n1782 ,
         \UART_TXFF/n1781 , \UART_TXFF/n1780 , \UART_TXFF/n1779 ,
         \UART_TXFF/n1778 , \UART_TXFF/n1777 , \UART_TXFF/n1776 ,
         \UART_TXFF/n1775 , \UART_TXFF/n1774 , \UART_TXFF/n1773 ,
         \UART_TXFF/n1772 , \UART_TXFF/n1771 , \UART_TXFF/n1770 ,
         \UART_TXFF/n1769 , \UART_TXFF/n1768 , \UART_TXFF/n1767 ,
         \UART_TXFF/n1766 , \UART_TXFF/n1765 , \UART_TXFF/n1764 ,
         \UART_TXFF/n1763 , \UART_TXFF/n1762 , \UART_TXFF/n1761 ,
         \UART_TXFF/n1760 , \UART_TXFF/n1759 , \UART_TXFF/n1758 ,
         \UART_TXFF/n1757 , \UART_TXFF/n1756 , \UART_TXFF/n1755 ,
         \UART_TXFF/n1754 , \UART_TXFF/n1753 , \UART_TXFF/n1752 ,
         \UART_TXFF/n1751 , \UART_TXFF/n1750 , \UART_TXFF/n1749 ,
         \UART_TXFF/n1748 , \UART_TXFF/n1747 , \UART_TXFF/n1746 ,
         \UART_TXFF/n1745 , \UART_TXFF/n1744 , \UART_TXFF/n1743 ,
         \UART_TXFF/n1742 , \UART_TXFF/n1741 , \UART_TXFF/n1740 ,
         \UART_TXFF/n1739 , \UART_TXFF/n1738 , \UART_TXFF/n1737 ,
         \UART_TXFF/n1736 , \UART_TXFF/n1735 , \UART_TXFF/n1734 ,
         \UART_TXFF/n1733 , \UART_TXFF/n1732 , \UART_TXFF/n1731 ,
         \UART_TXFF/n1730 , \UART_TXFF/n1729 , \UART_TXFF/n1728 ,
         \UART_TXFF/n1727 , \UART_TXFF/n1726 , \UART_TXFF/n1725 ,
         \UART_TXFF/n1724 , \UART_TXFF/n1723 , \UART_TXFF/n1722 ,
         \UART_TXFF/n1721 , \UART_TXFF/n1720 , \UART_TXFF/n1719 ,
         \UART_TXFF/n1718 , \UART_TXFF/n1717 , \UART_TXFF/n1716 ,
         \UART_TXFF/n1715 , \UART_TXFF/n1714 , \UART_TXFF/n1713 ,
         \UART_TXFF/n1712 , \UART_TXFF/n1711 , \UART_TXFF/n1710 ,
         \UART_TXFF/n1709 , \UART_TXFF/n1708 , \UART_TXFF/n1707 ,
         \UART_TXFF/n1706 , \UART_TXFF/n1705 , \UART_TXFF/n1704 ,
         \UART_TXFF/n1703 , \UART_TXFF/n1702 , \UART_TXFF/n1701 ,
         \UART_TXFF/n1700 , \UART_TXFF/n1699 , \UART_TXFF/n1698 ,
         \UART_TXFF/n1697 , \UART_TXFF/n1696 , \UART_TXFF/n1695 ,
         \UART_TXFF/n1694 , \UART_TXFF/n1693 , \UART_TXFF/n1692 ,
         \UART_TXFF/n1691 , \UART_TXFF/n1690 , \UART_TXFF/n1689 ,
         \UART_TXFF/n1688 , \UART_TXFF/n1687 , \UART_TXFF/n1686 ,
         \UART_TXFF/n1685 , \UART_TXFF/n1684 , \UART_TXFF/n1683 ,
         \UART_TXFF/n1682 , \UART_TXFF/n1681 , \UART_TXFF/n1680 ,
         \UART_TXFF/n1679 , \UART_TXFF/n1678 , \UART_TXFF/n1677 ,
         \UART_TXFF/n1676 , \UART_TXFF/n1675 , \UART_TXFF/n1674 ,
         \UART_TXFF/n1673 , \UART_TXFF/n1672 , \UART_TXFF/n1671 ,
         \UART_TXFF/n1670 , \UART_TXFF/n1669 , \UART_TXFF/n1668 ,
         \UART_TXFF/n1667 , \UART_TXFF/n1666 , \UART_TXFF/n1665 ,
         \UART_TXFF/n1664 , \UART_TXFF/n1663 , \UART_TXFF/n1662 ,
         \UART_TXFF/n1661 , \UART_TXFF/n1660 , \UART_TXFF/n1659 ,
         \UART_TXFF/n1658 , \UART_TXFF/n1657 , \UART_TXFF/n1656 ,
         \UART_TXFF/n1655 , \UART_TXFF/n1654 , \UART_TXFF/n1653 ,
         \UART_TXFF/n1652 , \UART_TXFF/n1651 , \UART_TXFF/n1650 ,
         \UART_TXFF/n1649 , \UART_TXFF/n1648 , \UART_TXFF/n1647 ,
         \UART_TXFF/n1646 , \UART_TXFF/n1645 , \UART_TXFF/n1644 ,
         \UART_TXFF/n1643 , \UART_TXFF/n1642 , \UART_TXFF/n1641 ,
         \UART_TXFF/n1640 , \UART_TXFF/n1639 , \UART_TXFF/n1638 ,
         \UART_TXFF/n1637 , \UART_TXFF/n1636 , \UART_TXFF/n1635 ,
         \UART_TXFF/n1634 , \UART_TXFF/n1633 , \UART_TXFF/n1632 ,
         \UART_TXFF/n1631 , \UART_TXFF/n1630 , \UART_TXFF/n1629 ,
         \UART_TXFF/n1628 , \UART_TXFF/n1627 , \UART_TXFF/n1626 ,
         \UART_TXFF/n1625 , \UART_TXFF/n1624 , \UART_TXFF/n1623 ,
         \UART_TXFF/n1622 , \UART_TXFF/n1621 , \UART_TXFF/n1620 ,
         \UART_TXFF/n1619 , \UART_TXFF/n1618 , \UART_TXFF/n1617 ,
         \UART_TXFF/n1616 , \UART_TXFF/n1615 , \UART_TXFF/n1614 ,
         \UART_TXFF/n1613 , \UART_TXFF/n1612 , \UART_TXFF/n1611 ,
         \UART_TXFF/n1610 , \UART_TXFF/n1609 , \UART_TXFF/n1608 ,
         \UART_TXFF/n1607 , \UART_TXFF/n1606 , \UART_TXFF/n1605 ,
         \UART_TXFF/n1604 , \UART_TXFF/n1603 , \UART_TXFF/n1602 ,
         \UART_TXFF/n1601 , \UART_TXFF/n1600 , \UART_TXFF/n1599 ,
         \UART_TXFF/n1598 , \UART_TXFF/n1597 , \UART_TXFF/n1596 ,
         \UART_TXFF/n1595 , \UART_TXFF/n1594 , \UART_TXFF/n1593 ,
         \UART_TXFF/n1592 , \UART_TXFF/n1591 , \UART_TXFF/n1590 ,
         \UART_TXFF/n1589 , \UART_TXFF/n1588 , \UART_TXFF/n1587 ,
         \UART_TXFF/n1586 , \UART_TXFF/n1585 , \UART_TXFF/n1584 ,
         \UART_TXFF/n1583 , \UART_TXFF/n1582 , \UART_TXFF/n1581 ,
         \UART_TXFF/n1580 , \UART_TXFF/n1579 , \UART_TXFF/n1578 ,
         \UART_TXFF/n1577 , \UART_TXFF/n1576 , \UART_TXFF/n1575 ,
         \UART_TXFF/n1574 , \UART_TXFF/n1573 , \UART_TXFF/n1572 ,
         \UART_TXFF/n1571 , \UART_TXFF/n1570 , \UART_TXFF/n1569 ,
         \UART_TXFF/n1568 , \UART_TXFF/n1567 , \UART_TXFF/n1566 ,
         \UART_TXFF/n1565 , \UART_TXFF/n1564 , \UART_TXFF/n1563 ,
         \UART_TXFF/n1562 , \UART_TXFF/n1561 , \UART_TXFF/n1560 ,
         \UART_TXFF/n1559 , \UART_TXFF/n1558 , \UART_TXFF/n1557 ,
         \UART_TXFF/n1556 , \UART_TXFF/n1555 , \UART_TXFF/n1554 ,
         \UART_TXFF/n1553 , \UART_TXFF/n1552 , \UART_TXFF/n1551 ,
         \UART_TXFF/n1550 , \UART_TXFF/n1549 , \UART_TXFF/n1548 ,
         \UART_TXFF/n1547 , \UART_TXFF/n1546 , \UART_TXFF/n1545 ,
         \UART_TXFF/n1544 , \UART_TXFF/n1543 , \UART_TXFF/n1542 ,
         \UART_TXFF/n1541 , \UART_TXFF/n1540 , \UART_TXFF/n1539 ,
         \UART_TXFF/n1538 , \UART_TXFF/n1537 , \UART_TXFF/n1536 ,
         \UART_TXFF/n1535 , \UART_TXFF/n1534 , \UART_TXFF/n1533 ,
         \UART_TXFF/n1532 , \UART_TXFF/n1531 , \UART_TXFF/n1530 ,
         \UART_TXFF/n1529 , \UART_TXFF/n1528 , \UART_TXFF/n1527 ,
         \UART_TXFF/n1526 , \UART_TXFF/n1525 , \UART_TXFF/n1524 ,
         \UART_TXFF/n1523 , \UART_TXFF/n1522 , \UART_TXFF/n1521 ,
         \UART_TXFF/n1520 , \UART_TXFF/n1519 , \UART_TXFF/n1518 ,
         \UART_TXFF/n1517 , \UART_TXFF/n1516 , \UART_TXFF/n1515 ,
         \UART_TXFF/n1514 , \UART_TXFF/n1513 , \UART_TXFF/n1512 ,
         \UART_TXFF/n1511 , \UART_TXFF/n1510 , \UART_TXFF/n1509 ,
         \UART_TXFF/n1508 , \UART_TXFF/n1507 , \UART_TXFF/n1506 ,
         \UART_TXFF/n1505 , \UART_TXFF/n1504 , \UART_TXFF/n1503 ,
         \UART_TXFF/n1502 , \UART_TXFF/n1501 , \UART_TXFF/n1500 ,
         \UART_TXFF/n1499 , \UART_TXFF/n1498 , \UART_TXFF/n1497 ,
         \UART_TXFF/n1496 , \UART_TXFF/n1495 , \UART_TXFF/n1494 ,
         \UART_TXFF/n1493 , \UART_TXFF/n1492 , \UART_TXFF/n1491 ,
         \UART_TXFF/n1490 , \UART_TXFF/n1489 , \UART_TXFF/n1488 ,
         \UART_TXFF/n1487 , \UART_TXFF/n1486 , \UART_TXFF/n1485 ,
         \UART_TXFF/n1484 , \UART_TXFF/n1483 , \UART_TXFF/n1482 ,
         \UART_TXFF/n1481 , \UART_TXFF/n1480 , \UART_TXFF/n1479 ,
         \UART_TXFF/n1478 , \UART_TXFF/n1477 , \UART_TXFF/n1476 ,
         \UART_TXFF/n1475 , \UART_TXFF/n1474 , \UART_TXFF/n1473 ,
         \UART_TXFF/n1472 , \UART_TXFF/n1471 , \UART_TXFF/n1470 ,
         \UART_TXFF/n1469 , \UART_TXFF/n1468 , \UART_TXFF/n1467 ,
         \UART_TXFF/n1466 , \UART_TXFF/n1465 , \UART_TXFF/n1464 ,
         \UART_TXFF/n1463 , \UART_TXFF/n1462 , \UART_TXFF/n1461 ,
         \UART_TXFF/n1460 , \UART_TXFF/n1459 , \UART_TXFF/n1458 ,
         \UART_TXFF/n1457 , \UART_TXFF/n1456 , \UART_TXFF/n1455 ,
         \UART_TXFF/n1454 , \UART_TXFF/n1453 , \UART_TXFF/n1452 ,
         \UART_TXFF/n1451 , \UART_TXFF/n1450 , \UART_TXFF/n1449 ,
         \UART_TXFF/n1448 , \UART_TXFF/n1447 , \UART_TXFF/n1446 ,
         \UART_TXFF/n1445 , \UART_TXFF/n1444 , \UART_TXFF/n1443 ,
         \UART_TXFF/n1442 , \UART_TXFF/n1441 , \UART_TXFF/n1440 ,
         \UART_TXFF/n1439 , \UART_TXFF/n1438 , \UART_TXFF/n1437 ,
         \UART_TXFF/n1436 , \UART_TXFF/n1435 , \UART_TXFF/n1434 ,
         \UART_TXFF/n1433 , \UART_TXFF/n1432 , \UART_TXFF/n1431 ,
         \UART_TXFF/n1430 , \UART_TXFF/n1429 , \UART_TXFF/n1428 ,
         \UART_TXFF/n1427 , \UART_TXFF/n1426 , \UART_TXFF/n1425 ,
         \UART_TXFF/n1424 , \UART_TXFF/n1423 , \UART_TXFF/n1422 ,
         \UART_TXFF/n1421 , \UART_TXFF/n1420 , \UART_TXFF/n1419 ,
         \UART_TXFF/n1418 , \UART_TXFF/n1417 , \UART_TXFF/n1416 ,
         \UART_TXFF/n1415 , \UART_TXFF/n1414 , \UART_TXFF/n1413 ,
         \UART_TXFF/n1412 , \UART_TXFF/n1411 , \UART_TXFF/n1410 ,
         \UART_TXFF/n1409 , \UART_TXFF/n1408 , \UART_TXFF/n1407 ,
         \UART_TXFF/n1406 , \UART_TXFF/n1405 , \UART_TXFF/n1404 ,
         \UART_TXFF/n1403 , \UART_TXFF/n1402 , \UART_TXFF/n1401 ,
         \UART_TXFF/n1400 , \UART_TXFF/n1399 , \UART_TXFF/n1398 ,
         \UART_TXFF/n1397 , \UART_TXFF/n1396 , \UART_TXFF/n1395 ,
         \UART_TXFF/n1394 , \UART_TXFF/n1393 , \UART_TXFF/n1392 ,
         \UART_TXFF/n1391 , \UART_TXFF/n1390 , \UART_TXFF/n1389 ,
         \UART_TXFF/n1388 , \UART_TXFF/n1387 , \UART_TXFF/n1386 ,
         \UART_TXFF/n1385 , \UART_TXFF/n1384 , \UART_TXFF/n1383 ,
         \UART_TXFF/n1382 , \UART_TXFF/n1381 , \UART_TXFF/n1380 ,
         \UART_TXFF/n1379 , \UART_TXFF/n1378 , \UART_TXFF/n1377 ,
         \UART_TXFF/n1376 , \UART_TXFF/n1375 , \UART_TXFF/n1374 ,
         \UART_TXFF/n1373 , \UART_TXFF/n1372 , \UART_TXFF/n1371 ,
         \UART_TXFF/n1370 , \UART_TXFF/n1369 , \UART_TXFF/n1368 ,
         \UART_TXFF/n1367 , \UART_TXFF/n1366 , \UART_TXFF/n1365 ,
         \UART_TXFF/n1364 , \UART_TXFF/n1363 , \UART_TXFF/n1362 ,
         \UART_TXFF/n1361 , \UART_TXFF/n1360 , \UART_TXFF/n1359 ,
         \UART_TXFF/n1358 , \UART_TXFF/n1357 , \UART_TXFF/n1356 ,
         \UART_TXFF/n1355 , \UART_TXFF/n1354 , \UART_TXFF/n1353 ,
         \UART_TXFF/n1352 , \UART_TXFF/n1351 , \UART_TXFF/n1350 ,
         \UART_TXFF/n1349 , \UART_TXFF/n1348 , \UART_TXFF/n1347 ,
         \UART_TXFF/n1346 , \UART_TXFF/n1345 , \UART_TXFF/n1344 ,
         \UART_TXFF/n1343 , \UART_TXFF/n1342 , \UART_TXFF/n1341 ,
         \UART_TXFF/n1340 , \UART_TXFF/n1339 , \UART_TXFF/n1338 ,
         \UART_TXFF/n1337 , \UART_TXFF/n1336 , \UART_TXFF/n1335 ,
         \UART_TXFF/n1334 , \UART_TXFF/n1333 , \UART_TXFF/n1332 ,
         \UART_TXFF/n1331 , \UART_TXFF/n1330 , \UART_TXFF/n1329 ,
         \UART_TXFF/n1328 , \UART_TXFF/n1327 , \UART_TXFF/n1326 ,
         \UART_TXFF/n1325 , \UART_TXFF/n1324 , \UART_TXFF/n1323 ,
         \UART_TXFF/n1322 , \UART_TXFF/n1321 , \UART_TXFF/n1320 ,
         \UART_TXFF/n1319 , \UART_TXFF/n1318 , \UART_TXFF/n1317 ,
         \UART_TXFF/n1316 , \UART_TXFF/n1315 , \UART_TXFF/n1314 ,
         \UART_TXFF/n1313 , \UART_TXFF/n1312 , \UART_TXFF/n1311 ,
         \UART_TXFF/n1310 , \UART_TXFF/n1309 , \UART_TXFF/n1308 ,
         \UART_TXFF/n1307 , \UART_TXFF/n1306 , \UART_TXFF/n1305 ,
         \UART_TXFF/n1304 , \UART_TXFF/n1303 , \UART_TXFF/n1302 ,
         \UART_TXFF/n1301 , \UART_TXFF/n1300 , \UART_TXFF/n1299 ,
         \UART_TXFF/n1298 , \UART_TXFF/n1297 , \UART_TXFF/n1296 ,
         \UART_TXFF/n1295 , \UART_TXFF/n1294 , \UART_TXFF/n1293 ,
         \UART_TXFF/n1292 , \UART_TXFF/n1291 , \UART_TXFF/n1290 ,
         \UART_TXFF/n1289 , \UART_TXFF/n1288 , \UART_TXFF/n1287 ,
         \UART_TXFF/n772 , \UART_TXFF/n770 , \UART_TXFF/n768 ,
         \UART_TXFF/n766 , \UART_TXFF/n764 , \UART_TXFF/n762 ,
         \UART_TXFF/n760 , \UART_TXFF/n758 , \UART_TXFF/N130 ,
         \UART_TXFF/N129 , \UART_TXFF/N128 , \UART_TXFF/N127 ,
         \UART_TXFF/N126 , \UART_TXFF/N125 , \UART_TXFF/N124 ,
         \UART_TXFF/N123 , \UART_TXFF/iFIFOMem[0][0] ,
         \UART_TXFF/iFIFOMem[0][1] , \UART_TXFF/iFIFOMem[0][2] ,
         \UART_TXFF/iFIFOMem[0][3] , \UART_TXFF/iFIFOMem[0][4] ,
         \UART_TXFF/iFIFOMem[0][5] , \UART_TXFF/iFIFOMem[0][6] ,
         \UART_TXFF/iFIFOMem[0][7] , \UART_TXFF/iFIFOMem[1][0] ,
         \UART_TXFF/iFIFOMem[1][1] , \UART_TXFF/iFIFOMem[1][2] ,
         \UART_TXFF/iFIFOMem[1][3] , \UART_TXFF/iFIFOMem[1][4] ,
         \UART_TXFF/iFIFOMem[1][5] , \UART_TXFF/iFIFOMem[1][6] ,
         \UART_TXFF/iFIFOMem[1][7] , \UART_TXFF/iFIFOMem[2][0] ,
         \UART_TXFF/iFIFOMem[2][1] , \UART_TXFF/iFIFOMem[2][2] ,
         \UART_TXFF/iFIFOMem[2][3] , \UART_TXFF/iFIFOMem[2][4] ,
         \UART_TXFF/iFIFOMem[2][5] , \UART_TXFF/iFIFOMem[2][6] ,
         \UART_TXFF/iFIFOMem[2][7] , \UART_TXFF/iFIFOMem[3][0] ,
         \UART_TXFF/iFIFOMem[3][1] , \UART_TXFF/iFIFOMem[3][2] ,
         \UART_TXFF/iFIFOMem[3][3] , \UART_TXFF/iFIFOMem[3][4] ,
         \UART_TXFF/iFIFOMem[3][5] , \UART_TXFF/iFIFOMem[3][6] ,
         \UART_TXFF/iFIFOMem[3][7] , \UART_TXFF/iFIFOMem[4][0] ,
         \UART_TXFF/iFIFOMem[4][1] , \UART_TXFF/iFIFOMem[4][2] ,
         \UART_TXFF/iFIFOMem[4][3] , \UART_TXFF/iFIFOMem[4][4] ,
         \UART_TXFF/iFIFOMem[4][5] , \UART_TXFF/iFIFOMem[4][6] ,
         \UART_TXFF/iFIFOMem[4][7] , \UART_TXFF/iFIFOMem[5][0] ,
         \UART_TXFF/iFIFOMem[5][1] , \UART_TXFF/iFIFOMem[5][2] ,
         \UART_TXFF/iFIFOMem[5][3] , \UART_TXFF/iFIFOMem[5][4] ,
         \UART_TXFF/iFIFOMem[5][5] , \UART_TXFF/iFIFOMem[5][6] ,
         \UART_TXFF/iFIFOMem[5][7] , \UART_TXFF/iFIFOMem[6][0] ,
         \UART_TXFF/iFIFOMem[6][1] , \UART_TXFF/iFIFOMem[6][2] ,
         \UART_TXFF/iFIFOMem[6][3] , \UART_TXFF/iFIFOMem[6][4] ,
         \UART_TXFF/iFIFOMem[6][5] , \UART_TXFF/iFIFOMem[6][6] ,
         \UART_TXFF/iFIFOMem[6][7] , \UART_TXFF/iFIFOMem[7][0] ,
         \UART_TXFF/iFIFOMem[7][1] , \UART_TXFF/iFIFOMem[7][2] ,
         \UART_TXFF/iFIFOMem[7][3] , \UART_TXFF/iFIFOMem[7][4] ,
         \UART_TXFF/iFIFOMem[7][5] , \UART_TXFF/iFIFOMem[7][6] ,
         \UART_TXFF/iFIFOMem[7][7] , \UART_TXFF/iFIFOMem[8][0] ,
         \UART_TXFF/iFIFOMem[8][1] , \UART_TXFF/iFIFOMem[8][2] ,
         \UART_TXFF/iFIFOMem[8][3] , \UART_TXFF/iFIFOMem[8][4] ,
         \UART_TXFF/iFIFOMem[8][5] , \UART_TXFF/iFIFOMem[8][6] ,
         \UART_TXFF/iFIFOMem[8][7] , \UART_TXFF/iFIFOMem[9][0] ,
         \UART_TXFF/iFIFOMem[9][1] , \UART_TXFF/iFIFOMem[9][2] ,
         \UART_TXFF/iFIFOMem[9][3] , \UART_TXFF/iFIFOMem[9][4] ,
         \UART_TXFF/iFIFOMem[9][5] , \UART_TXFF/iFIFOMem[9][6] ,
         \UART_TXFF/iFIFOMem[9][7] , \UART_TXFF/iFIFOMem[10][0] ,
         \UART_TXFF/iFIFOMem[10][1] , \UART_TXFF/iFIFOMem[10][2] ,
         \UART_TXFF/iFIFOMem[10][3] , \UART_TXFF/iFIFOMem[10][4] ,
         \UART_TXFF/iFIFOMem[10][5] , \UART_TXFF/iFIFOMem[10][6] ,
         \UART_TXFF/iFIFOMem[10][7] , \UART_TXFF/iFIFOMem[11][0] ,
         \UART_TXFF/iFIFOMem[11][1] , \UART_TXFF/iFIFOMem[11][2] ,
         \UART_TXFF/iFIFOMem[11][3] , \UART_TXFF/iFIFOMem[11][4] ,
         \UART_TXFF/iFIFOMem[11][5] , \UART_TXFF/iFIFOMem[11][6] ,
         \UART_TXFF/iFIFOMem[11][7] , \UART_TXFF/iFIFOMem[12][0] ,
         \UART_TXFF/iFIFOMem[12][1] , \UART_TXFF/iFIFOMem[12][2] ,
         \UART_TXFF/iFIFOMem[12][3] , \UART_TXFF/iFIFOMem[12][4] ,
         \UART_TXFF/iFIFOMem[12][5] , \UART_TXFF/iFIFOMem[12][6] ,
         \UART_TXFF/iFIFOMem[12][7] , \UART_TXFF/iFIFOMem[13][0] ,
         \UART_TXFF/iFIFOMem[13][1] , \UART_TXFF/iFIFOMem[13][2] ,
         \UART_TXFF/iFIFOMem[13][3] , \UART_TXFF/iFIFOMem[13][4] ,
         \UART_TXFF/iFIFOMem[13][5] , \UART_TXFF/iFIFOMem[13][6] ,
         \UART_TXFF/iFIFOMem[13][7] , \UART_TXFF/iFIFOMem[14][0] ,
         \UART_TXFF/iFIFOMem[14][1] , \UART_TXFF/iFIFOMem[14][2] ,
         \UART_TXFF/iFIFOMem[14][3] , \UART_TXFF/iFIFOMem[14][4] ,
         \UART_TXFF/iFIFOMem[14][5] , \UART_TXFF/iFIFOMem[14][6] ,
         \UART_TXFF/iFIFOMem[14][7] , \UART_TXFF/iFIFOMem[15][0] ,
         \UART_TXFF/iFIFOMem[15][1] , \UART_TXFF/iFIFOMem[15][2] ,
         \UART_TXFF/iFIFOMem[15][3] , \UART_TXFF/iFIFOMem[15][4] ,
         \UART_TXFF/iFIFOMem[15][5] , \UART_TXFF/iFIFOMem[15][6] ,
         \UART_TXFF/iFIFOMem[15][7] , \UART_TXFF/iFIFOMem[16][0] ,
         \UART_TXFF/iFIFOMem[16][1] , \UART_TXFF/iFIFOMem[16][2] ,
         \UART_TXFF/iFIFOMem[16][3] , \UART_TXFF/iFIFOMem[16][4] ,
         \UART_TXFF/iFIFOMem[16][5] , \UART_TXFF/iFIFOMem[16][6] ,
         \UART_TXFF/iFIFOMem[16][7] , \UART_TXFF/iFIFOMem[17][0] ,
         \UART_TXFF/iFIFOMem[17][1] , \UART_TXFF/iFIFOMem[17][2] ,
         \UART_TXFF/iFIFOMem[17][3] , \UART_TXFF/iFIFOMem[17][4] ,
         \UART_TXFF/iFIFOMem[17][5] , \UART_TXFF/iFIFOMem[17][6] ,
         \UART_TXFF/iFIFOMem[17][7] , \UART_TXFF/iFIFOMem[18][0] ,
         \UART_TXFF/iFIFOMem[18][1] , \UART_TXFF/iFIFOMem[18][2] ,
         \UART_TXFF/iFIFOMem[18][3] , \UART_TXFF/iFIFOMem[18][4] ,
         \UART_TXFF/iFIFOMem[18][5] , \UART_TXFF/iFIFOMem[18][6] ,
         \UART_TXFF/iFIFOMem[18][7] , \UART_TXFF/iFIFOMem[19][0] ,
         \UART_TXFF/iFIFOMem[19][1] , \UART_TXFF/iFIFOMem[19][2] ,
         \UART_TXFF/iFIFOMem[19][3] , \UART_TXFF/iFIFOMem[19][4] ,
         \UART_TXFF/iFIFOMem[19][5] , \UART_TXFF/iFIFOMem[19][6] ,
         \UART_TXFF/iFIFOMem[19][7] , \UART_TXFF/iFIFOMem[20][0] ,
         \UART_TXFF/iFIFOMem[20][1] , \UART_TXFF/iFIFOMem[20][2] ,
         \UART_TXFF/iFIFOMem[20][3] , \UART_TXFF/iFIFOMem[20][4] ,
         \UART_TXFF/iFIFOMem[20][5] , \UART_TXFF/iFIFOMem[20][6] ,
         \UART_TXFF/iFIFOMem[20][7] , \UART_TXFF/iFIFOMem[21][0] ,
         \UART_TXFF/iFIFOMem[21][1] , \UART_TXFF/iFIFOMem[21][2] ,
         \UART_TXFF/iFIFOMem[21][3] , \UART_TXFF/iFIFOMem[21][4] ,
         \UART_TXFF/iFIFOMem[21][5] , \UART_TXFF/iFIFOMem[21][6] ,
         \UART_TXFF/iFIFOMem[21][7] , \UART_TXFF/iFIFOMem[22][0] ,
         \UART_TXFF/iFIFOMem[22][1] , \UART_TXFF/iFIFOMem[22][2] ,
         \UART_TXFF/iFIFOMem[22][3] , \UART_TXFF/iFIFOMem[22][4] ,
         \UART_TXFF/iFIFOMem[22][5] , \UART_TXFF/iFIFOMem[22][6] ,
         \UART_TXFF/iFIFOMem[22][7] , \UART_TXFF/iFIFOMem[23][0] ,
         \UART_TXFF/iFIFOMem[23][1] , \UART_TXFF/iFIFOMem[23][2] ,
         \UART_TXFF/iFIFOMem[23][3] , \UART_TXFF/iFIFOMem[23][4] ,
         \UART_TXFF/iFIFOMem[23][5] , \UART_TXFF/iFIFOMem[23][6] ,
         \UART_TXFF/iFIFOMem[23][7] , \UART_TXFF/iFIFOMem[24][0] ,
         \UART_TXFF/iFIFOMem[24][1] , \UART_TXFF/iFIFOMem[24][2] ,
         \UART_TXFF/iFIFOMem[24][3] , \UART_TXFF/iFIFOMem[24][4] ,
         \UART_TXFF/iFIFOMem[24][5] , \UART_TXFF/iFIFOMem[24][6] ,
         \UART_TXFF/iFIFOMem[24][7] , \UART_TXFF/iFIFOMem[25][0] ,
         \UART_TXFF/iFIFOMem[25][1] , \UART_TXFF/iFIFOMem[25][2] ,
         \UART_TXFF/iFIFOMem[25][3] , \UART_TXFF/iFIFOMem[25][4] ,
         \UART_TXFF/iFIFOMem[25][5] , \UART_TXFF/iFIFOMem[25][6] ,
         \UART_TXFF/iFIFOMem[25][7] , \UART_TXFF/iFIFOMem[26][0] ,
         \UART_TXFF/iFIFOMem[26][1] , \UART_TXFF/iFIFOMem[26][2] ,
         \UART_TXFF/iFIFOMem[26][3] , \UART_TXFF/iFIFOMem[26][4] ,
         \UART_TXFF/iFIFOMem[26][5] , \UART_TXFF/iFIFOMem[26][6] ,
         \UART_TXFF/iFIFOMem[26][7] , \UART_TXFF/iFIFOMem[27][0] ,
         \UART_TXFF/iFIFOMem[27][1] , \UART_TXFF/iFIFOMem[27][2] ,
         \UART_TXFF/iFIFOMem[27][3] , \UART_TXFF/iFIFOMem[27][4] ,
         \UART_TXFF/iFIFOMem[27][5] , \UART_TXFF/iFIFOMem[27][6] ,
         \UART_TXFF/iFIFOMem[27][7] , \UART_TXFF/iFIFOMem[28][0] ,
         \UART_TXFF/iFIFOMem[28][1] , \UART_TXFF/iFIFOMem[28][2] ,
         \UART_TXFF/iFIFOMem[28][3] , \UART_TXFF/iFIFOMem[28][4] ,
         \UART_TXFF/iFIFOMem[28][5] , \UART_TXFF/iFIFOMem[28][6] ,
         \UART_TXFF/iFIFOMem[28][7] , \UART_TXFF/iFIFOMem[29][0] ,
         \UART_TXFF/iFIFOMem[29][1] , \UART_TXFF/iFIFOMem[29][2] ,
         \UART_TXFF/iFIFOMem[29][3] , \UART_TXFF/iFIFOMem[29][4] ,
         \UART_TXFF/iFIFOMem[29][5] , \UART_TXFF/iFIFOMem[29][6] ,
         \UART_TXFF/iFIFOMem[29][7] , \UART_TXFF/iFIFOMem[30][0] ,
         \UART_TXFF/iFIFOMem[30][1] , \UART_TXFF/iFIFOMem[30][2] ,
         \UART_TXFF/iFIFOMem[30][3] , \UART_TXFF/iFIFOMem[30][4] ,
         \UART_TXFF/iFIFOMem[30][5] , \UART_TXFF/iFIFOMem[30][6] ,
         \UART_TXFF/iFIFOMem[30][7] , \UART_TXFF/iFIFOMem[31][0] ,
         \UART_TXFF/iFIFOMem[31][1] , \UART_TXFF/iFIFOMem[31][2] ,
         \UART_TXFF/iFIFOMem[31][3] , \UART_TXFF/iFIFOMem[31][4] ,
         \UART_TXFF/iFIFOMem[31][5] , \UART_TXFF/iFIFOMem[31][6] ,
         \UART_TXFF/iFIFOMem[31][7] , \UART_TXFF/iFIFOMem[32][0] ,
         \UART_TXFF/iFIFOMem[32][1] , \UART_TXFF/iFIFOMem[32][2] ,
         \UART_TXFF/iFIFOMem[32][3] , \UART_TXFF/iFIFOMem[32][4] ,
         \UART_TXFF/iFIFOMem[32][5] , \UART_TXFF/iFIFOMem[32][6] ,
         \UART_TXFF/iFIFOMem[32][7] , \UART_TXFF/iFIFOMem[33][0] ,
         \UART_TXFF/iFIFOMem[33][1] , \UART_TXFF/iFIFOMem[33][2] ,
         \UART_TXFF/iFIFOMem[33][3] , \UART_TXFF/iFIFOMem[33][4] ,
         \UART_TXFF/iFIFOMem[33][5] , \UART_TXFF/iFIFOMem[33][6] ,
         \UART_TXFF/iFIFOMem[33][7] , \UART_TXFF/iFIFOMem[34][0] ,
         \UART_TXFF/iFIFOMem[34][1] , \UART_TXFF/iFIFOMem[34][2] ,
         \UART_TXFF/iFIFOMem[34][3] , \UART_TXFF/iFIFOMem[34][4] ,
         \UART_TXFF/iFIFOMem[34][5] , \UART_TXFF/iFIFOMem[34][6] ,
         \UART_TXFF/iFIFOMem[34][7] , \UART_TXFF/iFIFOMem[35][0] ,
         \UART_TXFF/iFIFOMem[35][1] , \UART_TXFF/iFIFOMem[35][2] ,
         \UART_TXFF/iFIFOMem[35][3] , \UART_TXFF/iFIFOMem[35][4] ,
         \UART_TXFF/iFIFOMem[35][5] , \UART_TXFF/iFIFOMem[35][6] ,
         \UART_TXFF/iFIFOMem[35][7] , \UART_TXFF/iFIFOMem[36][0] ,
         \UART_TXFF/iFIFOMem[36][1] , \UART_TXFF/iFIFOMem[36][2] ,
         \UART_TXFF/iFIFOMem[36][3] , \UART_TXFF/iFIFOMem[36][4] ,
         \UART_TXFF/iFIFOMem[36][5] , \UART_TXFF/iFIFOMem[36][6] ,
         \UART_TXFF/iFIFOMem[36][7] , \UART_TXFF/iFIFOMem[37][0] ,
         \UART_TXFF/iFIFOMem[37][1] , \UART_TXFF/iFIFOMem[37][2] ,
         \UART_TXFF/iFIFOMem[37][3] , \UART_TXFF/iFIFOMem[37][4] ,
         \UART_TXFF/iFIFOMem[37][5] , \UART_TXFF/iFIFOMem[37][6] ,
         \UART_TXFF/iFIFOMem[37][7] , \UART_TXFF/iFIFOMem[38][0] ,
         \UART_TXFF/iFIFOMem[38][1] , \UART_TXFF/iFIFOMem[38][2] ,
         \UART_TXFF/iFIFOMem[38][3] , \UART_TXFF/iFIFOMem[38][4] ,
         \UART_TXFF/iFIFOMem[38][5] , \UART_TXFF/iFIFOMem[38][6] ,
         \UART_TXFF/iFIFOMem[38][7] , \UART_TXFF/iFIFOMem[39][0] ,
         \UART_TXFF/iFIFOMem[39][1] , \UART_TXFF/iFIFOMem[39][2] ,
         \UART_TXFF/iFIFOMem[39][3] , \UART_TXFF/iFIFOMem[39][4] ,
         \UART_TXFF/iFIFOMem[39][5] , \UART_TXFF/iFIFOMem[39][6] ,
         \UART_TXFF/iFIFOMem[39][7] , \UART_TXFF/iFIFOMem[40][0] ,
         \UART_TXFF/iFIFOMem[40][1] , \UART_TXFF/iFIFOMem[40][2] ,
         \UART_TXFF/iFIFOMem[40][3] , \UART_TXFF/iFIFOMem[40][4] ,
         \UART_TXFF/iFIFOMem[40][5] , \UART_TXFF/iFIFOMem[40][6] ,
         \UART_TXFF/iFIFOMem[40][7] , \UART_TXFF/iFIFOMem[41][0] ,
         \UART_TXFF/iFIFOMem[41][1] , \UART_TXFF/iFIFOMem[41][2] ,
         \UART_TXFF/iFIFOMem[41][3] , \UART_TXFF/iFIFOMem[41][4] ,
         \UART_TXFF/iFIFOMem[41][5] , \UART_TXFF/iFIFOMem[41][6] ,
         \UART_TXFF/iFIFOMem[41][7] , \UART_TXFF/iFIFOMem[42][0] ,
         \UART_TXFF/iFIFOMem[42][1] , \UART_TXFF/iFIFOMem[42][2] ,
         \UART_TXFF/iFIFOMem[42][3] , \UART_TXFF/iFIFOMem[42][4] ,
         \UART_TXFF/iFIFOMem[42][5] , \UART_TXFF/iFIFOMem[42][6] ,
         \UART_TXFF/iFIFOMem[42][7] , \UART_TXFF/iFIFOMem[43][0] ,
         \UART_TXFF/iFIFOMem[43][1] , \UART_TXFF/iFIFOMem[43][2] ,
         \UART_TXFF/iFIFOMem[43][3] , \UART_TXFF/iFIFOMem[43][4] ,
         \UART_TXFF/iFIFOMem[43][5] , \UART_TXFF/iFIFOMem[43][6] ,
         \UART_TXFF/iFIFOMem[43][7] , \UART_TXFF/iFIFOMem[44][0] ,
         \UART_TXFF/iFIFOMem[44][1] , \UART_TXFF/iFIFOMem[44][2] ,
         \UART_TXFF/iFIFOMem[44][3] , \UART_TXFF/iFIFOMem[44][4] ,
         \UART_TXFF/iFIFOMem[44][5] , \UART_TXFF/iFIFOMem[44][6] ,
         \UART_TXFF/iFIFOMem[44][7] , \UART_TXFF/iFIFOMem[45][0] ,
         \UART_TXFF/iFIFOMem[45][1] , \UART_TXFF/iFIFOMem[45][2] ,
         \UART_TXFF/iFIFOMem[45][3] , \UART_TXFF/iFIFOMem[45][4] ,
         \UART_TXFF/iFIFOMem[45][5] , \UART_TXFF/iFIFOMem[45][6] ,
         \UART_TXFF/iFIFOMem[45][7] , \UART_TXFF/iFIFOMem[46][0] ,
         \UART_TXFF/iFIFOMem[46][1] , \UART_TXFF/iFIFOMem[46][2] ,
         \UART_TXFF/iFIFOMem[46][3] , \UART_TXFF/iFIFOMem[46][4] ,
         \UART_TXFF/iFIFOMem[46][5] , \UART_TXFF/iFIFOMem[46][6] ,
         \UART_TXFF/iFIFOMem[46][7] , \UART_TXFF/iFIFOMem[47][0] ,
         \UART_TXFF/iFIFOMem[47][1] , \UART_TXFF/iFIFOMem[47][2] ,
         \UART_TXFF/iFIFOMem[47][3] , \UART_TXFF/iFIFOMem[47][4] ,
         \UART_TXFF/iFIFOMem[47][5] , \UART_TXFF/iFIFOMem[47][6] ,
         \UART_TXFF/iFIFOMem[47][7] , \UART_TXFF/iFIFOMem[48][0] ,
         \UART_TXFF/iFIFOMem[48][1] , \UART_TXFF/iFIFOMem[48][2] ,
         \UART_TXFF/iFIFOMem[48][3] , \UART_TXFF/iFIFOMem[48][4] ,
         \UART_TXFF/iFIFOMem[48][5] , \UART_TXFF/iFIFOMem[48][6] ,
         \UART_TXFF/iFIFOMem[48][7] , \UART_TXFF/iFIFOMem[49][0] ,
         \UART_TXFF/iFIFOMem[49][1] , \UART_TXFF/iFIFOMem[49][2] ,
         \UART_TXFF/iFIFOMem[49][3] , \UART_TXFF/iFIFOMem[49][4] ,
         \UART_TXFF/iFIFOMem[49][5] , \UART_TXFF/iFIFOMem[49][6] ,
         \UART_TXFF/iFIFOMem[49][7] , \UART_TXFF/iFIFOMem[50][0] ,
         \UART_TXFF/iFIFOMem[50][1] , \UART_TXFF/iFIFOMem[50][2] ,
         \UART_TXFF/iFIFOMem[50][3] , \UART_TXFF/iFIFOMem[50][4] ,
         \UART_TXFF/iFIFOMem[50][5] , \UART_TXFF/iFIFOMem[50][6] ,
         \UART_TXFF/iFIFOMem[50][7] , \UART_TXFF/iFIFOMem[51][0] ,
         \UART_TXFF/iFIFOMem[51][1] , \UART_TXFF/iFIFOMem[51][2] ,
         \UART_TXFF/iFIFOMem[51][3] , \UART_TXFF/iFIFOMem[51][4] ,
         \UART_TXFF/iFIFOMem[51][5] , \UART_TXFF/iFIFOMem[51][6] ,
         \UART_TXFF/iFIFOMem[51][7] , \UART_TXFF/iFIFOMem[52][0] ,
         \UART_TXFF/iFIFOMem[52][1] , \UART_TXFF/iFIFOMem[52][2] ,
         \UART_TXFF/iFIFOMem[52][3] , \UART_TXFF/iFIFOMem[52][4] ,
         \UART_TXFF/iFIFOMem[52][5] , \UART_TXFF/iFIFOMem[52][6] ,
         \UART_TXFF/iFIFOMem[52][7] , \UART_TXFF/iFIFOMem[53][0] ,
         \UART_TXFF/iFIFOMem[53][1] , \UART_TXFF/iFIFOMem[53][2] ,
         \UART_TXFF/iFIFOMem[53][3] , \UART_TXFF/iFIFOMem[53][4] ,
         \UART_TXFF/iFIFOMem[53][5] , \UART_TXFF/iFIFOMem[53][6] ,
         \UART_TXFF/iFIFOMem[53][7] , \UART_TXFF/iFIFOMem[54][0] ,
         \UART_TXFF/iFIFOMem[54][1] , \UART_TXFF/iFIFOMem[54][2] ,
         \UART_TXFF/iFIFOMem[54][3] , \UART_TXFF/iFIFOMem[54][4] ,
         \UART_TXFF/iFIFOMem[54][5] , \UART_TXFF/iFIFOMem[54][6] ,
         \UART_TXFF/iFIFOMem[54][7] , \UART_TXFF/iFIFOMem[55][0] ,
         \UART_TXFF/iFIFOMem[55][1] , \UART_TXFF/iFIFOMem[55][2] ,
         \UART_TXFF/iFIFOMem[55][3] , \UART_TXFF/iFIFOMem[55][4] ,
         \UART_TXFF/iFIFOMem[55][5] , \UART_TXFF/iFIFOMem[55][6] ,
         \UART_TXFF/iFIFOMem[55][7] , \UART_TXFF/iFIFOMem[56][0] ,
         \UART_TXFF/iFIFOMem[56][1] , \UART_TXFF/iFIFOMem[56][2] ,
         \UART_TXFF/iFIFOMem[56][3] , \UART_TXFF/iFIFOMem[56][4] ,
         \UART_TXFF/iFIFOMem[56][5] , \UART_TXFF/iFIFOMem[56][6] ,
         \UART_TXFF/iFIFOMem[56][7] , \UART_TXFF/iFIFOMem[57][0] ,
         \UART_TXFF/iFIFOMem[57][1] , \UART_TXFF/iFIFOMem[57][2] ,
         \UART_TXFF/iFIFOMem[57][3] , \UART_TXFF/iFIFOMem[57][4] ,
         \UART_TXFF/iFIFOMem[57][5] , \UART_TXFF/iFIFOMem[57][6] ,
         \UART_TXFF/iFIFOMem[57][7] , \UART_TXFF/iFIFOMem[58][0] ,
         \UART_TXFF/iFIFOMem[58][1] , \UART_TXFF/iFIFOMem[58][2] ,
         \UART_TXFF/iFIFOMem[58][3] , \UART_TXFF/iFIFOMem[58][4] ,
         \UART_TXFF/iFIFOMem[58][5] , \UART_TXFF/iFIFOMem[58][6] ,
         \UART_TXFF/iFIFOMem[58][7] , \UART_TXFF/iFIFOMem[59][0] ,
         \UART_TXFF/iFIFOMem[59][1] , \UART_TXFF/iFIFOMem[59][2] ,
         \UART_TXFF/iFIFOMem[59][3] , \UART_TXFF/iFIFOMem[59][4] ,
         \UART_TXFF/iFIFOMem[59][5] , \UART_TXFF/iFIFOMem[59][6] ,
         \UART_TXFF/iFIFOMem[59][7] , \UART_TXFF/iFIFOMem[60][0] ,
         \UART_TXFF/iFIFOMem[60][1] , \UART_TXFF/iFIFOMem[60][2] ,
         \UART_TXFF/iFIFOMem[60][3] , \UART_TXFF/iFIFOMem[60][4] ,
         \UART_TXFF/iFIFOMem[60][5] , \UART_TXFF/iFIFOMem[60][6] ,
         \UART_TXFF/iFIFOMem[60][7] , \UART_TXFF/iFIFOMem[61][0] ,
         \UART_TXFF/iFIFOMem[61][1] , \UART_TXFF/iFIFOMem[61][2] ,
         \UART_TXFF/iFIFOMem[61][3] , \UART_TXFF/iFIFOMem[61][4] ,
         \UART_TXFF/iFIFOMem[61][5] , \UART_TXFF/iFIFOMem[61][6] ,
         \UART_TXFF/iFIFOMem[61][7] , \UART_TXFF/iFIFOMem[62][0] ,
         \UART_TXFF/iFIFOMem[62][1] , \UART_TXFF/iFIFOMem[62][2] ,
         \UART_TXFF/iFIFOMem[62][3] , \UART_TXFF/iFIFOMem[62][4] ,
         \UART_TXFF/iFIFOMem[62][5] , \UART_TXFF/iFIFOMem[62][6] ,
         \UART_TXFF/iFIFOMem[62][7] , \UART_TXFF/iFIFOMem[63][0] ,
         \UART_TXFF/iFIFOMem[63][1] , \UART_TXFF/iFIFOMem[63][2] ,
         \UART_TXFF/iFIFOMem[63][3] , \UART_TXFF/iFIFOMem[63][4] ,
         \UART_TXFF/iFIFOMem[63][5] , \UART_TXFF/iFIFOMem[63][6] ,
         \UART_TXFF/iFIFOMem[63][7] , \UART_TXFF/N56 , \UART_TXFF/N38 ,
         \UART_TXFF/N37 , \UART_TXFF/N36 , \UART_TXFF/N35 , \UART_TXFF/N34 ,
         \UART_TXFF/N33 , \UART_TXFF/N30 , \UART_TXFF/N29 , \UART_TXFF/N28 ,
         \UART_TXFF/N27 , \UART_TXFF/N26 , \UART_TXFF/N25 ,
         \UART_TXFF/iWRAddr[0] , \UART_TXFF/iWRAddr[1] ,
         \UART_TXFF/iWRAddr[2] , \UART_TXFF/iWRAddr[3] ,
         \UART_TXFF/iWRAddr[4] , \UART_TXFF/iWRAddr[5] ,
         \UART_TXFF/iWRAddr[6] , \UART_TXFF/iRDAddr[6] , \UART_TXFF/USAGE[0] ,
         \UART_TXFF/USAGE[1] , \UART_TXFF/USAGE[2] , \UART_TXFF/USAGE[3] ,
         \UART_TXFF/N17 , \UART_TXFF/N16 , \UART_TXFF/N15 , \UART_TXFF/N14 ,
         \UART_TXFF/N13 , \UART_TXFF/N12 , \UART_RXFF/n451 , \UART_RXFF/n450 ,
         \UART_RXFF/n449 , \UART_RXFF/n448 , \UART_RXFF/n447 ,
         \UART_RXFF/n446 , \UART_RXFF/n445 , \UART_RXFF/n444 ,
         \UART_RXFF/n443 , \UART_RXFF/n442 , \UART_RXFF/n441 ,
         \UART_RXFF/n440 , \UART_RXFF/n439 , \UART_RXFF/n438 ,
         \UART_RXFF/n437 , \UART_RXFF/n436 , \UART_RXFF/n435 ,
         \UART_RXFF/n434 , \UART_RXFF/n433 , \UART_RXFF/n432 ,
         \UART_RXFF/n431 , \UART_RXFF/n430 , \UART_RXFF/n429 ,
         \UART_RXFF/n428 , \UART_RXFF/n427 , \UART_RXFF/n426 ,
         \UART_RXFF/n425 , \UART_RXFF/n424 , \UART_RXFF/n423 ,
         \UART_RXFF/n422 , \UART_RXFF/n421 , \UART_RXFF/n420 ,
         \UART_RXFF/n419 , \UART_RXFF/n418 , \UART_RXFF/n417 ,
         \UART_RXFF/n416 , \UART_RXFF/n415 , \UART_RXFF/n414 ,
         \UART_RXFF/n413 , \UART_RXFF/n412 , \UART_RXFF/n411 ,
         \UART_RXFF/n410 , \UART_RXFF/n409 , \UART_RXFF/n408 ,
         \UART_RXFF/n407 , \UART_RXFF/n406 , \UART_RXFF/n405 ,
         \UART_RXFF/n404 , \UART_RXFF/n403 , \UART_RXFF/n402 ,
         \UART_RXFF/n401 , \UART_RXFF/n400 , \UART_RXFF/n399 ,
         \UART_RXFF/n398 , \UART_RXFF/n397 , \UART_RXFF/n396 ,
         \UART_RXFF/n395 , \UART_RXFF/n394 , \UART_RXFF/n393 ,
         \UART_RXFF/n392 , \UART_RXFF/n391 , \UART_RXFF/n390 ,
         \UART_RXFF/n389 , \UART_RXFF/n388 , \UART_RXFF/n387 ,
         \UART_RXFF/n386 , \UART_RXFF/n385 , \UART_RXFF/n384 ,
         \UART_RXFF/n383 , \UART_RXFF/n382 , \UART_RXFF/n381 ,
         \UART_RXFF/n380 , \UART_RXFF/n379 , \UART_RXFF/n378 ,
         \UART_RXFF/n377 , \UART_RXFF/n376 , \UART_RXFF/n375 ,
         \UART_RXFF/n374 , \UART_RXFF/n373 , \UART_RXFF/n372 ,
         \UART_RXFF/n371 , \UART_RXFF/n370 , \UART_RXFF/n369 ,
         \UART_RXFF/n368 , \UART_RXFF/n367 , \UART_RXFF/n366 ,
         \UART_RXFF/n365 , \UART_RXFF/n364 , \UART_RXFF/n363 ,
         \UART_RXFF/n362 , \UART_RXFF/n361 , \UART_RXFF/n360 ,
         \UART_RXFF/n359 , \UART_RXFF/n358 , \UART_RXFF/n357 ,
         \UART_RXFF/n356 , \UART_RXFF/n355 , \UART_RXFF/n354 ,
         \UART_RXFF/n353 , \UART_RXFF/n352 , \UART_RXFF/n351 ,
         \UART_RXFF/n350 , \UART_RXFF/n349 , \UART_RXFF/n348 ,
         \UART_RXFF/n347 , \UART_RXFF/n346 , \UART_RXFF/n345 ,
         \UART_RXFF/n344 , \UART_RXFF/n343 , \UART_RXFF/n342 ,
         \UART_RXFF/n341 , \UART_RXFF/n340 , \UART_RXFF/n339 ,
         \UART_RXFF/n338 , \UART_RXFF/n337 , \UART_RXFF/n336 ,
         \UART_RXFF/n335 , \UART_RXFF/n334 , \UART_RXFF/n333 ,
         \UART_RXFF/n332 , \UART_RXFF/n331 , \UART_RXFF/n330 ,
         \UART_RXFF/n329 , \UART_RXFF/n328 , \UART_RXFF/n327 ,
         \UART_RXFF/n326 , \UART_RXFF/n325 , \UART_RXFF/n324 ,
         \UART_RXFF/n323 , \UART_RXFF/n322 , \UART_RXFF/n321 ,
         \UART_RXFF/n320 , \UART_RXFF/n318 , \UART_RXFF/n317 ,
         \UART_RXFF/n316 , \UART_RXFF/n315 , \UART_RXFF/n314 ,
         \UART_RXFF/n313 , \UART_RXFF/n312 , \UART_RXFF/n311 ,
         \UART_RXFF/n310 , \UART_RXFF/n309 , \UART_RXFF/n308 ,
         \UART_RXFF/n307 , \UART_RXFF/n306 , \UART_RXFF/n305 ,
         \UART_RXFF/n304 , \UART_RXFF/n303 , \UART_RXFF/n302 ,
         \UART_RXFF/n301 , \UART_RXFF/n300 , \UART_RXFF/n299 ,
         \UART_RXFF/n298 , \UART_RXFF/n297 , \UART_RXFF/n296 ,
         \UART_RXFF/n295 , \UART_RXFF/n294 , \UART_RXFF/n293 ,
         \UART_RXFF/n292 , \UART_RXFF/n291 , \UART_RXFF/n290 ,
         \UART_RXFF/n289 , \UART_RXFF/n288 , \UART_RXFF/n287 ,
         \UART_RXFF/n286 , \UART_RXFF/n285 , \UART_RXFF/n284 ,
         \UART_RXFF/n283 , \UART_RXFF/n282 , \UART_RXFF/n281 ,
         \UART_RXFF/n280 , \UART_RXFF/n279 , \UART_RXFF/n278 ,
         \UART_RXFF/n277 , \UART_RXFF/n276 , \UART_RXFF/n275 ,
         \UART_RXFF/n274 , \UART_RXFF/n273 , \UART_RXFF/n272 ,
         \UART_RXFF/n271 , \UART_RXFF/n270 , \UART_RXFF/n269 ,
         \UART_RXFF/n268 , \UART_RXFF/n267 , \UART_RXFF/n266 ,
         \UART_RXFF/n265 , \UART_RXFF/n264 , \UART_RXFF/n263 ,
         \UART_RXFF/n262 , \UART_RXFF/n261 , \UART_RXFF/n260 ,
         \UART_RXFF/n259 , \UART_RXFF/n258 , \UART_RXFF/n257 ,
         \UART_RXFF/n256 , \UART_RXFF/n255 , \UART_RXFF/n254 ,
         \UART_RXFF/n253 , \UART_RXFF/n252 , \UART_RXFF/n251 ,
         \UART_RXFF/n250 , \UART_RXFF/n249 , \UART_RXFF/n248 ,
         \UART_RXFF/n247 , \UART_RXFF/n246 , \UART_RXFF/n245 ,
         \UART_RXFF/n244 , \UART_RXFF/n243 , \UART_RXFF/n242 ,
         \UART_RXFF/n241 , \UART_RXFF/n240 , \UART_RXFF/n239 ,
         \UART_RXFF/n238 , \UART_RXFF/n237 , \UART_RXFF/n236 ,
         \UART_RXFF/n235 , \UART_RXFF/n234 , \UART_RXFF/n233 ,
         \UART_RXFF/n232 , \UART_RXFF/n231 , \UART_RXFF/n230 ,
         \UART_RXFF/n229 , \UART_RXFF/n228 , \UART_RXFF/n227 ,
         \UART_RXFF/n226 , \UART_RXFF/n225 , \UART_RXFF/n224 ,
         \UART_RXFF/n223 , \UART_RXFF/n222 , \UART_RXFF/n221 ,
         \UART_RXFF/n220 , \UART_RXFF/n219 , \UART_RXFF/n218 ,
         \UART_RXFF/n217 , \UART_RXFF/n216 , \UART_RXFF/n215 ,
         \UART_RXFF/n214 , \UART_RXFF/n213 , \UART_RXFF/n212 ,
         \UART_RXFF/n211 , \UART_RXFF/n210 , \UART_RXFF/n209 ,
         \UART_RXFF/n208 , \UART_RXFF/n207 , \UART_RXFF/n206 ,
         \UART_RXFF/n205 , \UART_RXFF/n204 , \UART_RXFF/n203 ,
         \UART_RXFF/n202 , \UART_RXFF/n201 , \UART_RXFF/n200 ,
         \UART_RXFF/n199 , \UART_RXFF/n198 , \UART_RXFF/n197 ,
         \UART_RXFF/n196 , \UART_RXFF/n195 , \UART_RXFF/n194 ,
         \UART_RXFF/n193 , \UART_RXFF/n192 , \UART_RXFF/n191 ,
         \UART_RXFF/n190 , \UART_RXFF/n189 , \UART_RXFF/n188 ,
         \UART_RXFF/n187 , \UART_RXFF/n186 , \UART_RXFF/n185 ,
         \UART_RXFF/n184 , \UART_RXFF/n183 , \UART_RXFF/n182 ,
         \UART_RXFF/n181 , \UART_RXFF/n180 , \UART_RXFF/n179 ,
         \UART_RXFF/n178 , \UART_RXFF/n177 , \UART_RXFF/n176 ,
         \UART_RXFF/n175 , \UART_RXFF/n174 , \UART_RXFF/n173 ,
         \UART_RXFF/n172 , \UART_RXFF/n171 , \UART_RXFF/n170 ,
         \UART_RXFF/n169 , \UART_RXFF/n168 , \UART_RXFF/n167 ,
         \UART_RXFF/n166 , \UART_RXFF/n165 , \UART_RXFF/n164 ,
         \UART_RXFF/n163 , \UART_RXFF/n162 , \UART_RXFF/n161 ,
         \UART_RXFF/n160 , \UART_RXFF/n159 , \UART_RXFF/n158 ,
         \UART_RXFF/n157 , \UART_RXFF/n156 , \UART_RXFF/n155 ,
         \UART_RXFF/n154 , \UART_RXFF/n153 , \UART_RXFF/n152 ,
         \UART_RXFF/n151 , \UART_RXFF/n150 , \UART_RXFF/n149 ,
         \UART_RXFF/n148 , \UART_RXFF/n147 , \UART_RXFF/n146 ,
         \UART_RXFF/n145 , \UART_RXFF/n144 , \UART_RXFF/n143 ,
         \UART_RXFF/n142 , \UART_RXFF/n141 , \UART_RXFF/n140 ,
         \UART_RXFF/n139 , \UART_RXFF/n138 , \UART_RXFF/n137 ,
         \UART_RXFF/n136 , \UART_RXFF/n135 , \UART_RXFF/n134 ,
         \UART_RXFF/n133 , \UART_RXFF/n132 , \UART_RXFF/n131 ,
         \UART_RXFF/n130 , \UART_RXFF/n129 , \UART_RXFF/n128 ,
         \UART_RXFF/n127 , \UART_RXFF/n126 , \UART_RXFF/n125 ,
         \UART_RXFF/n124 , \UART_RXFF/n123 , \UART_RXFF/n122 ,
         \UART_RXFF/n121 , \UART_RXFF/n120 , \UART_RXFF/n119 ,
         \UART_RXFF/n118 , \UART_RXFF/n117 , \UART_RXFF/n116 ,
         \UART_RXFF/n115 , \UART_RXFF/n114 , \UART_RXFF/n113 ,
         \UART_RXFF/n112 , \UART_RXFF/n111 , \UART_RXFF/n110 ,
         \UART_RXFF/n109 , \UART_RXFF/n108 , \UART_RXFF/n107 ,
         \UART_RXFF/n106 , \UART_RXFF/n105 , \UART_RXFF/n104 ,
         \UART_RXFF/n103 , \UART_RXFF/n102 , \UART_RXFF/n101 ,
         \UART_RXFF/n100 , \UART_RXFF/n99 , \UART_RXFF/n98 , \UART_RXFF/n97 ,
         \UART_RXFF/n96 , \UART_RXFF/n95 , \UART_RXFF/n94 , \UART_RXFF/n93 ,
         \UART_RXFF/n92 , \UART_RXFF/n91 , \UART_RXFF/n90 , \UART_RXFF/n89 ,
         \UART_RXFF/n88 , \UART_RXFF/n87 , \UART_RXFF/n86 , \UART_RXFF/n85 ,
         \UART_RXFF/n84 , \UART_RXFF/n83 , \UART_RXFF/n82 , \UART_RXFF/n81 ,
         \UART_RXFF/n80 , \UART_RXFF/n79 , \UART_RXFF/n78 , \UART_RXFF/n77 ,
         \UART_RXFF/n76 , \UART_RXFF/n75 , \UART_RXFF/n74 , \UART_RXFF/n73 ,
         \UART_RXFF/n72 , \UART_RXFF/n71 , \UART_RXFF/n70 , \UART_RXFF/n69 ,
         \UART_RXFF/n68 , \UART_RXFF/n67 , \UART_RXFF/n66 , \UART_RXFF/n65 ,
         \UART_RXFF/n64 , \UART_RXFF/n63 , \UART_RXFF/n62 , \UART_RXFF/n61 ,
         \UART_RXFF/n60 , \UART_RXFF/n59 , \UART_RXFF/n58 , \UART_RXFF/n57 ,
         \UART_RXFF/n56 , \UART_RXFF/n55 , \UART_RXFF/n54 , \UART_RXFF/n53 ,
         \UART_RXFF/n52 , \UART_RXFF/n51 , \UART_RXFF/n50 , \UART_RXFF/n49 ,
         \UART_RXFF/n48 , \UART_RXFF/n47 , \UART_RXFF/n46 , \UART_RXFF/n44 ,
         \UART_RXFF/n43 , \UART_RXFF/n42 , \UART_RXFF/n40 , \UART_RXFF/n39 ,
         \UART_RXFF/n38 , \UART_RXFF/n37 , \UART_RXFF/n36 , \UART_RXFF/n35 ,
         \UART_RXFF/n34 , \UART_RXFF/n33 , \UART_RXFF/n32 , \UART_RXFF/n31 ,
         \UART_RXFF/n30 , \UART_RXFF/n29 , \UART_RXFF/n28 , \UART_RXFF/n27 ,
         \UART_RXFF/n26 , \UART_RXFF/n25 , \UART_RXFF/n24 , \UART_RXFF/n23 ,
         \UART_RXFF/n22 , \UART_RXFF/n21 , \UART_RXFF/n20 , \UART_RXFF/n19 ,
         \UART_RXFF/n18 , \UART_RXFF/n17 , \UART_RXFF/n16 , \UART_RXFF/n15 ,
         \UART_RXFF/n14 , \UART_RXFF/n13 , \UART_RXFF/n12 , \UART_RXFF/n11 ,
         \UART_RXFF/n10 , \UART_RXFF/n9 , \UART_RXFF/n8 , \UART_RXFF/n7 ,
         \UART_RXFF/n6 , \UART_RXFF/n5 , \UART_RXFF/n4 , \UART_RXFF/n3 ,
         \UART_RXFF/n2 , \UART_RXFF/n1 , \UART_RXFF/n2408 , \UART_RXFF/n2407 ,
         \UART_RXFF/n2406 , \UART_RXFF/n2405 , \UART_RXFF/n2404 ,
         \UART_RXFF/n2403 , \UART_RXFF/n2402 , \UART_RXFF/n2401 ,
         \UART_RXFF/n2400 , \UART_RXFF/n2399 , \UART_RXFF/n2398 ,
         \UART_RXFF/n2397 , \UART_RXFF/n2396 , \UART_RXFF/n2395 ,
         \UART_RXFF/n2394 , \UART_RXFF/n2393 , \UART_RXFF/n2392 ,
         \UART_RXFF/n2391 , \UART_RXFF/n2390 , \UART_RXFF/n2389 ,
         \UART_RXFF/n2388 , \UART_RXFF/n2387 , \UART_RXFF/n2386 ,
         \UART_RXFF/n2385 , \UART_RXFF/n2384 , \UART_RXFF/n2383 ,
         \UART_RXFF/n2382 , \UART_RXFF/n2381 , \UART_RXFF/n2380 ,
         \UART_RXFF/n2379 , \UART_RXFF/n2378 , \UART_RXFF/n2377 ,
         \UART_RXFF/n2376 , \UART_RXFF/n2375 , \UART_RXFF/n2374 ,
         \UART_RXFF/n2373 , \UART_RXFF/n2372 , \UART_RXFF/n2371 ,
         \UART_RXFF/n2370 , \UART_RXFF/n2369 , \UART_RXFF/n2368 ,
         \UART_RXFF/n2367 , \UART_RXFF/n2366 , \UART_RXFF/n2365 ,
         \UART_RXFF/n2364 , \UART_RXFF/n2363 , \UART_RXFF/n2362 ,
         \UART_RXFF/n2361 , \UART_RXFF/n2360 , \UART_RXFF/n2359 ,
         \UART_RXFF/n2358 , \UART_RXFF/n2357 , \UART_RXFF/n2356 ,
         \UART_RXFF/n2355 , \UART_RXFF/n2354 , \UART_RXFF/n2353 ,
         \UART_RXFF/n2352 , \UART_RXFF/n2351 , \UART_RXFF/n2350 ,
         \UART_RXFF/n2349 , \UART_RXFF/n2348 , \UART_RXFF/n2347 ,
         \UART_RXFF/n2346 , \UART_RXFF/n2345 , \UART_RXFF/n2344 ,
         \UART_RXFF/n2343 , \UART_RXFF/n2342 , \UART_RXFF/n2341 ,
         \UART_RXFF/n2340 , \UART_RXFF/n2339 , \UART_RXFF/n2338 ,
         \UART_RXFF/n2337 , \UART_RXFF/n2336 , \UART_RXFF/n2335 ,
         \UART_RXFF/n2334 , \UART_RXFF/n2333 , \UART_RXFF/n2332 ,
         \UART_RXFF/n2331 , \UART_RXFF/n2330 , \UART_RXFF/n2329 ,
         \UART_RXFF/n2328 , \UART_RXFF/n2327 , \UART_RXFF/n2326 ,
         \UART_RXFF/n2325 , \UART_RXFF/n2324 , \UART_RXFF/n2323 ,
         \UART_RXFF/n2322 , \UART_RXFF/n2321 , \UART_RXFF/n2320 ,
         \UART_RXFF/n2319 , \UART_RXFF/n2318 , \UART_RXFF/n2317 ,
         \UART_RXFF/n2316 , \UART_RXFF/n2315 , \UART_RXFF/n2314 ,
         \UART_RXFF/n2313 , \UART_RXFF/n2312 , \UART_RXFF/n2311 ,
         \UART_RXFF/n2310 , \UART_RXFF/n2309 , \UART_RXFF/n2308 ,
         \UART_RXFF/n2307 , \UART_RXFF/n2306 , \UART_RXFF/n2305 ,
         \UART_RXFF/n2304 , \UART_RXFF/n2303 , \UART_RXFF/n2302 ,
         \UART_RXFF/n2301 , \UART_RXFF/n2300 , \UART_RXFF/n2299 ,
         \UART_RXFF/n2298 , \UART_RXFF/n2297 , \UART_RXFF/n2296 ,
         \UART_RXFF/n2295 , \UART_RXFF/n2294 , \UART_RXFF/n2293 ,
         \UART_RXFF/n2292 , \UART_RXFF/n2291 , \UART_RXFF/n2290 ,
         \UART_RXFF/n2289 , \UART_RXFF/n2288 , \UART_RXFF/n2287 ,
         \UART_RXFF/n2286 , \UART_RXFF/n2285 , \UART_RXFF/n2284 ,
         \UART_RXFF/n2283 , \UART_RXFF/n2282 , \UART_RXFF/n2281 ,
         \UART_RXFF/n2280 , \UART_RXFF/n2279 , \UART_RXFF/n2278 ,
         \UART_RXFF/n2277 , \UART_RXFF/n2276 , \UART_RXFF/n2275 ,
         \UART_RXFF/n2274 , \UART_RXFF/n2273 , \UART_RXFF/n2272 ,
         \UART_RXFF/n2271 , \UART_RXFF/n2270 , \UART_RXFF/n2269 ,
         \UART_RXFF/n2268 , \UART_RXFF/n2267 , \UART_RXFF/n2266 ,
         \UART_RXFF/n2265 , \UART_RXFF/n2264 , \UART_RXFF/n2263 ,
         \UART_RXFF/n2262 , \UART_RXFF/n2261 , \UART_RXFF/n2260 ,
         \UART_RXFF/n2259 , \UART_RXFF/n2258 , \UART_RXFF/n2257 ,
         \UART_RXFF/n2256 , \UART_RXFF/n2255 , \UART_RXFF/n2254 ,
         \UART_RXFF/n2253 , \UART_RXFF/n2252 , \UART_RXFF/n2251 ,
         \UART_RXFF/n2250 , \UART_RXFF/n2249 , \UART_RXFF/n2248 ,
         \UART_RXFF/n2247 , \UART_RXFF/n2246 , \UART_RXFF/n2245 ,
         \UART_RXFF/n2244 , \UART_RXFF/n2243 , \UART_RXFF/n2242 ,
         \UART_RXFF/n2241 , \UART_RXFF/n2240 , \UART_RXFF/n2239 ,
         \UART_RXFF/n2238 , \UART_RXFF/n2237 , \UART_RXFF/n2236 ,
         \UART_RXFF/n2235 , \UART_RXFF/n2234 , \UART_RXFF/n2233 ,
         \UART_RXFF/n2232 , \UART_RXFF/n2231 , \UART_RXFF/n2230 ,
         \UART_RXFF/n2229 , \UART_RXFF/n2228 , \UART_RXFF/n2227 ,
         \UART_RXFF/n2226 , \UART_RXFF/n2225 , \UART_RXFF/n2224 ,
         \UART_RXFF/n2223 , \UART_RXFF/n2222 , \UART_RXFF/n2221 ,
         \UART_RXFF/n2220 , \UART_RXFF/n2219 , \UART_RXFF/n2218 ,
         \UART_RXFF/n2217 , \UART_RXFF/n2216 , \UART_RXFF/n2215 ,
         \UART_RXFF/n2214 , \UART_RXFF/n2213 , \UART_RXFF/n2212 ,
         \UART_RXFF/n2211 , \UART_RXFF/n2210 , \UART_RXFF/n2209 ,
         \UART_RXFF/n2208 , \UART_RXFF/n2207 , \UART_RXFF/n2206 ,
         \UART_RXFF/n2205 , \UART_RXFF/n2204 , \UART_RXFF/n2203 ,
         \UART_RXFF/n2202 , \UART_RXFF/n2201 , \UART_RXFF/n2200 ,
         \UART_RXFF/n2199 , \UART_RXFF/n2198 , \UART_RXFF/n2197 ,
         \UART_RXFF/n2196 , \UART_RXFF/n2195 , \UART_RXFF/n2194 ,
         \UART_RXFF/n2193 , \UART_RXFF/n2192 , \UART_RXFF/n2191 ,
         \UART_RXFF/n2190 , \UART_RXFF/n2189 , \UART_RXFF/n2188 ,
         \UART_RXFF/n2187 , \UART_RXFF/n2186 , \UART_RXFF/n2185 ,
         \UART_RXFF/n2184 , \UART_RXFF/n2183 , \UART_RXFF/n2182 ,
         \UART_RXFF/n2181 , \UART_RXFF/n2180 , \UART_RXFF/n2179 ,
         \UART_RXFF/n2178 , \UART_RXFF/n2177 , \UART_RXFF/n2176 ,
         \UART_RXFF/n2175 , \UART_RXFF/n2174 , \UART_RXFF/n2173 ,
         \UART_RXFF/n2172 , \UART_RXFF/n2171 , \UART_RXFF/n2170 ,
         \UART_RXFF/n2169 , \UART_RXFF/n2168 , \UART_RXFF/n2167 ,
         \UART_RXFF/n2166 , \UART_RXFF/n2165 , \UART_RXFF/n2164 ,
         \UART_RXFF/n2163 , \UART_RXFF/n2162 , \UART_RXFF/n2161 ,
         \UART_RXFF/n2160 , \UART_RXFF/n2159 , \UART_RXFF/n2158 ,
         \UART_RXFF/n2157 , \UART_RXFF/n2156 , \UART_RXFF/n2155 ,
         \UART_RXFF/n2154 , \UART_RXFF/n2153 , \UART_RXFF/n2152 ,
         \UART_RXFF/n2151 , \UART_RXFF/n2150 , \UART_RXFF/n2149 ,
         \UART_RXFF/n2148 , \UART_RXFF/n2147 , \UART_RXFF/n2146 ,
         \UART_RXFF/n2145 , \UART_RXFF/n2144 , \UART_RXFF/n2143 ,
         \UART_RXFF/n2142 , \UART_RXFF/n2141 , \UART_RXFF/n2140 ,
         \UART_RXFF/n2139 , \UART_RXFF/n2138 , \UART_RXFF/n2137 ,
         \UART_RXFF/n2136 , \UART_RXFF/n2135 , \UART_RXFF/n2134 ,
         \UART_RXFF/n2133 , \UART_RXFF/n2132 , \UART_RXFF/n2131 ,
         \UART_RXFF/n2130 , \UART_RXFF/n2129 , \UART_RXFF/n2128 ,
         \UART_RXFF/n2127 , \UART_RXFF/n2126 , \UART_RXFF/n2125 ,
         \UART_RXFF/n2124 , \UART_RXFF/n2123 , \UART_RXFF/n2122 ,
         \UART_RXFF/n2121 , \UART_RXFF/n2120 , \UART_RXFF/n2119 ,
         \UART_RXFF/n2118 , \UART_RXFF/n2117 , \UART_RXFF/n2116 ,
         \UART_RXFF/n2115 , \UART_RXFF/n2114 , \UART_RXFF/n2113 ,
         \UART_RXFF/n2112 , \UART_RXFF/n2111 , \UART_RXFF/n2110 ,
         \UART_RXFF/n2109 , \UART_RXFF/n2108 , \UART_RXFF/n2107 ,
         \UART_RXFF/n2106 , \UART_RXFF/n2105 , \UART_RXFF/n2104 ,
         \UART_RXFF/n2103 , \UART_RXFF/n2102 , \UART_RXFF/n2101 ,
         \UART_RXFF/n2100 , \UART_RXFF/n2099 , \UART_RXFF/n2098 ,
         \UART_RXFF/n2097 , \UART_RXFF/n2096 , \UART_RXFF/n2095 ,
         \UART_RXFF/n2094 , \UART_RXFF/n2093 , \UART_RXFF/n2092 ,
         \UART_RXFF/n2091 , \UART_RXFF/n2090 , \UART_RXFF/n2089 ,
         \UART_RXFF/n2088 , \UART_RXFF/n2087 , \UART_RXFF/n2086 ,
         \UART_RXFF/n2085 , \UART_RXFF/n2084 , \UART_RXFF/n2083 ,
         \UART_RXFF/n2082 , \UART_RXFF/n2081 , \UART_RXFF/n2080 ,
         \UART_RXFF/n2079 , \UART_RXFF/n2078 , \UART_RXFF/n2077 ,
         \UART_RXFF/n2076 , \UART_RXFF/n2075 , \UART_RXFF/n2074 ,
         \UART_RXFF/n2073 , \UART_RXFF/n2072 , \UART_RXFF/n2071 ,
         \UART_RXFF/n2070 , \UART_RXFF/n2069 , \UART_RXFF/n2068 ,
         \UART_RXFF/n2067 , \UART_RXFF/n2066 , \UART_RXFF/n2065 ,
         \UART_RXFF/n2064 , \UART_RXFF/n2063 , \UART_RXFF/n2062 ,
         \UART_RXFF/n2061 , \UART_RXFF/n2060 , \UART_RXFF/n2059 ,
         \UART_RXFF/n2058 , \UART_RXFF/n2057 , \UART_RXFF/n2056 ,
         \UART_RXFF/n2055 , \UART_RXFF/n2054 , \UART_RXFF/n2053 ,
         \UART_RXFF/n2052 , \UART_RXFF/n2051 , \UART_RXFF/n2050 ,
         \UART_RXFF/n2049 , \UART_RXFF/n2048 , \UART_RXFF/n2047 ,
         \UART_RXFF/n2046 , \UART_RXFF/n2045 , \UART_RXFF/n2044 ,
         \UART_RXFF/n2043 , \UART_RXFF/n2042 , \UART_RXFF/n2041 ,
         \UART_RXFF/n2040 , \UART_RXFF/n2039 , \UART_RXFF/n2038 ,
         \UART_RXFF/n2037 , \UART_RXFF/n2036 , \UART_RXFF/n2035 ,
         \UART_RXFF/n2034 , \UART_RXFF/n2033 , \UART_RXFF/n2032 ,
         \UART_RXFF/n2031 , \UART_RXFF/n2030 , \UART_RXFF/n2029 ,
         \UART_RXFF/n2028 , \UART_RXFF/n2027 , \UART_RXFF/n2026 ,
         \UART_RXFF/n2025 , \UART_RXFF/n2024 , \UART_RXFF/n2023 ,
         \UART_RXFF/n2022 , \UART_RXFF/n2021 , \UART_RXFF/n2020 ,
         \UART_RXFF/n2019 , \UART_RXFF/n2018 , \UART_RXFF/n2017 ,
         \UART_RXFF/n2016 , \UART_RXFF/n2015 , \UART_RXFF/n2014 ,
         \UART_RXFF/n2013 , \UART_RXFF/n2012 , \UART_RXFF/n2011 ,
         \UART_RXFF/n2010 , \UART_RXFF/n2009 , \UART_RXFF/n2008 ,
         \UART_RXFF/n2007 , \UART_RXFF/n2006 , \UART_RXFF/n2005 ,
         \UART_RXFF/n2004 , \UART_RXFF/n2003 , \UART_RXFF/n2002 ,
         \UART_RXFF/n2001 , \UART_RXFF/n2000 , \UART_RXFF/n1999 ,
         \UART_RXFF/n1998 , \UART_RXFF/n1997 , \UART_RXFF/n1996 ,
         \UART_RXFF/n1995 , \UART_RXFF/n1994 , \UART_RXFF/n1993 ,
         \UART_RXFF/n1992 , \UART_RXFF/n1991 , \UART_RXFF/n1990 ,
         \UART_RXFF/n1989 , \UART_RXFF/n1988 , \UART_RXFF/n1987 ,
         \UART_RXFF/n1986 , \UART_RXFF/n1985 , \UART_RXFF/n1984 ,
         \UART_RXFF/n1983 , \UART_RXFF/n1982 , \UART_RXFF/n1981 ,
         \UART_RXFF/n1980 , \UART_RXFF/n1979 , \UART_RXFF/n1978 ,
         \UART_RXFF/n1977 , \UART_RXFF/n1976 , \UART_RXFF/n1975 ,
         \UART_RXFF/n1974 , \UART_RXFF/n1973 , \UART_RXFF/n1972 ,
         \UART_RXFF/n1971 , \UART_RXFF/n1970 , \UART_RXFF/n1969 ,
         \UART_RXFF/n1968 , \UART_RXFF/n1967 , \UART_RXFF/n1966 ,
         \UART_RXFF/n1965 , \UART_RXFF/n1964 , \UART_RXFF/n1963 ,
         \UART_RXFF/n1962 , \UART_RXFF/n1961 , \UART_RXFF/n1960 ,
         \UART_RXFF/n1959 , \UART_RXFF/n1958 , \UART_RXFF/n1957 ,
         \UART_RXFF/n1956 , \UART_RXFF/n1955 , \UART_RXFF/n1954 ,
         \UART_RXFF/n1953 , \UART_RXFF/n1952 , \UART_RXFF/n1951 ,
         \UART_RXFF/n1950 , \UART_RXFF/n1949 , \UART_RXFF/n1948 ,
         \UART_RXFF/n1947 , \UART_RXFF/n1946 , \UART_RXFF/n1945 ,
         \UART_RXFF/n1944 , \UART_RXFF/n1943 , \UART_RXFF/n1942 ,
         \UART_RXFF/n1941 , \UART_RXFF/n1940 , \UART_RXFF/n1939 ,
         \UART_RXFF/n1938 , \UART_RXFF/n1937 , \UART_RXFF/n1936 ,
         \UART_RXFF/n1935 , \UART_RXFF/n1934 , \UART_RXFF/n1933 ,
         \UART_RXFF/n1932 , \UART_RXFF/n1931 , \UART_RXFF/n1930 ,
         \UART_RXFF/n1929 , \UART_RXFF/n1928 , \UART_RXFF/n1927 ,
         \UART_RXFF/n1926 , \UART_RXFF/n1925 , \UART_RXFF/n1924 ,
         \UART_RXFF/n1923 , \UART_RXFF/n1922 , \UART_RXFF/n1921 ,
         \UART_RXFF/n1920 , \UART_RXFF/n1919 , \UART_RXFF/n1918 ,
         \UART_RXFF/n1917 , \UART_RXFF/n1916 , \UART_RXFF/n1915 ,
         \UART_RXFF/n1914 , \UART_RXFF/n1913 , \UART_RXFF/n1912 ,
         \UART_RXFF/n1911 , \UART_RXFF/n1910 , \UART_RXFF/n1909 ,
         \UART_RXFF/n1908 , \UART_RXFF/n1907 , \UART_RXFF/n1906 ,
         \UART_RXFF/n1905 , \UART_RXFF/n1904 , \UART_RXFF/n1903 ,
         \UART_RXFF/n1902 , \UART_RXFF/n1901 , \UART_RXFF/n1900 ,
         \UART_RXFF/n1899 , \UART_RXFF/n1898 , \UART_RXFF/n1897 ,
         \UART_RXFF/n1896 , \UART_RXFF/n1895 , \UART_RXFF/n1894 ,
         \UART_RXFF/n1893 , \UART_RXFF/n1892 , \UART_RXFF/n1891 ,
         \UART_RXFF/n1890 , \UART_RXFF/n1889 , \UART_RXFF/n1888 ,
         \UART_RXFF/n1887 , \UART_RXFF/n1886 , \UART_RXFF/n1885 ,
         \UART_RXFF/n1884 , \UART_RXFF/n1883 , \UART_RXFF/n1882 ,
         \UART_RXFF/n1881 , \UART_RXFF/n1880 , \UART_RXFF/n1879 ,
         \UART_RXFF/n1878 , \UART_RXFF/n1877 , \UART_RXFF/n1876 ,
         \UART_RXFF/n1875 , \UART_RXFF/n1874 , \UART_RXFF/n1873 ,
         \UART_RXFF/n1872 , \UART_RXFF/n1871 , \UART_RXFF/n1870 ,
         \UART_RXFF/n1869 , \UART_RXFF/n1868 , \UART_RXFF/n1867 ,
         \UART_RXFF/n1866 , \UART_RXFF/n1865 , \UART_RXFF/n1864 ,
         \UART_RXFF/n1863 , \UART_RXFF/n1862 , \UART_RXFF/n1861 ,
         \UART_RXFF/n1860 , \UART_RXFF/n1859 , \UART_RXFF/n1858 ,
         \UART_RXFF/n1857 , \UART_RXFF/n1856 , \UART_RXFF/n1855 ,
         \UART_RXFF/n1854 , \UART_RXFF/n1853 , \UART_RXFF/n1852 ,
         \UART_RXFF/n1851 , \UART_RXFF/n1850 , \UART_RXFF/n1849 ,
         \UART_RXFF/n1848 , \UART_RXFF/n1847 , \UART_RXFF/n1846 ,
         \UART_RXFF/n1845 , \UART_RXFF/n1844 , \UART_RXFF/n1843 ,
         \UART_RXFF/n1842 , \UART_RXFF/n1841 , \UART_RXFF/n1840 ,
         \UART_RXFF/n1839 , \UART_RXFF/n1838 , \UART_RXFF/n1837 ,
         \UART_RXFF/n1836 , \UART_RXFF/n1835 , \UART_RXFF/n1834 ,
         \UART_RXFF/n1833 , \UART_RXFF/n1832 , \UART_RXFF/n1831 ,
         \UART_RXFF/n1830 , \UART_RXFF/n1829 , \UART_RXFF/n1828 ,
         \UART_RXFF/n1827 , \UART_RXFF/n1826 , \UART_RXFF/n1825 ,
         \UART_RXFF/n1824 , \UART_RXFF/n1823 , \UART_RXFF/n1822 ,
         \UART_RXFF/n1821 , \UART_RXFF/n1820 , \UART_RXFF/n1819 ,
         \UART_RXFF/n1818 , \UART_RXFF/n1817 , \UART_RXFF/n1816 ,
         \UART_RXFF/n1815 , \UART_RXFF/n1814 , \UART_RXFF/n1813 ,
         \UART_RXFF/n1812 , \UART_RXFF/n1811 , \UART_RXFF/n1810 ,
         \UART_RXFF/n1809 , \UART_RXFF/n1808 , \UART_RXFF/n1807 ,
         \UART_RXFF/n1806 , \UART_RXFF/n1805 , \UART_RXFF/n1804 ,
         \UART_RXFF/n1803 , \UART_RXFF/n1802 , \UART_RXFF/n1801 ,
         \UART_RXFF/n1800 , \UART_RXFF/n1799 , \UART_RXFF/n1798 ,
         \UART_RXFF/n1797 , \UART_RXFF/n1796 , \UART_RXFF/n1795 ,
         \UART_RXFF/n1794 , \UART_RXFF/n1793 , \UART_RXFF/n1792 ,
         \UART_RXFF/n1791 , \UART_RXFF/n1790 , \UART_RXFF/n1789 ,
         \UART_RXFF/n1788 , \UART_RXFF/n1787 , \UART_RXFF/n1786 ,
         \UART_RXFF/n1785 , \UART_RXFF/n1784 , \UART_RXFF/n1783 ,
         \UART_RXFF/n1782 , \UART_RXFF/n1781 , \UART_RXFF/n1780 ,
         \UART_RXFF/n1779 , \UART_RXFF/n1778 , \UART_RXFF/n1777 ,
         \UART_RXFF/n1776 , \UART_RXFF/n1775 , \UART_RXFF/n1774 ,
         \UART_RXFF/n1773 , \UART_RXFF/n1772 , \UART_RXFF/n1771 ,
         \UART_RXFF/n1770 , \UART_RXFF/n1769 , \UART_RXFF/n1768 ,
         \UART_RXFF/n1767 , \UART_RXFF/n1766 , \UART_RXFF/n1765 ,
         \UART_RXFF/n1764 , \UART_RXFF/n1763 , \UART_RXFF/n1762 ,
         \UART_RXFF/n1761 , \UART_RXFF/n1760 , \UART_RXFF/n1759 ,
         \UART_RXFF/n1758 , \UART_RXFF/n1757 , \UART_RXFF/n1756 ,
         \UART_RXFF/n1755 , \UART_RXFF/n1754 , \UART_RXFF/n1753 ,
         \UART_RXFF/n1752 , \UART_RXFF/n1751 , \UART_RXFF/n1750 ,
         \UART_RXFF/n1749 , \UART_RXFF/n1748 , \UART_RXFF/n1747 ,
         \UART_RXFF/n1746 , \UART_RXFF/n1745 , \UART_RXFF/n1744 ,
         \UART_RXFF/n1743 , \UART_RXFF/n1742 , \UART_RXFF/n1741 ,
         \UART_RXFF/n1740 , \UART_RXFF/n1739 , \UART_RXFF/n1738 ,
         \UART_RXFF/n1737 , \UART_RXFF/n1736 , \UART_RXFF/n1735 ,
         \UART_RXFF/n1734 , \UART_RXFF/n1733 , \UART_RXFF/n1732 ,
         \UART_RXFF/n1731 , \UART_RXFF/n1730 , \UART_RXFF/n1729 ,
         \UART_RXFF/n1728 , \UART_RXFF/n1727 , \UART_RXFF/n1726 ,
         \UART_RXFF/n1725 , \UART_RXFF/n1724 , \UART_RXFF/n1723 ,
         \UART_RXFF/n1722 , \UART_RXFF/n1721 , \UART_RXFF/n1720 ,
         \UART_RXFF/n1719 , \UART_RXFF/n1718 , \UART_RXFF/n1717 ,
         \UART_RXFF/n1716 , \UART_RXFF/n1715 , \UART_RXFF/n1714 ,
         \UART_RXFF/n1713 , \UART_RXFF/n1712 , \UART_RXFF/n1711 ,
         \UART_RXFF/n1710 , \UART_RXFF/n1709 , \UART_RXFF/n1708 ,
         \UART_RXFF/n1707 , \UART_RXFF/n1706 , \UART_RXFF/n1705 ,
         \UART_RXFF/n1704 , \UART_RXFF/n1703 , \UART_RXFF/n1702 ,
         \UART_RXFF/n1701 , \UART_RXFF/n1700 , \UART_RXFF/n1699 ,
         \UART_RXFF/n1698 , \UART_RXFF/n1697 , \UART_RXFF/n1696 ,
         \UART_RXFF/n1695 , \UART_RXFF/n1694 , \UART_RXFF/n1693 ,
         \UART_RXFF/n1692 , \UART_RXFF/n1691 , \UART_RXFF/n1690 ,
         \UART_RXFF/n1689 , \UART_RXFF/n1688 , \UART_RXFF/n1687 ,
         \UART_RXFF/n1686 , \UART_RXFF/n1685 , \UART_RXFF/n979 ,
         \UART_RXFF/n977 , \UART_RXFF/n975 , \UART_RXFF/n973 ,
         \UART_RXFF/n971 , \UART_RXFF/n969 , \UART_RXFF/n967 ,
         \UART_RXFF/n965 , \UART_RXFF/n963 , \UART_RXFF/n961 ,
         \UART_RXFF/n959 , \UART_RXFF/N133 , \UART_RXFF/N132 ,
         \UART_RXFF/N131 , \UART_RXFF/N130 , \UART_RXFF/N129 ,
         \UART_RXFF/N128 , \UART_RXFF/N127 , \UART_RXFF/N126 ,
         \UART_RXFF/N125 , \UART_RXFF/N124 , \UART_RXFF/N123 ,
         \UART_RXFF/iFIFOMem[0][0] , \UART_RXFF/iFIFOMem[0][1] ,
         \UART_RXFF/iFIFOMem[0][2] , \UART_RXFF/iFIFOMem[0][3] ,
         \UART_RXFF/iFIFOMem[0][4] , \UART_RXFF/iFIFOMem[0][5] ,
         \UART_RXFF/iFIFOMem[0][6] , \UART_RXFF/iFIFOMem[0][7] ,
         \UART_RXFF/iFIFOMem[0][8] , \UART_RXFF/iFIFOMem[0][9] ,
         \UART_RXFF/iFIFOMem[0][10] , \UART_RXFF/iFIFOMem[1][0] ,
         \UART_RXFF/iFIFOMem[1][1] , \UART_RXFF/iFIFOMem[1][2] ,
         \UART_RXFF/iFIFOMem[1][3] , \UART_RXFF/iFIFOMem[1][4] ,
         \UART_RXFF/iFIFOMem[1][5] , \UART_RXFF/iFIFOMem[1][6] ,
         \UART_RXFF/iFIFOMem[1][7] , \UART_RXFF/iFIFOMem[1][8] ,
         \UART_RXFF/iFIFOMem[1][9] , \UART_RXFF/iFIFOMem[1][10] ,
         \UART_RXFF/iFIFOMem[2][0] , \UART_RXFF/iFIFOMem[2][1] ,
         \UART_RXFF/iFIFOMem[2][2] , \UART_RXFF/iFIFOMem[2][3] ,
         \UART_RXFF/iFIFOMem[2][4] , \UART_RXFF/iFIFOMem[2][5] ,
         \UART_RXFF/iFIFOMem[2][6] , \UART_RXFF/iFIFOMem[2][7] ,
         \UART_RXFF/iFIFOMem[2][8] , \UART_RXFF/iFIFOMem[2][9] ,
         \UART_RXFF/iFIFOMem[2][10] , \UART_RXFF/iFIFOMem[3][0] ,
         \UART_RXFF/iFIFOMem[3][1] , \UART_RXFF/iFIFOMem[3][2] ,
         \UART_RXFF/iFIFOMem[3][3] , \UART_RXFF/iFIFOMem[3][4] ,
         \UART_RXFF/iFIFOMem[3][5] , \UART_RXFF/iFIFOMem[3][6] ,
         \UART_RXFF/iFIFOMem[3][7] , \UART_RXFF/iFIFOMem[3][8] ,
         \UART_RXFF/iFIFOMem[3][9] , \UART_RXFF/iFIFOMem[3][10] ,
         \UART_RXFF/iFIFOMem[4][0] , \UART_RXFF/iFIFOMem[4][1] ,
         \UART_RXFF/iFIFOMem[4][2] , \UART_RXFF/iFIFOMem[4][3] ,
         \UART_RXFF/iFIFOMem[4][4] , \UART_RXFF/iFIFOMem[4][5] ,
         \UART_RXFF/iFIFOMem[4][6] , \UART_RXFF/iFIFOMem[4][7] ,
         \UART_RXFF/iFIFOMem[4][8] , \UART_RXFF/iFIFOMem[4][9] ,
         \UART_RXFF/iFIFOMem[4][10] , \UART_RXFF/iFIFOMem[5][0] ,
         \UART_RXFF/iFIFOMem[5][1] , \UART_RXFF/iFIFOMem[5][2] ,
         \UART_RXFF/iFIFOMem[5][3] , \UART_RXFF/iFIFOMem[5][4] ,
         \UART_RXFF/iFIFOMem[5][5] , \UART_RXFF/iFIFOMem[5][6] ,
         \UART_RXFF/iFIFOMem[5][7] , \UART_RXFF/iFIFOMem[5][8] ,
         \UART_RXFF/iFIFOMem[5][9] , \UART_RXFF/iFIFOMem[5][10] ,
         \UART_RXFF/iFIFOMem[6][0] , \UART_RXFF/iFIFOMem[6][1] ,
         \UART_RXFF/iFIFOMem[6][2] , \UART_RXFF/iFIFOMem[6][3] ,
         \UART_RXFF/iFIFOMem[6][4] , \UART_RXFF/iFIFOMem[6][5] ,
         \UART_RXFF/iFIFOMem[6][6] , \UART_RXFF/iFIFOMem[6][7] ,
         \UART_RXFF/iFIFOMem[6][8] , \UART_RXFF/iFIFOMem[6][9] ,
         \UART_RXFF/iFIFOMem[6][10] , \UART_RXFF/iFIFOMem[7][0] ,
         \UART_RXFF/iFIFOMem[7][1] , \UART_RXFF/iFIFOMem[7][2] ,
         \UART_RXFF/iFIFOMem[7][3] , \UART_RXFF/iFIFOMem[7][4] ,
         \UART_RXFF/iFIFOMem[7][5] , \UART_RXFF/iFIFOMem[7][6] ,
         \UART_RXFF/iFIFOMem[7][7] , \UART_RXFF/iFIFOMem[7][8] ,
         \UART_RXFF/iFIFOMem[7][9] , \UART_RXFF/iFIFOMem[7][10] ,
         \UART_RXFF/iFIFOMem[8][0] , \UART_RXFF/iFIFOMem[8][1] ,
         \UART_RXFF/iFIFOMem[8][2] , \UART_RXFF/iFIFOMem[8][3] ,
         \UART_RXFF/iFIFOMem[8][4] , \UART_RXFF/iFIFOMem[8][5] ,
         \UART_RXFF/iFIFOMem[8][6] , \UART_RXFF/iFIFOMem[8][7] ,
         \UART_RXFF/iFIFOMem[8][8] , \UART_RXFF/iFIFOMem[8][9] ,
         \UART_RXFF/iFIFOMem[8][10] , \UART_RXFF/iFIFOMem[9][0] ,
         \UART_RXFF/iFIFOMem[9][1] , \UART_RXFF/iFIFOMem[9][2] ,
         \UART_RXFF/iFIFOMem[9][3] , \UART_RXFF/iFIFOMem[9][4] ,
         \UART_RXFF/iFIFOMem[9][5] , \UART_RXFF/iFIFOMem[9][6] ,
         \UART_RXFF/iFIFOMem[9][7] , \UART_RXFF/iFIFOMem[9][8] ,
         \UART_RXFF/iFIFOMem[9][9] , \UART_RXFF/iFIFOMem[9][10] ,
         \UART_RXFF/iFIFOMem[10][0] , \UART_RXFF/iFIFOMem[10][1] ,
         \UART_RXFF/iFIFOMem[10][2] , \UART_RXFF/iFIFOMem[10][3] ,
         \UART_RXFF/iFIFOMem[10][4] , \UART_RXFF/iFIFOMem[10][5] ,
         \UART_RXFF/iFIFOMem[10][6] , \UART_RXFF/iFIFOMem[10][7] ,
         \UART_RXFF/iFIFOMem[10][8] , \UART_RXFF/iFIFOMem[10][9] ,
         \UART_RXFF/iFIFOMem[10][10] , \UART_RXFF/iFIFOMem[11][0] ,
         \UART_RXFF/iFIFOMem[11][1] , \UART_RXFF/iFIFOMem[11][2] ,
         \UART_RXFF/iFIFOMem[11][3] , \UART_RXFF/iFIFOMem[11][4] ,
         \UART_RXFF/iFIFOMem[11][5] , \UART_RXFF/iFIFOMem[11][6] ,
         \UART_RXFF/iFIFOMem[11][7] , \UART_RXFF/iFIFOMem[11][8] ,
         \UART_RXFF/iFIFOMem[11][9] , \UART_RXFF/iFIFOMem[11][10] ,
         \UART_RXFF/iFIFOMem[12][0] , \UART_RXFF/iFIFOMem[12][1] ,
         \UART_RXFF/iFIFOMem[12][2] , \UART_RXFF/iFIFOMem[12][3] ,
         \UART_RXFF/iFIFOMem[12][4] , \UART_RXFF/iFIFOMem[12][5] ,
         \UART_RXFF/iFIFOMem[12][6] , \UART_RXFF/iFIFOMem[12][7] ,
         \UART_RXFF/iFIFOMem[12][8] , \UART_RXFF/iFIFOMem[12][9] ,
         \UART_RXFF/iFIFOMem[12][10] , \UART_RXFF/iFIFOMem[13][0] ,
         \UART_RXFF/iFIFOMem[13][1] , \UART_RXFF/iFIFOMem[13][2] ,
         \UART_RXFF/iFIFOMem[13][3] , \UART_RXFF/iFIFOMem[13][4] ,
         \UART_RXFF/iFIFOMem[13][5] , \UART_RXFF/iFIFOMem[13][6] ,
         \UART_RXFF/iFIFOMem[13][7] , \UART_RXFF/iFIFOMem[13][8] ,
         \UART_RXFF/iFIFOMem[13][9] , \UART_RXFF/iFIFOMem[13][10] ,
         \UART_RXFF/iFIFOMem[14][0] , \UART_RXFF/iFIFOMem[14][1] ,
         \UART_RXFF/iFIFOMem[14][2] , \UART_RXFF/iFIFOMem[14][3] ,
         \UART_RXFF/iFIFOMem[14][4] , \UART_RXFF/iFIFOMem[14][5] ,
         \UART_RXFF/iFIFOMem[14][6] , \UART_RXFF/iFIFOMem[14][7] ,
         \UART_RXFF/iFIFOMem[14][8] , \UART_RXFF/iFIFOMem[14][9] ,
         \UART_RXFF/iFIFOMem[14][10] , \UART_RXFF/iFIFOMem[15][0] ,
         \UART_RXFF/iFIFOMem[15][1] , \UART_RXFF/iFIFOMem[15][2] ,
         \UART_RXFF/iFIFOMem[15][3] , \UART_RXFF/iFIFOMem[15][4] ,
         \UART_RXFF/iFIFOMem[15][5] , \UART_RXFF/iFIFOMem[15][6] ,
         \UART_RXFF/iFIFOMem[15][7] , \UART_RXFF/iFIFOMem[15][8] ,
         \UART_RXFF/iFIFOMem[15][9] , \UART_RXFF/iFIFOMem[15][10] ,
         \UART_RXFF/iFIFOMem[16][0] , \UART_RXFF/iFIFOMem[16][1] ,
         \UART_RXFF/iFIFOMem[16][2] , \UART_RXFF/iFIFOMem[16][3] ,
         \UART_RXFF/iFIFOMem[16][4] , \UART_RXFF/iFIFOMem[16][5] ,
         \UART_RXFF/iFIFOMem[16][6] , \UART_RXFF/iFIFOMem[16][7] ,
         \UART_RXFF/iFIFOMem[16][8] , \UART_RXFF/iFIFOMem[16][9] ,
         \UART_RXFF/iFIFOMem[16][10] , \UART_RXFF/iFIFOMem[17][0] ,
         \UART_RXFF/iFIFOMem[17][1] , \UART_RXFF/iFIFOMem[17][2] ,
         \UART_RXFF/iFIFOMem[17][3] , \UART_RXFF/iFIFOMem[17][4] ,
         \UART_RXFF/iFIFOMem[17][5] , \UART_RXFF/iFIFOMem[17][6] ,
         \UART_RXFF/iFIFOMem[17][7] , \UART_RXFF/iFIFOMem[17][8] ,
         \UART_RXFF/iFIFOMem[17][9] , \UART_RXFF/iFIFOMem[17][10] ,
         \UART_RXFF/iFIFOMem[18][0] , \UART_RXFF/iFIFOMem[18][1] ,
         \UART_RXFF/iFIFOMem[18][2] , \UART_RXFF/iFIFOMem[18][3] ,
         \UART_RXFF/iFIFOMem[18][4] , \UART_RXFF/iFIFOMem[18][5] ,
         \UART_RXFF/iFIFOMem[18][6] , \UART_RXFF/iFIFOMem[18][7] ,
         \UART_RXFF/iFIFOMem[18][8] , \UART_RXFF/iFIFOMem[18][9] ,
         \UART_RXFF/iFIFOMem[18][10] , \UART_RXFF/iFIFOMem[19][0] ,
         \UART_RXFF/iFIFOMem[19][1] , \UART_RXFF/iFIFOMem[19][2] ,
         \UART_RXFF/iFIFOMem[19][3] , \UART_RXFF/iFIFOMem[19][4] ,
         \UART_RXFF/iFIFOMem[19][5] , \UART_RXFF/iFIFOMem[19][6] ,
         \UART_RXFF/iFIFOMem[19][7] , \UART_RXFF/iFIFOMem[19][8] ,
         \UART_RXFF/iFIFOMem[19][9] , \UART_RXFF/iFIFOMem[19][10] ,
         \UART_RXFF/iFIFOMem[20][0] , \UART_RXFF/iFIFOMem[20][1] ,
         \UART_RXFF/iFIFOMem[20][2] , \UART_RXFF/iFIFOMem[20][3] ,
         \UART_RXFF/iFIFOMem[20][4] , \UART_RXFF/iFIFOMem[20][5] ,
         \UART_RXFF/iFIFOMem[20][6] , \UART_RXFF/iFIFOMem[20][7] ,
         \UART_RXFF/iFIFOMem[20][8] , \UART_RXFF/iFIFOMem[20][9] ,
         \UART_RXFF/iFIFOMem[20][10] , \UART_RXFF/iFIFOMem[21][0] ,
         \UART_RXFF/iFIFOMem[21][1] , \UART_RXFF/iFIFOMem[21][2] ,
         \UART_RXFF/iFIFOMem[21][3] , \UART_RXFF/iFIFOMem[21][4] ,
         \UART_RXFF/iFIFOMem[21][5] , \UART_RXFF/iFIFOMem[21][6] ,
         \UART_RXFF/iFIFOMem[21][7] , \UART_RXFF/iFIFOMem[21][8] ,
         \UART_RXFF/iFIFOMem[21][9] , \UART_RXFF/iFIFOMem[21][10] ,
         \UART_RXFF/iFIFOMem[22][0] , \UART_RXFF/iFIFOMem[22][1] ,
         \UART_RXFF/iFIFOMem[22][2] , \UART_RXFF/iFIFOMem[22][3] ,
         \UART_RXFF/iFIFOMem[22][4] , \UART_RXFF/iFIFOMem[22][5] ,
         \UART_RXFF/iFIFOMem[22][6] , \UART_RXFF/iFIFOMem[22][7] ,
         \UART_RXFF/iFIFOMem[22][8] , \UART_RXFF/iFIFOMem[22][9] ,
         \UART_RXFF/iFIFOMem[22][10] , \UART_RXFF/iFIFOMem[23][0] ,
         \UART_RXFF/iFIFOMem[23][1] , \UART_RXFF/iFIFOMem[23][2] ,
         \UART_RXFF/iFIFOMem[23][3] , \UART_RXFF/iFIFOMem[23][4] ,
         \UART_RXFF/iFIFOMem[23][5] , \UART_RXFF/iFIFOMem[23][6] ,
         \UART_RXFF/iFIFOMem[23][7] , \UART_RXFF/iFIFOMem[23][8] ,
         \UART_RXFF/iFIFOMem[23][9] , \UART_RXFF/iFIFOMem[23][10] ,
         \UART_RXFF/iFIFOMem[24][0] , \UART_RXFF/iFIFOMem[24][1] ,
         \UART_RXFF/iFIFOMem[24][2] , \UART_RXFF/iFIFOMem[24][3] ,
         \UART_RXFF/iFIFOMem[24][4] , \UART_RXFF/iFIFOMem[24][5] ,
         \UART_RXFF/iFIFOMem[24][6] , \UART_RXFF/iFIFOMem[24][7] ,
         \UART_RXFF/iFIFOMem[24][8] , \UART_RXFF/iFIFOMem[24][9] ,
         \UART_RXFF/iFIFOMem[24][10] , \UART_RXFF/iFIFOMem[25][0] ,
         \UART_RXFF/iFIFOMem[25][1] , \UART_RXFF/iFIFOMem[25][2] ,
         \UART_RXFF/iFIFOMem[25][3] , \UART_RXFF/iFIFOMem[25][4] ,
         \UART_RXFF/iFIFOMem[25][5] , \UART_RXFF/iFIFOMem[25][6] ,
         \UART_RXFF/iFIFOMem[25][7] , \UART_RXFF/iFIFOMem[25][8] ,
         \UART_RXFF/iFIFOMem[25][9] , \UART_RXFF/iFIFOMem[25][10] ,
         \UART_RXFF/iFIFOMem[26][0] , \UART_RXFF/iFIFOMem[26][1] ,
         \UART_RXFF/iFIFOMem[26][2] , \UART_RXFF/iFIFOMem[26][3] ,
         \UART_RXFF/iFIFOMem[26][4] , \UART_RXFF/iFIFOMem[26][5] ,
         \UART_RXFF/iFIFOMem[26][6] , \UART_RXFF/iFIFOMem[26][7] ,
         \UART_RXFF/iFIFOMem[26][8] , \UART_RXFF/iFIFOMem[26][9] ,
         \UART_RXFF/iFIFOMem[26][10] , \UART_RXFF/iFIFOMem[27][0] ,
         \UART_RXFF/iFIFOMem[27][1] , \UART_RXFF/iFIFOMem[27][2] ,
         \UART_RXFF/iFIFOMem[27][3] , \UART_RXFF/iFIFOMem[27][4] ,
         \UART_RXFF/iFIFOMem[27][5] , \UART_RXFF/iFIFOMem[27][6] ,
         \UART_RXFF/iFIFOMem[27][7] , \UART_RXFF/iFIFOMem[27][8] ,
         \UART_RXFF/iFIFOMem[27][9] , \UART_RXFF/iFIFOMem[27][10] ,
         \UART_RXFF/iFIFOMem[28][0] , \UART_RXFF/iFIFOMem[28][1] ,
         \UART_RXFF/iFIFOMem[28][2] , \UART_RXFF/iFIFOMem[28][3] ,
         \UART_RXFF/iFIFOMem[28][4] , \UART_RXFF/iFIFOMem[28][5] ,
         \UART_RXFF/iFIFOMem[28][6] , \UART_RXFF/iFIFOMem[28][7] ,
         \UART_RXFF/iFIFOMem[28][8] , \UART_RXFF/iFIFOMem[28][9] ,
         \UART_RXFF/iFIFOMem[28][10] , \UART_RXFF/iFIFOMem[29][0] ,
         \UART_RXFF/iFIFOMem[29][1] , \UART_RXFF/iFIFOMem[29][2] ,
         \UART_RXFF/iFIFOMem[29][3] , \UART_RXFF/iFIFOMem[29][4] ,
         \UART_RXFF/iFIFOMem[29][5] , \UART_RXFF/iFIFOMem[29][6] ,
         \UART_RXFF/iFIFOMem[29][7] , \UART_RXFF/iFIFOMem[29][8] ,
         \UART_RXFF/iFIFOMem[29][9] , \UART_RXFF/iFIFOMem[29][10] ,
         \UART_RXFF/iFIFOMem[30][0] , \UART_RXFF/iFIFOMem[30][1] ,
         \UART_RXFF/iFIFOMem[30][2] , \UART_RXFF/iFIFOMem[30][3] ,
         \UART_RXFF/iFIFOMem[30][4] , \UART_RXFF/iFIFOMem[30][5] ,
         \UART_RXFF/iFIFOMem[30][6] , \UART_RXFF/iFIFOMem[30][7] ,
         \UART_RXFF/iFIFOMem[30][8] , \UART_RXFF/iFIFOMem[30][9] ,
         \UART_RXFF/iFIFOMem[30][10] , \UART_RXFF/iFIFOMem[31][0] ,
         \UART_RXFF/iFIFOMem[31][1] , \UART_RXFF/iFIFOMem[31][2] ,
         \UART_RXFF/iFIFOMem[31][3] , \UART_RXFF/iFIFOMem[31][4] ,
         \UART_RXFF/iFIFOMem[31][5] , \UART_RXFF/iFIFOMem[31][6] ,
         \UART_RXFF/iFIFOMem[31][7] , \UART_RXFF/iFIFOMem[31][8] ,
         \UART_RXFF/iFIFOMem[31][9] , \UART_RXFF/iFIFOMem[31][10] ,
         \UART_RXFF/iFIFOMem[32][0] , \UART_RXFF/iFIFOMem[32][1] ,
         \UART_RXFF/iFIFOMem[32][2] , \UART_RXFF/iFIFOMem[32][3] ,
         \UART_RXFF/iFIFOMem[32][4] , \UART_RXFF/iFIFOMem[32][5] ,
         \UART_RXFF/iFIFOMem[32][6] , \UART_RXFF/iFIFOMem[32][7] ,
         \UART_RXFF/iFIFOMem[32][8] , \UART_RXFF/iFIFOMem[32][9] ,
         \UART_RXFF/iFIFOMem[32][10] , \UART_RXFF/iFIFOMem[33][0] ,
         \UART_RXFF/iFIFOMem[33][1] , \UART_RXFF/iFIFOMem[33][2] ,
         \UART_RXFF/iFIFOMem[33][3] , \UART_RXFF/iFIFOMem[33][4] ,
         \UART_RXFF/iFIFOMem[33][5] , \UART_RXFF/iFIFOMem[33][6] ,
         \UART_RXFF/iFIFOMem[33][7] , \UART_RXFF/iFIFOMem[33][8] ,
         \UART_RXFF/iFIFOMem[33][9] , \UART_RXFF/iFIFOMem[33][10] ,
         \UART_RXFF/iFIFOMem[34][0] , \UART_RXFF/iFIFOMem[34][1] ,
         \UART_RXFF/iFIFOMem[34][2] , \UART_RXFF/iFIFOMem[34][3] ,
         \UART_RXFF/iFIFOMem[34][4] , \UART_RXFF/iFIFOMem[34][5] ,
         \UART_RXFF/iFIFOMem[34][6] , \UART_RXFF/iFIFOMem[34][7] ,
         \UART_RXFF/iFIFOMem[34][8] , \UART_RXFF/iFIFOMem[34][9] ,
         \UART_RXFF/iFIFOMem[34][10] , \UART_RXFF/iFIFOMem[35][0] ,
         \UART_RXFF/iFIFOMem[35][1] , \UART_RXFF/iFIFOMem[35][2] ,
         \UART_RXFF/iFIFOMem[35][3] , \UART_RXFF/iFIFOMem[35][4] ,
         \UART_RXFF/iFIFOMem[35][5] , \UART_RXFF/iFIFOMem[35][6] ,
         \UART_RXFF/iFIFOMem[35][7] , \UART_RXFF/iFIFOMem[35][8] ,
         \UART_RXFF/iFIFOMem[35][9] , \UART_RXFF/iFIFOMem[35][10] ,
         \UART_RXFF/iFIFOMem[36][0] , \UART_RXFF/iFIFOMem[36][1] ,
         \UART_RXFF/iFIFOMem[36][2] , \UART_RXFF/iFIFOMem[36][3] ,
         \UART_RXFF/iFIFOMem[36][4] , \UART_RXFF/iFIFOMem[36][5] ,
         \UART_RXFF/iFIFOMem[36][6] , \UART_RXFF/iFIFOMem[36][7] ,
         \UART_RXFF/iFIFOMem[36][8] , \UART_RXFF/iFIFOMem[36][9] ,
         \UART_RXFF/iFIFOMem[36][10] , \UART_RXFF/iFIFOMem[37][0] ,
         \UART_RXFF/iFIFOMem[37][1] , \UART_RXFF/iFIFOMem[37][2] ,
         \UART_RXFF/iFIFOMem[37][3] , \UART_RXFF/iFIFOMem[37][4] ,
         \UART_RXFF/iFIFOMem[37][5] , \UART_RXFF/iFIFOMem[37][6] ,
         \UART_RXFF/iFIFOMem[37][7] , \UART_RXFF/iFIFOMem[37][8] ,
         \UART_RXFF/iFIFOMem[37][9] , \UART_RXFF/iFIFOMem[37][10] ,
         \UART_RXFF/iFIFOMem[38][0] , \UART_RXFF/iFIFOMem[38][1] ,
         \UART_RXFF/iFIFOMem[38][2] , \UART_RXFF/iFIFOMem[38][3] ,
         \UART_RXFF/iFIFOMem[38][4] , \UART_RXFF/iFIFOMem[38][5] ,
         \UART_RXFF/iFIFOMem[38][6] , \UART_RXFF/iFIFOMem[38][7] ,
         \UART_RXFF/iFIFOMem[38][8] , \UART_RXFF/iFIFOMem[38][9] ,
         \UART_RXFF/iFIFOMem[38][10] , \UART_RXFF/iFIFOMem[39][0] ,
         \UART_RXFF/iFIFOMem[39][1] , \UART_RXFF/iFIFOMem[39][2] ,
         \UART_RXFF/iFIFOMem[39][3] , \UART_RXFF/iFIFOMem[39][4] ,
         \UART_RXFF/iFIFOMem[39][5] , \UART_RXFF/iFIFOMem[39][6] ,
         \UART_RXFF/iFIFOMem[39][7] , \UART_RXFF/iFIFOMem[39][8] ,
         \UART_RXFF/iFIFOMem[39][9] , \UART_RXFF/iFIFOMem[39][10] ,
         \UART_RXFF/iFIFOMem[40][0] , \UART_RXFF/iFIFOMem[40][1] ,
         \UART_RXFF/iFIFOMem[40][2] , \UART_RXFF/iFIFOMem[40][3] ,
         \UART_RXFF/iFIFOMem[40][4] , \UART_RXFF/iFIFOMem[40][5] ,
         \UART_RXFF/iFIFOMem[40][6] , \UART_RXFF/iFIFOMem[40][7] ,
         \UART_RXFF/iFIFOMem[40][8] , \UART_RXFF/iFIFOMem[40][9] ,
         \UART_RXFF/iFIFOMem[40][10] , \UART_RXFF/iFIFOMem[41][0] ,
         \UART_RXFF/iFIFOMem[41][1] , \UART_RXFF/iFIFOMem[41][2] ,
         \UART_RXFF/iFIFOMem[41][3] , \UART_RXFF/iFIFOMem[41][4] ,
         \UART_RXFF/iFIFOMem[41][5] , \UART_RXFF/iFIFOMem[41][6] ,
         \UART_RXFF/iFIFOMem[41][7] , \UART_RXFF/iFIFOMem[41][8] ,
         \UART_RXFF/iFIFOMem[41][9] , \UART_RXFF/iFIFOMem[41][10] ,
         \UART_RXFF/iFIFOMem[42][0] , \UART_RXFF/iFIFOMem[42][1] ,
         \UART_RXFF/iFIFOMem[42][2] , \UART_RXFF/iFIFOMem[42][3] ,
         \UART_RXFF/iFIFOMem[42][4] , \UART_RXFF/iFIFOMem[42][5] ,
         \UART_RXFF/iFIFOMem[42][6] , \UART_RXFF/iFIFOMem[42][7] ,
         \UART_RXFF/iFIFOMem[42][8] , \UART_RXFF/iFIFOMem[42][9] ,
         \UART_RXFF/iFIFOMem[42][10] , \UART_RXFF/iFIFOMem[43][0] ,
         \UART_RXFF/iFIFOMem[43][1] , \UART_RXFF/iFIFOMem[43][2] ,
         \UART_RXFF/iFIFOMem[43][3] , \UART_RXFF/iFIFOMem[43][4] ,
         \UART_RXFF/iFIFOMem[43][5] , \UART_RXFF/iFIFOMem[43][6] ,
         \UART_RXFF/iFIFOMem[43][7] , \UART_RXFF/iFIFOMem[43][8] ,
         \UART_RXFF/iFIFOMem[43][9] , \UART_RXFF/iFIFOMem[43][10] ,
         \UART_RXFF/iFIFOMem[44][0] , \UART_RXFF/iFIFOMem[44][1] ,
         \UART_RXFF/iFIFOMem[44][2] , \UART_RXFF/iFIFOMem[44][3] ,
         \UART_RXFF/iFIFOMem[44][4] , \UART_RXFF/iFIFOMem[44][5] ,
         \UART_RXFF/iFIFOMem[44][6] , \UART_RXFF/iFIFOMem[44][7] ,
         \UART_RXFF/iFIFOMem[44][8] , \UART_RXFF/iFIFOMem[44][9] ,
         \UART_RXFF/iFIFOMem[44][10] , \UART_RXFF/iFIFOMem[45][0] ,
         \UART_RXFF/iFIFOMem[45][1] , \UART_RXFF/iFIFOMem[45][2] ,
         \UART_RXFF/iFIFOMem[45][3] , \UART_RXFF/iFIFOMem[45][4] ,
         \UART_RXFF/iFIFOMem[45][5] , \UART_RXFF/iFIFOMem[45][6] ,
         \UART_RXFF/iFIFOMem[45][7] , \UART_RXFF/iFIFOMem[45][8] ,
         \UART_RXFF/iFIFOMem[45][9] , \UART_RXFF/iFIFOMem[45][10] ,
         \UART_RXFF/iFIFOMem[46][0] , \UART_RXFF/iFIFOMem[46][1] ,
         \UART_RXFF/iFIFOMem[46][2] , \UART_RXFF/iFIFOMem[46][3] ,
         \UART_RXFF/iFIFOMem[46][4] , \UART_RXFF/iFIFOMem[46][5] ,
         \UART_RXFF/iFIFOMem[46][6] , \UART_RXFF/iFIFOMem[46][7] ,
         \UART_RXFF/iFIFOMem[46][8] , \UART_RXFF/iFIFOMem[46][9] ,
         \UART_RXFF/iFIFOMem[46][10] , \UART_RXFF/iFIFOMem[47][0] ,
         \UART_RXFF/iFIFOMem[47][1] , \UART_RXFF/iFIFOMem[47][2] ,
         \UART_RXFF/iFIFOMem[47][3] , \UART_RXFF/iFIFOMem[47][4] ,
         \UART_RXFF/iFIFOMem[47][5] , \UART_RXFF/iFIFOMem[47][6] ,
         \UART_RXFF/iFIFOMem[47][7] , \UART_RXFF/iFIFOMem[47][8] ,
         \UART_RXFF/iFIFOMem[47][9] , \UART_RXFF/iFIFOMem[47][10] ,
         \UART_RXFF/iFIFOMem[48][0] , \UART_RXFF/iFIFOMem[48][1] ,
         \UART_RXFF/iFIFOMem[48][2] , \UART_RXFF/iFIFOMem[48][3] ,
         \UART_RXFF/iFIFOMem[48][4] , \UART_RXFF/iFIFOMem[48][5] ,
         \UART_RXFF/iFIFOMem[48][6] , \UART_RXFF/iFIFOMem[48][7] ,
         \UART_RXFF/iFIFOMem[48][8] , \UART_RXFF/iFIFOMem[48][9] ,
         \UART_RXFF/iFIFOMem[48][10] , \UART_RXFF/iFIFOMem[49][0] ,
         \UART_RXFF/iFIFOMem[49][1] , \UART_RXFF/iFIFOMem[49][2] ,
         \UART_RXFF/iFIFOMem[49][3] , \UART_RXFF/iFIFOMem[49][4] ,
         \UART_RXFF/iFIFOMem[49][5] , \UART_RXFF/iFIFOMem[49][6] ,
         \UART_RXFF/iFIFOMem[49][7] , \UART_RXFF/iFIFOMem[49][8] ,
         \UART_RXFF/iFIFOMem[49][9] , \UART_RXFF/iFIFOMem[49][10] ,
         \UART_RXFF/iFIFOMem[50][0] , \UART_RXFF/iFIFOMem[50][1] ,
         \UART_RXFF/iFIFOMem[50][2] , \UART_RXFF/iFIFOMem[50][3] ,
         \UART_RXFF/iFIFOMem[50][4] , \UART_RXFF/iFIFOMem[50][5] ,
         \UART_RXFF/iFIFOMem[50][6] , \UART_RXFF/iFIFOMem[50][7] ,
         \UART_RXFF/iFIFOMem[50][8] , \UART_RXFF/iFIFOMem[50][9] ,
         \UART_RXFF/iFIFOMem[50][10] , \UART_RXFF/iFIFOMem[51][0] ,
         \UART_RXFF/iFIFOMem[51][1] , \UART_RXFF/iFIFOMem[51][2] ,
         \UART_RXFF/iFIFOMem[51][3] , \UART_RXFF/iFIFOMem[51][4] ,
         \UART_RXFF/iFIFOMem[51][5] , \UART_RXFF/iFIFOMem[51][6] ,
         \UART_RXFF/iFIFOMem[51][7] , \UART_RXFF/iFIFOMem[51][8] ,
         \UART_RXFF/iFIFOMem[51][9] , \UART_RXFF/iFIFOMem[51][10] ,
         \UART_RXFF/iFIFOMem[52][0] , \UART_RXFF/iFIFOMem[52][1] ,
         \UART_RXFF/iFIFOMem[52][2] , \UART_RXFF/iFIFOMem[52][3] ,
         \UART_RXFF/iFIFOMem[52][4] , \UART_RXFF/iFIFOMem[52][5] ,
         \UART_RXFF/iFIFOMem[52][6] , \UART_RXFF/iFIFOMem[52][7] ,
         \UART_RXFF/iFIFOMem[52][8] , \UART_RXFF/iFIFOMem[52][9] ,
         \UART_RXFF/iFIFOMem[52][10] , \UART_RXFF/iFIFOMem[53][0] ,
         \UART_RXFF/iFIFOMem[53][1] , \UART_RXFF/iFIFOMem[53][2] ,
         \UART_RXFF/iFIFOMem[53][3] , \UART_RXFF/iFIFOMem[53][4] ,
         \UART_RXFF/iFIFOMem[53][5] , \UART_RXFF/iFIFOMem[53][6] ,
         \UART_RXFF/iFIFOMem[53][7] , \UART_RXFF/iFIFOMem[53][8] ,
         \UART_RXFF/iFIFOMem[53][9] , \UART_RXFF/iFIFOMem[53][10] ,
         \UART_RXFF/iFIFOMem[54][0] , \UART_RXFF/iFIFOMem[54][1] ,
         \UART_RXFF/iFIFOMem[54][2] , \UART_RXFF/iFIFOMem[54][3] ,
         \UART_RXFF/iFIFOMem[54][4] , \UART_RXFF/iFIFOMem[54][5] ,
         \UART_RXFF/iFIFOMem[54][6] , \UART_RXFF/iFIFOMem[54][7] ,
         \UART_RXFF/iFIFOMem[54][8] , \UART_RXFF/iFIFOMem[54][9] ,
         \UART_RXFF/iFIFOMem[54][10] , \UART_RXFF/iFIFOMem[55][0] ,
         \UART_RXFF/iFIFOMem[55][1] , \UART_RXFF/iFIFOMem[55][2] ,
         \UART_RXFF/iFIFOMem[55][3] , \UART_RXFF/iFIFOMem[55][4] ,
         \UART_RXFF/iFIFOMem[55][5] , \UART_RXFF/iFIFOMem[55][6] ,
         \UART_RXFF/iFIFOMem[55][7] , \UART_RXFF/iFIFOMem[55][8] ,
         \UART_RXFF/iFIFOMem[55][9] , \UART_RXFF/iFIFOMem[55][10] ,
         \UART_RXFF/iFIFOMem[56][0] , \UART_RXFF/iFIFOMem[56][1] ,
         \UART_RXFF/iFIFOMem[56][2] , \UART_RXFF/iFIFOMem[56][3] ,
         \UART_RXFF/iFIFOMem[56][4] , \UART_RXFF/iFIFOMem[56][5] ,
         \UART_RXFF/iFIFOMem[56][6] , \UART_RXFF/iFIFOMem[56][7] ,
         \UART_RXFF/iFIFOMem[56][8] , \UART_RXFF/iFIFOMem[56][9] ,
         \UART_RXFF/iFIFOMem[56][10] , \UART_RXFF/iFIFOMem[57][0] ,
         \UART_RXFF/iFIFOMem[57][1] , \UART_RXFF/iFIFOMem[57][2] ,
         \UART_RXFF/iFIFOMem[57][3] , \UART_RXFF/iFIFOMem[57][4] ,
         \UART_RXFF/iFIFOMem[57][5] , \UART_RXFF/iFIFOMem[57][6] ,
         \UART_RXFF/iFIFOMem[57][7] , \UART_RXFF/iFIFOMem[57][8] ,
         \UART_RXFF/iFIFOMem[57][9] , \UART_RXFF/iFIFOMem[57][10] ,
         \UART_RXFF/iFIFOMem[58][0] , \UART_RXFF/iFIFOMem[58][1] ,
         \UART_RXFF/iFIFOMem[58][2] , \UART_RXFF/iFIFOMem[58][3] ,
         \UART_RXFF/iFIFOMem[58][4] , \UART_RXFF/iFIFOMem[58][5] ,
         \UART_RXFF/iFIFOMem[58][6] , \UART_RXFF/iFIFOMem[58][7] ,
         \UART_RXFF/iFIFOMem[58][8] , \UART_RXFF/iFIFOMem[58][9] ,
         \UART_RXFF/iFIFOMem[58][10] , \UART_RXFF/iFIFOMem[59][0] ,
         \UART_RXFF/iFIFOMem[59][1] , \UART_RXFF/iFIFOMem[59][2] ,
         \UART_RXFF/iFIFOMem[59][3] , \UART_RXFF/iFIFOMem[59][4] ,
         \UART_RXFF/iFIFOMem[59][5] , \UART_RXFF/iFIFOMem[59][6] ,
         \UART_RXFF/iFIFOMem[59][7] , \UART_RXFF/iFIFOMem[59][8] ,
         \UART_RXFF/iFIFOMem[59][9] , \UART_RXFF/iFIFOMem[59][10] ,
         \UART_RXFF/iFIFOMem[60][0] , \UART_RXFF/iFIFOMem[60][1] ,
         \UART_RXFF/iFIFOMem[60][2] , \UART_RXFF/iFIFOMem[60][3] ,
         \UART_RXFF/iFIFOMem[60][4] , \UART_RXFF/iFIFOMem[60][5] ,
         \UART_RXFF/iFIFOMem[60][6] , \UART_RXFF/iFIFOMem[60][7] ,
         \UART_RXFF/iFIFOMem[60][8] , \UART_RXFF/iFIFOMem[60][9] ,
         \UART_RXFF/iFIFOMem[60][10] , \UART_RXFF/iFIFOMem[61][0] ,
         \UART_RXFF/iFIFOMem[61][1] , \UART_RXFF/iFIFOMem[61][2] ,
         \UART_RXFF/iFIFOMem[61][3] , \UART_RXFF/iFIFOMem[61][4] ,
         \UART_RXFF/iFIFOMem[61][5] , \UART_RXFF/iFIFOMem[61][6] ,
         \UART_RXFF/iFIFOMem[61][7] , \UART_RXFF/iFIFOMem[61][8] ,
         \UART_RXFF/iFIFOMem[61][9] , \UART_RXFF/iFIFOMem[61][10] ,
         \UART_RXFF/iFIFOMem[62][0] , \UART_RXFF/iFIFOMem[62][1] ,
         \UART_RXFF/iFIFOMem[62][2] , \UART_RXFF/iFIFOMem[62][3] ,
         \UART_RXFF/iFIFOMem[62][4] , \UART_RXFF/iFIFOMem[62][5] ,
         \UART_RXFF/iFIFOMem[62][6] , \UART_RXFF/iFIFOMem[62][7] ,
         \UART_RXFF/iFIFOMem[62][8] , \UART_RXFF/iFIFOMem[62][9] ,
         \UART_RXFF/iFIFOMem[62][10] , \UART_RXFF/iFIFOMem[63][0] ,
         \UART_RXFF/iFIFOMem[63][1] , \UART_RXFF/iFIFOMem[63][2] ,
         \UART_RXFF/iFIFOMem[63][3] , \UART_RXFF/iFIFOMem[63][4] ,
         \UART_RXFF/iFIFOMem[63][5] , \UART_RXFF/iFIFOMem[63][6] ,
         \UART_RXFF/iFIFOMem[63][7] , \UART_RXFF/iFIFOMem[63][8] ,
         \UART_RXFF/iFIFOMem[63][9] , \UART_RXFF/iFIFOMem[63][10] ,
         \UART_RXFF/N56 , \UART_RXFF/N38 , \UART_RXFF/N37 , \UART_RXFF/N36 ,
         \UART_RXFF/N35 , \UART_RXFF/N34 , \UART_RXFF/N33 , \UART_RXFF/N30 ,
         \UART_RXFF/N29 , \UART_RXFF/N28 , \UART_RXFF/N27 , \UART_RXFF/N26 ,
         \UART_RXFF/N25 , \UART_RXFF/iWRAddr[0] , \UART_RXFF/iWRAddr[1] ,
         \UART_RXFF/iWRAddr[2] , \UART_RXFF/iWRAddr[3] ,
         \UART_RXFF/iWRAddr[4] , \UART_RXFF/iWRAddr[5] ,
         \UART_RXFF/iWRAddr[6] , \UART_RXFF/iRDAddr[6] , \UART_RXFF/USAGE[0] ,
         \UART_RXFF/N17 , \UART_RXFF/N16 , \UART_RXFF/N15 , \UART_RXFF/N14 ,
         \UART_RXFF/N13 , \UART_RXFF/N12 , \UART_TX/n84 , \UART_TX/n83 ,
         \UART_TX/n82 , \UART_TX/n81 , \UART_TX/n80 , \UART_TX/n79 ,
         \UART_TX/n78 , \UART_TX/n77 , \UART_TX/n76 , \UART_TX/n75 ,
         \UART_TX/n74 , \UART_TX/n73 , \UART_TX/n72 , \UART_TX/n71 ,
         \UART_TX/n70 , \UART_TX/n69 , \UART_TX/n68 , \UART_TX/n67 ,
         \UART_TX/n66 , \UART_TX/n65 , \UART_TX/n64 , \UART_TX/n63 ,
         \UART_TX/n62 , \UART_TX/n61 , \UART_TX/n60 , \UART_TX/n59 ,
         \UART_TX/n58 , \UART_TX/n57 , \UART_TX/n56 , \UART_TX/n54 ,
         \UART_TX/n53 , \UART_TX/n52 , \UART_TX/n51 , \UART_TX/n50 ,
         \UART_TX/n49 , \UART_TX/n48 , \UART_TX/n47 , \UART_TX/n46 ,
         \UART_TX/n45 , \UART_TX/n44 , \UART_TX/n43 , \UART_TX/n42 ,
         \UART_TX/n41 , \UART_TX/n40 , \UART_TX/n39 , \UART_TX/n38 ,
         \UART_TX/n37 , \UART_TX/n36 , \UART_TX/n35 , \UART_TX/n34 ,
         \UART_TX/n33 , \UART_TX/n32 , \UART_TX/n31 , \UART_TX/n30 ,
         \UART_TX/n29 , \UART_TX/n28 , \UART_TX/n27 , \UART_TX/n26 ,
         \UART_TX/n25 , \UART_TX/n24 , \UART_TX/n23 , \UART_TX/n22 ,
         \UART_TX/n21 , \UART_TX/n20 , \UART_TX/n19 , \UART_TX/n18 ,
         \UART_TX/n17 , \UART_TX/n16 , \UART_TX/n15 , \UART_TX/n14 ,
         \UART_TX/n13 , \UART_TX/n12 , \UART_TX/n11 , \UART_TX/n10 ,
         \UART_TX/n9 , \UART_TX/n8 , \UART_TX/n7 , \UART_TX/n6 , \UART_TX/n5 ,
         \UART_TX/n4 , \UART_TX/n3 , \UART_TX/n2 , \UART_TX/n1 , \UART_TX/n93 ,
         \UART_TX/n92 , \UART_TX/n90 , \UART_TX/n89 , \UART_TX/n88 ,
         \UART_TX/n87 , \UART_TX/N127 , \UART_TX/iLast , \UART_TX/iTx2 ,
         \UART_TX/CState[0] , \UART_TX/CState[1] , \UART_TX/CState[2] ,
         \UART_TX/CState[3] , \UART_RX/n85 , \UART_RX/n84 , \UART_RX/n83 ,
         \UART_RX/n82 , \UART_RX/n81 , \UART_RX/n80 , \UART_RX/n79 ,
         \UART_RX/n78 , \UART_RX/n77 , \UART_RX/n76 , \UART_RX/n75 ,
         \UART_RX/n74 , \UART_RX/n73 , \UART_RX/n72 , \UART_RX/n70 ,
         \UART_RX/n69 , \UART_RX/n68 , \UART_RX/n67 , \UART_RX/n66 ,
         \UART_RX/n65 , \UART_RX/n64 , \UART_RX/n63 , \UART_RX/n62 ,
         \UART_RX/n61 , \UART_RX/n59 , \UART_RX/n58 , \UART_RX/n57 ,
         \UART_RX/n56 , \UART_RX/n55 , \UART_RX/n54 , \UART_RX/n53 ,
         \UART_RX/n52 , \UART_RX/n51 , \UART_RX/n50 , \UART_RX/n49 ,
         \UART_RX/n48 , \UART_RX/n47 , \UART_RX/n46 , \UART_RX/n45 ,
         \UART_RX/n44 , \UART_RX/n43 , \UART_RX/n42 , \UART_RX/n41 ,
         \UART_RX/n40 , \UART_RX/n39 , \UART_RX/n38 , \UART_RX/n37 ,
         \UART_RX/n36 , \UART_RX/n35 , \UART_RX/n34 , \UART_RX/n33 ,
         \UART_RX/n32 , \UART_RX/n31 , \UART_RX/n30 , \UART_RX/n29 ,
         \UART_RX/n28 , \UART_RX/n27 , \UART_RX/n26 , \UART_RX/n25 ,
         \UART_RX/n24 , \UART_RX/n23 , \UART_RX/n22 , \UART_RX/n21 ,
         \UART_RX/n20 , \UART_RX/n19 , \UART_RX/n18 , \UART_RX/n17 ,
         \UART_RX/n16 , \UART_RX/n15 , \UART_RX/n14 , \UART_RX/n13 ,
         \UART_RX/n12 , \UART_RX/n11 , \UART_RX/n10 , \UART_RX/n9 ,
         \UART_RX/n8 , \UART_RX/n7 , \UART_RX/n6 , \UART_RX/n5 , \UART_RX/n4 ,
         \UART_RX/n3 , \UART_RX/n2 , \UART_RX/n1 , \UART_RX/n117 ,
         \UART_RX/n116 , \UART_RX/n115 , \UART_RX/n114 , \UART_RX/n113 ,
         \UART_RX/n112 , \UART_RX/n111 , \UART_RX/n110 , \UART_RX/n109 ,
         \UART_RX/n108 , \UART_RX/n107 , \UART_RX/n106 , \UART_RX/n105 ,
         \UART_RX/N106 , \UART_RX/iParityReceived , \UART_RX/N75 ,
         \UART_RX/CState[0] , \UART_RX/CState[1] , \UART_RX/CState[2] ,
         \UART_RX/iDataCount[0] , \UART_RX/iDataCount[1] ,
         \UART_RX/iDataCount[2] , \UART_RX/iDataCount[3] ,
         \UART_RX/iBaudStepD , \UART_RX/iFStopBit , \UART_RX/iFSIN ,
         \UART_RX/iFilterClear , \UART_RX/iBaudStep , \UART_RX/iBaudCount[3] ,
         \UART_RX/RX_BRC/n23 , \UART_RX/RX_BRC/n22 , \UART_RX/RX_BRC/n21 ,
         \UART_RX/RX_BRC/n18 , \UART_RX/RX_BRC/n17 , \UART_RX/RX_BRC/n13 ,
         \UART_RX/RX_BRC/n12 , \UART_RX/RX_BRC/n9 , \UART_RX/RX_BRC/n8 ,
         \UART_RX/RX_BRC/n7 , \UART_RX/RX_BRC/n6 , \UART_RX/RX_BRC/n5 ,
         \UART_RX/RX_BRC/n1 , \UART_RX/RX_BRC/n30 , \UART_RX/RX_BRC/n29 ,
         \UART_RX/RX_BRC/n28 , \UART_RX/RX_BRC/n27 , \UART_RX/RX_BRC/n26 ,
         \UART_RX/RX_BRC/Q[0] , \UART_RX/RX_BRC/Q[1] , \UART_RX/RX_BRC/Q[2] ,
         \UART_RX/RX_MVF/n18 , \UART_RX/RX_MVF/n17 , \UART_RX/RX_MVF/n16 ,
         \UART_RX/RX_MVF/n15 , \UART_RX/RX_MVF/n14 , \UART_RX/RX_MVF/n13 ,
         \UART_RX/RX_MVF/n12 , \UART_RX/RX_MVF/n11 , \UART_RX/RX_MVF/n10 ,
         \UART_RX/RX_MVF/n9 , \UART_RX/RX_MVF/n8 , \UART_RX/RX_MVF/n7 ,
         \UART_RX/RX_MVF/n6 , \UART_RX/RX_MVF/n5 , \UART_RX/RX_MVF/n3 ,
         \UART_RX/RX_MVF/n2 , \UART_RX/RX_MVF/n1 , \UART_RX/RX_MVF/n26 ,
         \UART_RX/RX_MVF/n24 , \UART_RX/RX_MVF/n23 , \UART_RX/RX_MVF/n22 ,
         \UART_RX/RX_MVF/n21 , \UART_RX/RX_MVF/iCounter[0] ,
         \UART_RX/RX_MVF/iCounter[1] , \UART_RX/RX_MVF/iCounter[2] ,
         \UART_RX/RX_MVF/iCounter[3] , \UART_RX/RX_IFSB/n18 ,
         \UART_RX/RX_IFSB/n17 , \UART_RX/RX_IFSB/n16 , \UART_RX/RX_IFSB/n15 ,
         \UART_RX/RX_IFSB/n14 , \UART_RX/RX_IFSB/n13 , \UART_RX/RX_IFSB/n12 ,
         \UART_RX/RX_IFSB/n11 , \UART_RX/RX_IFSB/n10 , \UART_RX/RX_IFSB/n9 ,
         \UART_RX/RX_IFSB/n8 , \UART_RX/RX_IFSB/n7 , \UART_RX/RX_IFSB/n6 ,
         \UART_RX/RX_IFSB/n5 , \UART_RX/RX_IFSB/n4 , \UART_RX/RX_IFSB/n3 ,
         \UART_RX/RX_IFSB/n2 , \UART_RX/RX_IFSB/n1 , \UART_RX/RX_IFSB/n33 ,
         \UART_RX/RX_IFSB/n32 , \UART_RX/RX_IFSB/n31 , \UART_RX/RX_IFSB/n30 ,
         \UART_RX/RX_IFSB/iCount[0] , \UART_RX/RX_IFSB/iCount[1] ,
         \UART_RX/RX_IFSB/iCount[2] , \r108/n1 , n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689;
  wire   [2:0] iA;
  wire   [7:0] iDIN;
  wire   [7:0] iDLL;
  wire   [7:0] iDLM;
  wire   [3:0] iIER;
  wire   [7:0] iLSR;
  wire   [7:0] iMSR;
  wire   [3:0] iIIR;
  wire   [5:0] iTimeoutCount;
  wire   [1:0] iFCR_RXTrigger;
  wire   [2:1] iFCR;
  wire   [7:0] iLCR;
  wire   [5:0] iMCR;
  wire   [6:0] iFECounter;
  wire   [10:0] iRXFIFOQ;
  wire   [10:0] iRXFIFOD;
  wire   [7:0] iSCR;
  wire   [7:0] iTXFIFOQ;
  wire   [5:1] iRXFIFOUsage;
  wire   [7:0] iTSR;
  wire   [7:0] iRXData;
  wire   [1:0] State;
  wire   [15:2] \UART_BG16/add_54/carry ;
  wire   [6:2] \UART_TXFF/add_73/carry ;
  wire   [6:2] \UART_TXFF/add_77/carry ;
  wire   [6:2] \UART_RXFF/add_73/carry ;
  wire   [6:2] \UART_RXFF/add_77/carry ;
  wire   [2:0] \UART_RX/NState ;
  wire   [6:0] \r108/carry ;

  notech_reg \iDIN_reg[7]  ( .D(DIN[7]), .CP(CLK), .CD(n416), .Q(iDIN[7]) );
  notech_reg \iDIN_reg[6]  ( .D(DIN[6]), .CP(CLK), .CD(n420), .Q(iDIN[6]) );
  notech_reg \iDIN_reg[5]  ( .D(DIN[5]), .CP(CLK), .CD(n419), .Q(iDIN[5]) );
  notech_reg \iDIN_reg[4]  ( .D(DIN[4]), .CP(CLK), .CD(n415), .Q(iDIN[4]) );
  notech_reg \iDIN_reg[3]  ( .D(DIN[3]), .CP(CLK), .CD(n420), .Q(iDIN[3]) );
  notech_reg \iDIN_reg[2]  ( .D(DIN[2]), .CP(CLK), .CD(n420), .Q(iDIN[2]) );
  notech_reg \iDIN_reg[1]  ( .D(DIN[1]), .CP(CLK), .CD(n415), .Q(iDIN[1]) );
  notech_reg \iDIN_reg[0]  ( .D(DIN[0]), .CP(CLK), .CD(n416), .Q(iDIN[0]) );
  notech_reg \iA_reg[2]  ( .D(A[2]), .CP(CLK), .CD(n416), .Q(iA[2]) );
  notech_reg \iA_reg[1]  ( .D(A[1]), .CP(CLK), .CD(n415), .Q(iA[1]) );
  notech_reg \iA_reg[0]  ( .D(A[0]), .CP(CLK), .CD(n420), .Q(iA[0]) );
  notech_reg \iFCR_RXTrigger_reg[1]  ( .D(n369), .CP(CLK), .CD(n420), .Q(
        iFCR_RXTrigger[1]) );
  notech_reg \iFCR_RXTrigger_reg[0]  ( .D(n368), .CP(CLK), .CD(n419), .Q(
        iFCR_RXTrigger[0]) );
  notech_reg iFCR_FIFOEnable_reg ( .D(n367), .CP(CLK), .CD(n416), .Q(iIIR_6)
         );
  notech_reg iFCR_RXFIFOReset_reg ( .D(N94), .CP(CLK), .CD(n418), .Q(iFCR[1])
         );
  notech_reg iFCR_TXFIFOReset_reg ( .D(N95), .CP(CLK), .CD(n417), .Q(iFCR[2])
         );
  notech_reg \iLCR_reg[7]  ( .D(n366), .CP(CLK), .CD(n417), .Q(iLCR[7]) );
  notech_reg \iDLL_reg[7]  ( .D(n365), .CP(CLK), .CD(n416), .Q(iDLL[7]) );
  notech_reg \iDLL_reg[6]  ( .D(n364), .CP(CLK), .CD(n419), .Q(iDLL[6]) );
  notech_reg \iDLL_reg[5]  ( .D(n363), .CP(CLK), .CD(n420), .Q(iDLL[5]) );
  notech_reg \iDLL_reg[4]  ( .D(n362), .CP(CLK), .CD(n418), .Q(iDLL[4]) );
  notech_reg \iDLL_reg[3]  ( .D(n361), .CP(CLK), .CD(n416), .Q(iDLL[3]) );
  notech_reg \iDLL_reg[2]  ( .D(n360), .CP(CLK), .CD(n418), .Q(iDLL[2]) );
  notech_reg \iDLL_reg[1]  ( .D(n359), .CP(CLK), .CD(n419), .Q(iDLL[1]) );
  notech_reg \iDLL_reg[0]  ( .D(n358), .CP(CLK), .CD(n415), .Q(iDLL[0]) );
  notech_reg \iDLM_reg[7]  ( .D(n357), .CP(CLK), .CD(n420), .Q(iDLM[7]) );
  notech_reg \iDLM_reg[6]  ( .D(n356), .CP(CLK), .CD(n417), .Q(iDLM[6]) );
  notech_reg \iDLM_reg[5]  ( .D(n355), .CP(CLK), .CD(n415), .Q(iDLM[5]) );
  notech_reg \iDLM_reg[4]  ( .D(n354), .CP(CLK), .CD(n418), .Q(iDLM[4]) );
  notech_reg \iDLM_reg[3]  ( .D(n353), .CP(CLK), .CD(n415), .Q(iDLM[3]) );
  notech_reg \iDLM_reg[2]  ( .D(n352), .CP(CLK), .CD(n416), .Q(iDLM[2]) );
  notech_reg \iDLM_reg[1]  ( .D(n351), .CP(CLK), .CD(n420), .Q(iDLM[1]) );
  notech_reg \iDLM_reg[0]  ( .D(n350), .CP(CLK), .CD(n415), .Q(iDLM[0]) );
  notech_reg iFCR_FIFO64E_reg ( .D(n412), .CP(CLK), .CD(n420), .Q(iFCR_5) );
  notech_reg \iIER_reg[3]  ( .D(n349), .CP(CLK), .CD(n420), .Q(iIER[3]) );
  notech_reg \iIER_reg[2]  ( .D(n348), .CP(CLK), .CD(n417), .Q(iIER[2]) );
  notech_reg \iIER_reg[1]  ( .D(n347), .CP(CLK), .CD(n419), .Q(iIER[1]) );
  notech_reg \iIER_reg[0]  ( .D(n346), .CP(CLK), .CD(n417), .Q(iIER[0]) );
  notech_reg \iLCR_reg[6]  ( .D(n345), .CP(CLK), .CD(n416), .Q(iLCR[6]) );
  notech_reg \iLCR_reg[5]  ( .D(n344), .CP(CLK), .CD(n418), .Q(iLCR[5]) );
  notech_reg \iLCR_reg[4]  ( .D(n343), .CP(CLK), .CD(n417), .Q(iLCR[4]) );
  notech_reg \iLCR_reg[3]  ( .D(n342), .CP(CLK), .CD(n416), .Q(iLCR[3]) );
  notech_reg \iLCR_reg[2]  ( .D(n341), .CP(CLK), .CD(n419), .Q(iLCR[2]) );
  notech_reg \iLCR_reg[1]  ( .D(n340), .CP(CLK), .CD(n419), .Q(iLCR[1]) );
  notech_reg \iLCR_reg[0]  ( .D(n339), .CP(CLK), .CD(n418), .Q(iLCR[0]) );
  notech_reg \iMCR_reg[5]  ( .D(n338), .CP(CLK), .CD(n417), .Q(iMCR[5]) );
  notech_reg \iMCR_reg[4]  ( .D(n337), .CP(CLK), .CD(n417), .Q(iMCR[4]) );
  notech_reg \iMCR_reg[3]  ( .D(n336), .CP(CLK), .CD(n420), .Q(iMCR[3]) );
  notech_reg \iMCR_reg[2]  ( .D(n335), .CP(CLK), .CD(n417), .Q(iMCR[2]) );
  notech_reg \iMCR_reg[1]  ( .D(n334), .CP(CLK), .CD(n418), .Q(iMCR[1]) );
  notech_reg \iMCR_reg[0]  ( .D(n333), .CP(CLK), .CD(n415), .Q(iMCR[0]) );
  notech_reg iMSR_dDCD_reg ( .D(n411), .CP(CLK), .CD(n419), .Q(iMSR[3]) );
  notech_reg iMSR_dDSR_reg ( .D(n410), .CP(CLK), .CD(n415), .Q(iMSR[1]) );
  notech_reg iMSR_TERI_reg ( .D(n409), .CP(CLK), .CD(n417), .Q(iMSR[2]) );
  notech_reg \iSCR_reg[7]  ( .D(n332), .CP(CLK), .CD(n416), .Q(iSCR[7]) );
  notech_reg \iSCR_reg[6]  ( .D(n331), .CP(CLK), .CD(n419), .Q(iSCR[6]) );
  notech_reg \iSCR_reg[5]  ( .D(n330), .CP(CLK), .CD(n418), .Q(iSCR[5]) );
  notech_reg \iSCR_reg[4]  ( .D(n329), .CP(CLK), .CD(n415), .Q(iSCR[4]) );
  notech_reg \iSCR_reg[3]  ( .D(n328), .CP(CLK), .CD(n415), .Q(iSCR[3]) );
  notech_reg \iSCR_reg[2]  ( .D(n327), .CP(CLK), .CD(n419), .Q(iSCR[2]) );
  notech_reg \iSCR_reg[1]  ( .D(n326), .CP(CLK), .CD(n416), .Q(iSCR[1]) );
  notech_reg \iSCR_reg[0]  ( .D(n325), .CP(CLK), .CD(n417), .Q(iSCR[0]) );
  notech_reg iRTS_reg ( .D(n408), .CP(CLK), .CD(n418), .Q(iRTS) );
  notech_reg iMSR_dCTS_reg ( .D(n407), .CP(CLK), .CD(n416), .Q(iMSR[0]) );
  notech_reg \State_reg[0]  ( .D(N181), .CP(CLK), .CD(n415), .Q(State[0]) );
  notech_reg iTXFIFORead_reg ( .D(n679), .CP(CLK), .CD(n416), .Q(iTXFIFORead)
         );
  notech_reg \iTSR_reg[7]  ( .D(n324), .CP(CLK), .CD(n415), .Q(iTSR[7]) );
  notech_reg \iTSR_reg[6]  ( .D(n323), .CP(CLK), .CD(n419), .Q(iTSR[6]) );
  notech_reg \iTSR_reg[5]  ( .D(n322), .CP(CLK), .CD(n418), .Q(iTSR[5]) );
  notech_reg \iTSR_reg[4]  ( .D(n321), .CP(CLK), .CD(n417), .Q(iTSR[4]) );
  notech_reg \iTSR_reg[3]  ( .D(n320), .CP(CLK), .CD(n418), .Q(iTSR[3]) );
  notech_reg \iTSR_reg[2]  ( .D(n319), .CP(CLK), .CD(n420), .Q(iTSR[2]) );
  notech_reg \iTSR_reg[1]  ( .D(n318), .CP(CLK), .CD(n419), .Q(iTSR[1]) );
  notech_reg \iTSR_reg[0]  ( .D(n317), .CP(CLK), .CD(n416), .Q(iTSR[0]) );
  notech_reg \State_reg[1]  ( .D(N182), .CP(CLK), .CD(n419), .Q(State[1]) );
  notech_reg iTXRunning_reg ( .D(n414), .CP(CLK), .CD(n416), .Q(iTXRunning) );
  notech_reg iTXStart_reg ( .D(N183), .CP(CLK), .CD(n418), .Q(iTXStart) );
  notech_reg iRXFIFOClear_reg ( .D(N190), .CP(CLK), .CD(n420), .Q(iRXFIFOClear) );
  notech_reg State_reg2 ( .D(n673), .CP(CLK), .CD(n420), .Q(State_snps_wire)
         );
  notech_reg \iRXFIFOD_reg[0]  ( .D(n406), .CP(CLK), .CD(n420), .Q(iRXFIFOD[0]) );
  notech_reg \iRXFIFOD_reg[1]  ( .D(n405), .CP(CLK), .CD(n419), .Q(iRXFIFOD[1]) );
  notech_reg \iRXFIFOD_reg[2]  ( .D(n404), .CP(CLK), .CD(n416), .Q(iRXFIFOD[2]) );
  notech_reg \iRXFIFOD_reg[3]  ( .D(n403), .CP(CLK), .CD(n418), .Q(iRXFIFOD[3]) );
  notech_reg \iRXFIFOD_reg[4]  ( .D(n402), .CP(CLK), .CD(n419), .Q(iRXFIFOD[4]) );
  notech_reg \iRXFIFOD_reg[5]  ( .D(n401), .CP(CLK), .CD(n418), .Q(iRXFIFOD[5]) );
  notech_reg \iRXFIFOD_reg[6]  ( .D(n400), .CP(CLK), .CD(n417), .Q(iRXFIFOD[6]) );
  notech_reg \iRXFIFOD_reg[7]  ( .D(n399), .CP(CLK), .CD(n415), .Q(iRXFIFOD[7]) );
  notech_reg \iRXFIFOD_reg[10]  ( .D(n398), .CP(CLK), .CD(n420), .Q(
        iRXFIFOD[10]) );
  notech_reg \iRXFIFOD_reg[9]  ( .D(n397), .CP(CLK), .CD(n417), .Q(iRXFIFOD[9]) );
  notech_reg \iRXFIFOD_reg[8]  ( .D(n396), .CP(CLK), .CD(n419), .Q(iRXFIFOD[8]) );
  notech_reg iRXFIFOWrite_reg ( .D(N191), .CP(CLK), .CD(n415), .Q(iRXFIFOWrite) );
  notech_reg iLSR_OE_reg ( .D(n395), .CP(CLK), .CD(n418), .Q(iLSR[1]) );
  notech_reg \iTimeoutCount_reg[5]  ( .D(n394), .CP(CLK), .CD(n417), .Q(
        iTimeoutCount[5]) );
  notech_reg \iTimeoutCount_reg[0]  ( .D(n393), .CP(CLK), .CD(n415), .Q(
        iTimeoutCount[0]) );
  notech_reg \iTimeoutCount_reg[1]  ( .D(n392), .CP(CLK), .CD(n416), .Q(
        iTimeoutCount[1]) );
  notech_reg \iTimeoutCount_reg[2]  ( .D(n391), .CP(CLK), .CD(n419), .Q(
        iTimeoutCount[2]) );
  notech_reg \iTimeoutCount_reg[3]  ( .D(n390), .CP(CLK), .CD(n419), .Q(
        iTimeoutCount[3]) );
  notech_reg \iTimeoutCount_reg[4]  ( .D(n389), .CP(CLK), .CD(n418), .Q(
        iTimeoutCount[4]) );
  notech_reg iCharTimeout_reg ( .D(n388), .CP(CLK), .CD(n420), .Q(iCharTimeout) );
  notech_reg iLSR_PE_reg ( .D(n387), .CP(CLK), .CD(n417), .Q(iLSR[2]) );
  notech_reg iLSR_FE_reg ( .D(n386), .CP(CLK), .CD(n415), .Q(iLSR[3]) );
  notech_reg iLSR_BI_reg ( .D(n377), .CP(CLK), .CD(n417), .Q(iLSR[4]) );
  notech_reg iTHRInterrupt_reg ( .D(n376), .CP(CLK), .CD(n420), .Q(
        iTHRInterrupt) );
  notech_reg \iFECounter_reg[6]  ( .D(n379), .CP(CLK), .CD(n418), .Q(
        iFECounter[6]) );
  notech_reg \iFECounter_reg[0]  ( .D(n385), .CP(CLK), .CD(n420), .Q(
        iFECounter[0]) );
  notech_reg \iFECounter_reg[1]  ( .D(n384), .CP(CLK), .CD(n416), .Q(
        iFECounter[1]) );
  notech_reg \iFECounter_reg[2]  ( .D(n383), .CP(CLK), .CD(n415), .Q(
        iFECounter[2]) );
  notech_reg \iFECounter_reg[3]  ( .D(n382), .CP(CLK), .CD(n415), .Q(
        iFECounter[3]) );
  notech_reg \iFECounter_reg[4]  ( .D(n381), .CP(CLK), .CD(n417), .Q(
        iFECounter[4]) );
  notech_reg \iFECounter_reg[5]  ( .D(n380), .CP(CLK), .CD(n417), .Q(
        iFECounter[5]) );
  notech_reg iLSR_FIFOERR_reg ( .D(n378), .CP(CLK), .CD(1'b1), .Q(iLSR_FIFOERR) );
  notech_reg_set SOUT_reg ( .D(N202), .CP(CLK), .SD(n418), .Q(SOUT) );
  notech_reg_set DDIS_reg ( .D(N197), .CP(CLK), .SD(n417), .Q(DDIS) );
  notech_reg_set BAUDOUTN_reg ( .D(n677), .CP(CLK), .SD(n419), .Q(BAUDOUTN) );
  notech_reg_set OUT1N_reg ( .D(N198), .CP(CLK), .SD(n418), .Q(OUT1N) );
  notech_reg_set OUT2N_reg ( .D(N199), .CP(CLK), .SD(n415), .Q(OUT2N) );
  notech_reg_set RTSN_reg ( .D(N200), .CP(CLK), .SD(n416), .Q(RTSN) );
  notech_reg_set DTRN_reg ( .D(N201), .CP(CLK), .SD(n416), .Q(DTRN) );
  notech_inv U447 ( .A(RST), .Z(n415) );
  notech_inv U448 ( .A(RST), .Z(n416) );
  notech_inv U449 ( .A(RST), .Z(n417) );
  notech_inv U450 ( .A(RST), .Z(n418) );
  notech_inv U451 ( .A(RST), .Z(n419) );
  notech_inv U452 ( .A(RST), .Z(n420) );
  notech_inv U453 ( .A(iBaudtick16x), .Z(n677) );
  notech_mux2 U454 ( .A(iFCR_5), .B(iDIN[5]), .S(n421), .Z(n412) );
  notech_and2 U455 ( .A(n422), .B(iLCR[7]), .Z(n421) );
  notech_nao3 U456 ( .C(iDCDnFE), .A(n685), .B(n424), .Z(n411) );
  notech_or2 U457 ( .A(n425), .B(n426), .Z(n424) );
  notech_nao3 U459 ( .C(iDSRnFE), .A(n684), .B(n428), .Z(n410) );
  notech_or2 U460 ( .A(n425), .B(n429), .Z(n428) );
  notech_or2 U462 ( .A(n430), .B(iRInFE), .Z(n409) );
  notech_nor2 U463 ( .A(n425), .B(n431), .Z(n430) );
  notech_and2 U464 ( .A(n432), .B(iMCR[1]), .Z(n408) );
  notech_or2 U465 ( .A(n433), .B(n434), .Z(n432) );
  notech_and2 U466 ( .A(n435), .B(n436), .Z(n433) );
  notech_nand2 U467 ( .A(n437), .B(n438), .Z(n436) );
  notech_nao3 U468 ( .C(iCTSnFE), .A(n683), .B(n440), .Z(n407) );
  notech_or2 U469 ( .A(n425), .B(n441), .Z(n440) );
  notech_and4 U470 ( .A(iA[2]), .B(iReadFE), .C(n442), .D(iA[1]), .Z(n425) );
  notech_mux2 U472 ( .A(iRXFIFOD[0]), .B(iRXData[0]), .S(n673), .Z(n406) );
  notech_mux2 U473 ( .A(iRXFIFOD[1]), .B(iRXData[1]), .S(n673), .Z(n405) );
  notech_mux2 U474 ( .A(iRXFIFOD[2]), .B(iRXData[2]), .S(n673), .Z(n404) );
  notech_mux2 U475 ( .A(iRXFIFOD[3]), .B(iRXData[3]), .S(n673), .Z(n403) );
  notech_mux2 U476 ( .A(iRXFIFOD[4]), .B(iRXData[4]), .S(n673), .Z(n402) );
  notech_mux2 U477 ( .A(iRXFIFOD[5]), .B(iRXData[5]), .S(n673), .Z(n401) );
  notech_mux2 U478 ( .A(iRXFIFOD[6]), .B(iRXData[6]), .S(n673), .Z(n400) );
  notech_mux2 U479 ( .A(iRXFIFOD[7]), .B(iRXData[7]), .S(n673), .Z(n399) );
  notech_mux2 U480 ( .A(iRXFIFOD[10]), .B(iRXBI), .S(n673), .Z(n398) );
  notech_mux2 U481 ( .A(iRXFIFOD[9]), .B(iRXFE), .S(n673), .Z(n397) );
  notech_mux2 U482 ( .A(iRXFIFOD[8]), .B(iRXPE), .S(n673), .Z(n396) );
  notech_nao4 U483 ( .A(n443), .B(n444), .C(n680), .D(n446), .Z(n395) );
  notech_inv U484 ( .A(n447), .Z(n446) );
  notech_mux2 U485 ( .A(n448), .B(n676), .S(n449), .Z(n447) );
  notech_inv U486 ( .A(n450), .Z(n676) );
  notech_nao4 U487 ( .A(n451), .B(n452), .C(n453), .D(n454), .Z(n394) );
  notech_mux2 U488 ( .A(n455), .B(n456), .S(n457), .Z(n393) );
  notech_mux2 U489 ( .A(n458), .B(n459), .S(iTimeoutCount[1]), .Z(n392) );
  notech_nor2 U490 ( .A(n460), .B(n457), .Z(n458) );
  notech_inv U491 ( .A(iTimeoutCount[0]), .Z(n457) );
  notech_mux2 U492 ( .A(n461), .B(n462), .S(iTimeoutCount[2]), .Z(n391) );
  notech_or2 U493 ( .A(n459), .B(n463), .Z(n462) );
  notech_nor2 U494 ( .A(n460), .B(iTimeoutCount[1]), .Z(n463) );
  notech_or2 U495 ( .A(n464), .B(n455), .Z(n459) );
  notech_nor2 U496 ( .A(n460), .B(iTimeoutCount[0]), .Z(n464) );
  notech_ao3 U497 ( .A(iTimeoutCount[1]), .B(iTimeoutCount[0]), .C(n460), .Z(
        n461) );
  notech_mux2 U498 ( .A(n465), .B(n466), .S(iTimeoutCount[3]), .Z(n390) );
  notech_and2 U499 ( .A(n456), .B(n467), .Z(n465) );
  notech_inv U500 ( .A(n460), .Z(n456) );
  notech_inv U501 ( .A(n468), .Z(n389) );
  notech_mux2 U502 ( .A(n451), .B(n453), .S(n454), .Z(n468) );
  notech_inv U503 ( .A(iTimeoutCount[4]), .Z(n454) );
  notech_nao3 U504 ( .C(n460), .A(iTimeoutCount[3]), .B(n467), .Z(n453) );
  notech_nor2 U505 ( .A(n466), .B(n469), .Z(n451) );
  notech_nor2 U506 ( .A(n460), .B(iTimeoutCount[3]), .Z(n469) );
  notech_or2 U507 ( .A(n470), .B(n455), .Z(n466) );
  notech_nor2 U508 ( .A(n460), .B(n467), .Z(n470) );
  notech_and3 U509 ( .A(iTimeoutCount[2]), .B(iTimeoutCount[1]), .C(
        iTimeoutCount[0]), .Z(n467) );
  notech_or2 U510 ( .A(n455), .B(n471), .Z(n460) );
  notech_nor2 U511 ( .A(n471), .B(n472), .Z(n455) );
  notech_and2 U512 ( .A(iBaudtick2x), .B(n452), .Z(n472) );
  notech_inv U513 ( .A(iTimeoutCount[5]), .Z(n452) );
  notech_nao3 U514 ( .C(n371), .A(n438), .B(\UART_RXFF/n441 ), .Z(n471) );
  notech_ao3 U515 ( .A(n474), .B(iIIR_6), .C(n371), .Z(n388) );
  notech_or2 U516 ( .A(iCharTimeout), .B(iTimeoutCount[5]), .Z(n474) );
  notech_or2 U517 ( .A(n475), .B(iPERE), .Z(n387) );
  notech_nor2 U518 ( .A(n443), .B(n476), .Z(n475) );
  notech_or2 U519 ( .A(n477), .B(iFERE), .Z(n386) );
  notech_nor2 U520 ( .A(n443), .B(n478), .Z(n477) );
  notech_inv U521 ( .A(n479), .Z(n385) );
  notech_mux2 U522 ( .A(n480), .B(n481), .S(iFECounter[0]), .Z(n479) );
  notech_nao4 U523 ( .A(n481), .B(n482), .C(n480), .D(n483), .Z(n384) );
  notech_inv U524 ( .A(N130), .Z(n483) );
  notech_inv U525 ( .A(iFECounter[1]), .Z(n482) );
  notech_nao4 U526 ( .A(n481), .B(n484), .C(n480), .D(n485), .Z(n383) );
  notech_inv U527 ( .A(N131), .Z(n485) );
  notech_inv U528 ( .A(iFECounter[2]), .Z(n484) );
  notech_nao4 U529 ( .A(n481), .B(n486), .C(n480), .D(n487), .Z(n382) );
  notech_inv U530 ( .A(N132), .Z(n487) );
  notech_inv U531 ( .A(iFECounter[3]), .Z(n486) );
  notech_nao4 U532 ( .A(n481), .B(n488), .C(n480), .D(n489), .Z(n381) );
  notech_inv U533 ( .A(N133), .Z(n489) );
  notech_inv U534 ( .A(iFECounter[4]), .Z(n488) );
  notech_nao4 U535 ( .A(n481), .B(n490), .C(n480), .D(n491), .Z(n380) );
  notech_inv U536 ( .A(N134), .Z(n491) );
  notech_inv U537 ( .A(iFECounter[5]), .Z(n490) );
  notech_nao4 U538 ( .A(n481), .B(n492), .C(n480), .D(n493), .Z(n379) );
  notech_inv U539 ( .A(N135), .Z(n493) );
  notech_nand2 U540 ( .A(n481), .B(\UART_RXFF/n308 ), .Z(n480) );
  notech_inv U541 ( .A(iFECounter[6]), .Z(n492) );
  notech_nand3 U542 ( .A(\UART_RXFF/n308 ), .B(\U3/U1/Z_0 ), .C(n495), .Z(n481) );
  notech_or4 U543 ( .A(n496), .B(n497), .C(iRXFIFOEmpty), .D(n498), .Z(n495)
         );
  notech_nor2 U544 ( .A(n499), .B(\UART_RXFF/n441 ), .Z(n497) );
  notech_mux2 U547 ( .A(iLSR_FIFOERR), .B(n500), .S(n501), .Z(n378) );
  notech_nor2 U548 ( .A(n502), .B(RST), .Z(n501) );
  notech_nor2 U549 ( .A(n503), .B(n500), .Z(n502) );
  notech_ao3 U550 ( .A(n504), .B(n505), .C(n674), .Z(n503) );
  notech_and2 U551 ( .A(iRXFIFOQ[10]), .B(n438), .Z(n674) );
  notech_inv U552 ( .A(N146), .Z(n505) );
  notech_inv U553 ( .A(n675), .Z(n504) );
  notech_and2 U554 ( .A(iRXFIFOQ[9]), .B(n438), .Z(n675) );
  notech_or2 U555 ( .A(n506), .B(iBIRE), .Z(n377) );
  notech_nor2 U556 ( .A(n443), .B(n507), .Z(n506) );
  notech_and4 U557 ( .A(iReadFE), .B(iA[0]), .C(n508), .D(iA[2]), .Z(n443) );
  notech_or4 U558 ( .A(n509), .B(n510), .C(iLSR_THRERE), .D(iFCR[2]), .Z(n376)
         );
  notech_and2 U559 ( .A(iTHRInterrupt), .B(n511), .Z(n510) );
  notech_nao3 U560 ( .C(iA[0]), .A(n512), .B(n513), .Z(n511) );
  notech_mux2 U561 ( .A(n514), .B(n515), .S(n508), .Z(n513) );
  notech_and2 U562 ( .A(n516), .B(iWriteFE), .Z(n515) );
  notech_and4 U563 ( .A(iIIR[1]), .B(iReadFE), .C(n517), .D(n518), .Z(n514) );
  notech_ao3 U564 ( .A(iDIN[1]), .B(n519), .C(n520), .Z(n509) );
  notech_ao3 U565 ( .A(iReadFE), .B(n521), .C(iA[0]), .Z(n371) );
  notech_mux2 U566 ( .A(iFCR_RXTrigger[1]), .B(iDIN[7]), .S(n422), .Z(n369) );
  notech_mux2 U567 ( .A(iFCR_RXTrigger[0]), .B(iDIN[6]), .S(n422), .Z(n368) );
  notech_mux2 U568 ( .A(iIIR_6), .B(iDIN[0]), .S(n422), .Z(n367) );
  notech_mux2 U569 ( .A(iLCR[7]), .B(iDIN[7]), .S(n522), .Z(n366) );
  notech_mux2 U570 ( .A(iDLL[7]), .B(iDIN[7]), .S(n523), .Z(n365) );
  notech_mux2 U571 ( .A(iDLL[6]), .B(iDIN[6]), .S(n523), .Z(n364) );
  notech_mux2 U572 ( .A(iDLL[5]), .B(iDIN[5]), .S(n523), .Z(n363) );
  notech_mux2 U573 ( .A(iDLL[4]), .B(iDIN[4]), .S(n523), .Z(n362) );
  notech_mux2 U574 ( .A(iDLL[3]), .B(iDIN[3]), .S(n523), .Z(n361) );
  notech_mux2 U575 ( .A(iDLL[2]), .B(iDIN[2]), .S(n523), .Z(n360) );
  notech_mux2 U576 ( .A(iDLL[1]), .B(iDIN[1]), .S(n523), .Z(n359) );
  notech_mux2 U577 ( .A(iDLL[0]), .B(iDIN[0]), .S(n523), .Z(n358) );
  notech_and2 U578 ( .A(n524), .B(n442), .Z(n523) );
  notech_mux2 U579 ( .A(iDLM[7]), .B(iDIN[7]), .S(n525), .Z(n357) );
  notech_mux2 U580 ( .A(iDLM[6]), .B(iDIN[6]), .S(n525), .Z(n356) );
  notech_mux2 U581 ( .A(iDLM[5]), .B(iDIN[5]), .S(n525), .Z(n355) );
  notech_mux2 U582 ( .A(iDLM[4]), .B(iDIN[4]), .S(n525), .Z(n354) );
  notech_mux2 U583 ( .A(iDLM[3]), .B(iDIN[3]), .S(n525), .Z(n353) );
  notech_mux2 U584 ( .A(iDLM[2]), .B(iDIN[2]), .S(n525), .Z(n352) );
  notech_mux2 U585 ( .A(iDLM[1]), .B(iDIN[1]), .S(n525), .Z(n351) );
  notech_mux2 U586 ( .A(iDLM[0]), .B(iDIN[0]), .S(n525), .Z(n350) );
  notech_and2 U587 ( .A(n524), .B(iA[0]), .Z(n525) );
  notech_and4 U588 ( .A(iWriteFE), .B(iLCR[7]), .C(n512), .D(n508), .Z(n524)
         );
  notech_mux2 U589 ( .A(iIER[3]), .B(iDIN[3]), .S(n519), .Z(n349) );
  notech_mux2 U590 ( .A(iIER[2]), .B(iDIN[2]), .S(n519), .Z(n348) );
  notech_mux2 U591 ( .A(iIER[1]), .B(iDIN[1]), .S(n519), .Z(n347) );
  notech_mux2 U592 ( .A(iIER[0]), .B(iDIN[0]), .S(n519), .Z(n346) );
  notech_and3 U593 ( .A(n521), .B(iWriteFE), .C(iA[0]), .Z(n519) );
  notech_mux2 U594 ( .A(iLCR[6]), .B(iDIN[6]), .S(n522), .Z(n345) );
  notech_mux2 U595 ( .A(iLCR[5]), .B(iDIN[5]), .S(n522), .Z(n344) );
  notech_mux2 U596 ( .A(iLCR[4]), .B(iDIN[4]), .S(n522), .Z(n343) );
  notech_mux2 U597 ( .A(iLCR[3]), .B(iDIN[3]), .S(n522), .Z(n342) );
  notech_mux2 U598 ( .A(iLCR[2]), .B(iDIN[2]), .S(n522), .Z(n341) );
  notech_mux2 U599 ( .A(iLCR[1]), .B(iDIN[1]), .S(n522), .Z(n340) );
  notech_mux2 U600 ( .A(iLCR[0]), .B(iDIN[0]), .S(n522), .Z(n339) );
  notech_and2 U601 ( .A(n526), .B(n512), .Z(n522) );
  notech_mux2 U602 ( .A(iMCR[5]), .B(iDIN[5]), .S(n527), .Z(n338) );
  notech_mux2 U603 ( .A(iMCR[4]), .B(iDIN[4]), .S(n527), .Z(n337) );
  notech_mux2 U604 ( .A(iMCR[3]), .B(iDIN[3]), .S(n527), .Z(n336) );
  notech_mux2 U605 ( .A(iMCR[2]), .B(iDIN[2]), .S(n527), .Z(n335) );
  notech_mux2 U606 ( .A(iMCR[1]), .B(iDIN[1]), .S(n527), .Z(n334) );
  notech_mux2 U607 ( .A(iMCR[0]), .B(iDIN[0]), .S(n527), .Z(n333) );
  notech_and3 U608 ( .A(n528), .B(n508), .C(iA[2]), .Z(n527) );
  notech_mux2 U609 ( .A(iSCR[7]), .B(iDIN[7]), .S(n529), .Z(n332) );
  notech_mux2 U610 ( .A(iSCR[6]), .B(iDIN[6]), .S(n529), .Z(n331) );
  notech_mux2 U611 ( .A(iSCR[5]), .B(iDIN[5]), .S(n529), .Z(n330) );
  notech_mux2 U612 ( .A(iSCR[4]), .B(iDIN[4]), .S(n529), .Z(n329) );
  notech_mux2 U613 ( .A(iSCR[3]), .B(iDIN[3]), .S(n529), .Z(n328) );
  notech_mux2 U614 ( .A(iSCR[2]), .B(iDIN[2]), .S(n529), .Z(n327) );
  notech_mux2 U615 ( .A(iSCR[1]), .B(iDIN[1]), .S(n529), .Z(n326) );
  notech_mux2 U616 ( .A(iSCR[0]), .B(iDIN[0]), .S(n529), .Z(n325) );
  notech_and2 U617 ( .A(n526), .B(iA[2]), .Z(n529) );
  notech_and3 U618 ( .A(iA[1]), .B(iWriteFE), .C(iA[0]), .Z(n526) );
  notech_mux2 U619 ( .A(iTSR[7]), .B(iTXFIFOQ[7]), .S(n679), .Z(n324) );
  notech_mux2 U620 ( .A(iTSR[6]), .B(iTXFIFOQ[6]), .S(n679), .Z(n323) );
  notech_mux2 U621 ( .A(iTSR[5]), .B(iTXFIFOQ[5]), .S(n679), .Z(n322) );
  notech_mux2 U622 ( .A(iTSR[4]), .B(iTXFIFOQ[4]), .S(n679), .Z(n321) );
  notech_mux2 U623 ( .A(iTSR[3]), .B(iTXFIFOQ[3]), .S(n679), .Z(n320) );
  notech_mux2 U624 ( .A(iTSR[2]), .B(iTXFIFOQ[2]), .S(n679), .Z(n319) );
  notech_mux2 U625 ( .A(iTSR[1]), .B(iTXFIFOQ[1]), .S(n679), .Z(n318) );
  notech_mux2 U626 ( .A(iTSR[0]), .B(iTXFIFOQ[0]), .S(n679), .Z(n317) );
  notech_mux2 U627 ( .A(iSOUT), .B(iSINr), .S(n530), .Z(iSIN) );
  notech_nao3 U628 ( .C(n499), .A(n531), .B(iRXFIFOWrite), .Z(\U3/U1/Z_0 ) );
  notech_nao3 U629 ( .C(n496), .A(n500), .B(n438), .Z(n531) );
  notech_inv U630 ( .A(n498), .Z(n500) );
  notech_nor4 U631 ( .A(iFECounter[2]), .B(iFECounter[1]), .C(iFECounter[0]), 
        .D(n532), .Z(n498) );
  notech_or4 U632 ( .A(iFECounter[4]), .B(iFECounter[3]), .C(iFECounter[6]), 
        .D(iFECounter[5]), .Z(n532) );
  notech_ao3 U633 ( .A(n533), .B(n534), .C(iFERE), .Z(n496) );
  notech_inv U634 ( .A(iPERE), .Z(n534) );
  notech_inv U635 ( .A(iBIRE), .Z(n533) );
  notech_ao3 U636 ( .A(n535), .B(\UART_RXFF/n37 ), .C(iRXFIFOD[8]), .Z(n499)
         );
  notech_inv U638 ( .A(iRXFIFOD[10]), .Z(n535) );
  notech_and2 U639 ( .A(n422), .B(n537), .Z(N95) );
  notech_or2 U640 ( .A(iDIN[2]), .B(n538), .Z(n537) );
  notech_and2 U641 ( .A(n422), .B(n539), .Z(N94) );
  notech_or2 U642 ( .A(iDIN[1]), .B(n538), .Z(n539) );
  notech_xor2 U643 ( .A(iDIN[0]), .B(iIIR_6), .Z(n538) );
  notech_ao3 U644 ( .A(n528), .B(iA[1]), .C(iA[2]), .Z(n422) );
  notech_inv U645 ( .A(n540), .Z(N66) );
  notech_mux2 U646 ( .A(n435), .B(n450), .S(n449), .Z(n540) );
  notech_ao3 U647 ( .A(n541), .B(n542), .C(n448), .Z(n435) );
  notech_nand2 U648 ( .A(n543), .B(n544), .Z(n542) );
  notech_xor2 U649 ( .A(iFCR_RXTrigger[1]), .B(iFCR_RXTrigger[0]), .Z(n544) );
  notech_mux2 U650 ( .A(iRXFIFOUsage[5]), .B(iRXFIFOUsage[3]), .S(n545), .Z(
        n543) );
  notech_mux2 U651 ( .A(n546), .B(n547), .S(iFCR_RXTrigger[0]), .Z(n541) );
  notech_nao4 U652 ( .A(iRXFIFOUsage[4]), .B(n548), .C(n549), .D(n550), .Z(
        n547) );
  notech_and2 U653 ( .A(n551), .B(iRXFIFOUsage[3]), .Z(n549) );
  notech_ao4 U654 ( .A(iRXFIFOUsage[5]), .B(n548), .C(iRXFIFOUsage[4]), .D(
        iRXFIFOUsage[1]), .Z(n551) );
  notech_and2 U655 ( .A(iRXFIFOUsage[2]), .B(n545), .Z(n548) );
  notech_nand2 U656 ( .A(n438), .B(n550), .Z(n546) );
  notech_inv U657 ( .A(iFCR_RXTrigger[1]), .Z(n550) );
  notech_and2 U658 ( .A(WR), .B(CS), .Z(N48) );
  notech_or2 U659 ( .A(iMCR[4]), .B(iSOUT), .Z(N202) );
  notech_nand2 U660 ( .A(n530), .B(iMCR[0]), .Z(N201) );
  notech_nand2 U661 ( .A(n530), .B(iRTS), .Z(N200) );
  notech_nand2 U662 ( .A(n530), .B(iMCR[3]), .Z(N199) );
  notech_nand2 U663 ( .A(n530), .B(iMCR[2]), .Z(N198) );
  notech_inv U664 ( .A(n678), .Z(N197) );
  notech_and2 U665 ( .A(RD), .B(CS), .Z(n678) );
  notech_and2 U666 ( .A(n552), .B(State_snps_wire), .Z(N191) );
  notech_nand2 U667 ( .A(n448), .B(iIIR_6), .Z(n552) );
  notech_mux2 U668 ( .A(iRXFIFO64Full), .B(iRXFIFOUsage[4]), .S(n545), .Z(n448) );
  notech_or2 U669 ( .A(n553), .B(iFCR[1]), .Z(N190) );
  notech_and2 U670 ( .A(n673), .B(n449), .Z(n553) );
  notech_nor2 U671 ( .A(n680), .B(State_snps_wire), .Z(n673) );
  notech_or2 U673 ( .A(n554), .B(N182), .Z(N183) );
  notech_or2 U674 ( .A(n679), .B(n414), .Z(N182) );
  notech_nor2 U675 ( .A(n555), .B(State[1]), .Z(n679) );
  notech_or2 U676 ( .A(n554), .B(n556), .Z(N181) );
  notech_and2 U677 ( .A(iTXFinished), .B(n414), .Z(n556) );
  notech_and2 U678 ( .A(State[1]), .B(n555), .Z(n414) );
  notech_inv U679 ( .A(State[0]), .Z(n555) );
  notech_nor4 U680 ( .A(State[0]), .B(n557), .C(iTXFIFOEmpty), .D(State[1]), 
        .Z(n554) );
  notech_and2 U681 ( .A(n558), .B(iMCR[5]), .Z(n557) );
  notech_ao3 U682 ( .A(n521), .B(n528), .C(n559), .Z(N169) );
  notech_mux2 U683 ( .A(n560), .B(n520), .S(n449), .Z(n559) );
  notech_mux2 U684 ( .A(iTXFIFO64Full), .B(\iTXFIFOUsage[4] ), .S(n545), .Z(
        n560) );
  notech_and2 U685 ( .A(n442), .B(iWriteFE), .Z(n528) );
  notech_inv U686 ( .A(iA[0]), .Z(n442) );
  notech_and3 U687 ( .A(n512), .B(n516), .C(n508), .Z(n521) );
  notech_inv U688 ( .A(iA[1]), .Z(n508) );
  notech_inv U689 ( .A(iA[2]), .Z(n512) );
  notech_inv U690 ( .A(n561), .Z(N157) );
  notech_inv U691 ( .A(n562), .Z(N156) );
  notech_inv U692 ( .A(n563), .Z(N155) );
  notech_inv U693 ( .A(n558), .Z(N154) );
  notech_and2 U694 ( .A(iRXFIFOQ[8]), .B(n438), .Z(N146) );
  notech_nand3 U695 ( .A(n564), .B(n565), .C(n566), .Z(DOUT[7]) );
  notech_and3 U696 ( .A(n567), .B(n568), .C(n569), .Z(n566) );
  notech_ao4 U697 ( .A(n561), .B(n570), .C(n516), .D(n571), .Z(n569) );
  notech_inv U698 ( .A(iLCR[7]), .Z(n516) );
  notech_mux2 U699 ( .A(n572), .B(iDCDn), .S(n530), .Z(n561) );
  notech_nao3 U700 ( .C(n449), .A(iLSR_FIFOERR), .B(n573), .Z(n567) );
  notech_ao4 U701 ( .A(n574), .B(n575), .C(n576), .D(n577), .Z(n565) );
  notech_inv U702 ( .A(iDLL[7]), .Z(n576) );
  notech_inv U703 ( .A(iDLM[7]), .Z(n574) );
  notech_ao4 U704 ( .A(n578), .B(n579), .C(n580), .D(n581), .Z(n564) );
  notech_inv U705 ( .A(iSCR[7]), .Z(n580) );
  notech_inv U706 ( .A(iRXFIFOQ[7]), .Z(n579) );
  notech_nand3 U707 ( .A(n582), .B(n583), .C(n584), .Z(DOUT[6]) );
  notech_and3 U708 ( .A(n585), .B(n568), .C(n586), .Z(n584) );
  notech_ao4 U709 ( .A(n562), .B(n570), .C(n587), .D(n571), .Z(n586) );
  notech_inv U710 ( .A(iLCR[6]), .Z(n587) );
  notech_mux2 U711 ( .A(n588), .B(iRIn), .S(n530), .Z(n562) );
  notech_nao3 U712 ( .C(iTXRunning), .A(iTXFIFOEmpty), .B(n573), .Z(n585) );
  notech_ao4 U713 ( .A(n589), .B(n575), .C(n590), .D(n577), .Z(n583) );
  notech_inv U714 ( .A(iDLL[6]), .Z(n590) );
  notech_inv U715 ( .A(iDLM[6]), .Z(n589) );
  notech_ao4 U716 ( .A(n578), .B(n591), .C(n592), .D(n581), .Z(n582) );
  notech_inv U717 ( .A(iSCR[6]), .Z(n592) );
  notech_inv U718 ( .A(iRXFIFOQ[6]), .Z(n591) );
  notech_or4 U719 ( .A(n593), .B(n594), .C(n595), .D(n596), .Z(DOUT[5]) );
  notech_nao4 U720 ( .A(n597), .B(n571), .C(n434), .D(n598), .Z(n596) );
  notech_inv U721 ( .A(iMCR[5]), .Z(n434) );
  notech_inv U722 ( .A(iLCR[5]), .Z(n597) );
  notech_nand2 U723 ( .A(n599), .B(n600), .Z(n595) );
  notech_or2 U724 ( .A(n601), .B(n520), .Z(n600) );
  notech_inv U725 ( .A(iTXFIFOEmpty), .Z(n520) );
  notech_ao4 U726 ( .A(n545), .B(n568), .C(n563), .D(n570), .Z(n599) );
  notech_mux2 U727 ( .A(n602), .B(iDSRn), .S(n530), .Z(n563) );
  notech_or2 U728 ( .A(n603), .B(n449), .Z(n568) );
  notech_inv U729 ( .A(iIIR_6), .Z(n449) );
  notech_inv U730 ( .A(iFCR_5), .Z(n545) );
  notech_nao4 U731 ( .A(n604), .B(n581), .C(n578), .D(n605), .Z(n594) );
  notech_inv U732 ( .A(iRXFIFOQ[5]), .Z(n605) );
  notech_inv U733 ( .A(iSCR[5]), .Z(n604) );
  notech_nao4 U734 ( .A(n606), .B(n577), .C(n607), .D(n575), .Z(n593) );
  notech_inv U735 ( .A(iDLM[5]), .Z(n607) );
  notech_inv U736 ( .A(iDLL[5]), .Z(n606) );
  notech_or4 U737 ( .A(n608), .B(n609), .C(n610), .D(n611), .Z(DOUT[4]) );
  notech_nao4 U738 ( .A(n612), .B(n571), .C(n530), .D(n598), .Z(n611) );
  notech_inv U739 ( .A(iLCR[4]), .Z(n612) );
  notech_nao4 U740 ( .A(n507), .B(n601), .C(n558), .D(n570), .Z(n610) );
  notech_mux2 U741 ( .A(n437), .B(iCTSn), .S(n530), .Z(n558) );
  notech_inv U742 ( .A(iMCR[4]), .Z(n530) );
  notech_inv U743 ( .A(iRTS), .Z(n437) );
  notech_inv U744 ( .A(iLSR[4]), .Z(n507) );
  notech_nao4 U745 ( .A(n613), .B(n581), .C(n578), .D(n614), .Z(n609) );
  notech_inv U746 ( .A(iRXFIFOQ[4]), .Z(n614) );
  notech_inv U747 ( .A(n615), .Z(n578) );
  notech_inv U748 ( .A(iSCR[4]), .Z(n613) );
  notech_nao4 U749 ( .A(n616), .B(n577), .C(n617), .D(n575), .Z(n608) );
  notech_inv U750 ( .A(iDLM[4]), .Z(n617) );
  notech_inv U751 ( .A(iDLL[4]), .Z(n616) );
  notech_or4 U752 ( .A(n618), .B(n619), .C(n620), .D(n621), .Z(DOUT[3]) );
  notech_nand3 U753 ( .A(n622), .B(n623), .C(n624), .Z(n621) );
  notech_ao4 U754 ( .A(\UART_RX/n47 ), .B(n571), .C(n603), .D(n518), .Z(n624)
         );
  notech_inv U755 ( .A(iIIR[3]), .Z(n518) );
  notech_or2 U757 ( .A(n598), .B(n572), .Z(n623) );
  notech_inv U758 ( .A(iMCR[3]), .Z(n572) );
  notech_ao4 U759 ( .A(n426), .B(n570), .C(n478), .D(n601), .Z(n622) );
  notech_inv U760 ( .A(iLSR[3]), .Z(n478) );
  notech_inv U761 ( .A(iMSR[3]), .Z(n426) );
  notech_nao4 U762 ( .A(n626), .B(n627), .C(n628), .D(n581), .Z(n620) );
  notech_inv U763 ( .A(iSCR[3]), .Z(n628) );
  notech_inv U764 ( .A(iIER[3]), .Z(n626) );
  notech_nao4 U765 ( .A(n629), .B(n577), .C(n630), .D(n575), .Z(n619) );
  notech_inv U766 ( .A(iDLM[3]), .Z(n630) );
  notech_inv U767 ( .A(iDLL[3]), .Z(n629) );
  notech_and2 U768 ( .A(iRXFIFOQ[3]), .B(n615), .Z(n618) );
  notech_or4 U769 ( .A(n631), .B(n632), .C(n633), .D(n634), .Z(DOUT[2]) );
  notech_nand3 U770 ( .A(n635), .B(n636), .C(n637), .Z(n634) );
  notech_ao4 U771 ( .A(n638), .B(n571), .C(n603), .D(n517), .Z(n637) );
  notech_inv U772 ( .A(iIIR[2]), .Z(n517) );
  notech_inv U773 ( .A(iLCR[2]), .Z(n638) );
  notech_or2 U774 ( .A(n598), .B(n588), .Z(n636) );
  notech_inv U775 ( .A(iMCR[2]), .Z(n588) );
  notech_ao4 U776 ( .A(n431), .B(n570), .C(n476), .D(n601), .Z(n635) );
  notech_inv U777 ( .A(iLSR[2]), .Z(n476) );
  notech_inv U778 ( .A(iMSR[2]), .Z(n431) );
  notech_nao4 U779 ( .A(n639), .B(n627), .C(n640), .D(n581), .Z(n633) );
  notech_inv U780 ( .A(iSCR[2]), .Z(n640) );
  notech_inv U781 ( .A(iIER[2]), .Z(n639) );
  notech_nao4 U782 ( .A(n641), .B(n577), .C(n642), .D(n575), .Z(n632) );
  notech_inv U783 ( .A(iDLM[2]), .Z(n642) );
  notech_inv U784 ( .A(iDLL[2]), .Z(n641) );
  notech_and2 U785 ( .A(iRXFIFOQ[2]), .B(n615), .Z(n631) );
  notech_or4 U786 ( .A(n643), .B(n644), .C(n645), .D(n646), .Z(DOUT[1]) );
  notech_nand3 U787 ( .A(n647), .B(n648), .C(n649), .Z(n646) );
  notech_ao4 U788 ( .A(\UART_TX/n37 ), .B(n571), .C(n651), .D(n603), .Z(n649)
         );
  notech_inv U789 ( .A(iIIR[1]), .Z(n651) );
  notech_nand2 U791 ( .A(n652), .B(iMCR[1]), .Z(n648) );
  notech_ao4 U792 ( .A(n429), .B(n570), .C(n444), .D(n601), .Z(n647) );
  notech_inv U793 ( .A(iLSR[1]), .Z(n444) );
  notech_inv U794 ( .A(iMSR[1]), .Z(n429) );
  notech_nao4 U795 ( .A(n653), .B(n627), .C(n654), .D(n581), .Z(n645) );
  notech_inv U796 ( .A(iSCR[1]), .Z(n654) );
  notech_inv U797 ( .A(iIER[1]), .Z(n653) );
  notech_nao4 U798 ( .A(n655), .B(n577), .C(n656), .D(n575), .Z(n644) );
  notech_inv U799 ( .A(iDLM[1]), .Z(n656) );
  notech_inv U800 ( .A(iDLL[1]), .Z(n655) );
  notech_and2 U801 ( .A(iRXFIFOQ[1]), .B(n615), .Z(n643) );
  notech_or4 U802 ( .A(n657), .B(n658), .C(n659), .D(n660), .Z(DOUT[0]) );
  notech_nand3 U803 ( .A(n661), .B(n662), .C(n663), .Z(n660) );
  notech_ao4 U804 ( .A(\UART_TX/n24 ), .B(n571), .C(n603), .D(INT), .Z(n663)
         );
  notech_nao3 U805 ( .C(n665), .A(n666), .B(n667), .Z(n603) );
  notech_nand3 U806 ( .A(n666), .B(A[1]), .C(A[0]), .Z(n571) );
  notech_or2 U808 ( .A(n598), .B(n602), .Z(n662) );
  notech_inv U809 ( .A(iMCR[0]), .Z(n602) );
  notech_inv U810 ( .A(n652), .Z(n598) );
  notech_ao3 U811 ( .A(A[2]), .B(n665), .C(A[0]), .Z(n652) );
  notech_ao4 U812 ( .A(n441), .B(n570), .C(n450), .D(n601), .Z(n661) );
  notech_inv U813 ( .A(n573), .Z(n601) );
  notech_ao3 U814 ( .A(A[2]), .B(A[0]), .C(A[1]), .Z(n573) );
  notech_nor2 U815 ( .A(n438), .B(iRXFIFOWrite), .Z(n450) );
  notech_inv U816 ( .A(iRXFIFOEmpty), .Z(n438) );
  notech_nand3 U817 ( .A(n667), .B(A[1]), .C(A[2]), .Z(n570) );
  notech_inv U818 ( .A(iMSR[0]), .Z(n441) );
  notech_nao4 U819 ( .A(n668), .B(n627), .C(n669), .D(n581), .Z(n659) );
  notech_nao3 U820 ( .C(n667), .A(A[1]), .B(A[2]), .Z(n581) );
  notech_inv U821 ( .A(iSCR[0]), .Z(n669) );
  notech_or4 U822 ( .A(A[1]), .B(n667), .C(iLCR[7]), .D(A[2]), .Z(n627) );
  notech_inv U823 ( .A(iIER[0]), .Z(n668) );
  notech_nao4 U824 ( .A(n670), .B(n577), .C(n671), .D(n575), .Z(n658) );
  notech_nand2 U825 ( .A(n672), .B(A[0]), .Z(n575) );
  notech_inv U826 ( .A(iDLM[0]), .Z(n671) );
  notech_nand2 U827 ( .A(n672), .B(n667), .Z(n577) );
  notech_inv U828 ( .A(A[0]), .Z(n667) );
  notech_and3 U829 ( .A(n665), .B(n666), .C(iLCR[7]), .Z(n672) );
  notech_inv U830 ( .A(A[2]), .Z(n666) );
  notech_inv U831 ( .A(A[1]), .Z(n665) );
  notech_inv U832 ( .A(iDLL[0]), .Z(n670) );
  notech_and2 U833 ( .A(iRXFIFOQ[0]), .B(n615), .Z(n657) );
  notech_nor4 U834 ( .A(A[1]), .B(A[0]), .C(iLCR[7]), .D(A[2]), .Z(n615) );
  notech_inv \UART_ED_WRITE/U6  ( .A(\UART_ED_WRITE/iDd ), .Z(
        \UART_ED_WRITE/n1 ) );
  notech_nor2 \UART_ED_WRITE/U4  ( .A(\UART_ED_WRITE/n1 ), .B(N48), .Z(
        iWriteFE) );
  notech_reg \UART_ED_WRITE/iDd_reg  ( .D(N48), .CP(CLK), .CD(\UART_IS_DSR/n1 ), .Q(\UART_ED_WRITE/iDd ) );
  notech_inv \UART_ED_READ/U6  ( .A(\UART_ED_READ/iDd ), .Z(\UART_ED_READ/n1 )
         );
  notech_nor2 \UART_ED_READ/U4  ( .A(\UART_ED_READ/n1 ), .B(n678), .Z(iReadFE)
         );
  notech_reg \UART_ED_READ/iDd_reg  ( .D(n678), .CP(CLK), .CD(\UART_IS_DSR/n1 ), .Q(\UART_ED_READ/iDd ) );
  notech_inv \UART_IS_SIN/U3  ( .A(RST), .Z(\UART_IS_SIN/n1 ) );
  notech_reg \UART_IS_SIN/iD_reg[1]  ( .D(\UART_IS_SIN/iD[0] ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(iSINr) );
  notech_reg \UART_IS_SIN/iD_reg[0]  ( .D(SIN), .CP(CLK), .CD(\UART_IS_SIN/n1 ), .Q(\UART_IS_SIN/iD[0] ) );
  notech_inv \UART_IS_CTS/U3  ( .A(RST), .Z(\UART_IS_CTS/n1 ) );
  notech_reg \UART_IS_CTS/iD_reg[1]  ( .D(\UART_IS_CTS/iD[0] ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(iCTSNs) );
  notech_reg \UART_IS_CTS/iD_reg[0]  ( .D(CTSN), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_IS_CTS/iD[0] ) );
  notech_inv \UART_IS_DSR/U3  ( .A(RST), .Z(\UART_IS_DSR/n1 ) );
  notech_reg \UART_IS_DSR/iD_reg[1]  ( .D(\UART_IS_DSR/iD[0] ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(iDSRNs) );
  notech_reg \UART_IS_DSR/iD_reg[0]  ( .D(DSRN), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_IS_DSR/iD[0] ) );
  notech_inv \UART_IS_DCD/U3  ( .A(RST), .Z(\UART_IS_DCD/n1 ) );
  notech_reg \UART_IS_DCD/iD_reg[1]  ( .D(\UART_IS_DCD/iD[0] ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(iDCDNs) );
  notech_reg \UART_IS_DCD/iD_reg[0]  ( .D(DCDN), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_IS_DCD/iD[0] ) );
  notech_inv \UART_IS_RI/U3  ( .A(RST), .Z(\UART_IS_RI/n1 ) );
  notech_reg \UART_IS_RI/iD_reg[1]  ( .D(\UART_IS_RI/iD[0] ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(iRINs) );
  notech_reg \UART_IS_RI/iD_reg[0]  ( .D(RIN), .CP(CLK), .CD(\UART_IS_RI/n1 ), 
        .Q(\UART_IS_RI/iD[0] ) );
  notech_mux2 \UART_IF_CTS/U13  ( .A(\UART_IF_CTS/iCount[1] ), .B(iCTSn), .S(
        \UART_IF_CTS/iCount[0] ), .Z(\UART_IF_CTS/n16 ) );
  notech_and3 \UART_IF_CTS/U12  ( .A(\UART_IF_CTS/iCount[0] ), .B(iCTSNs), .C(
        iBaudtick2x), .Z(\UART_IF_CTS/n5 ) );
  notech_xor2 \UART_IF_CTS/U10  ( .A(\UART_IF_CTS/iCount[0] ), .B(iCTSNs), .Z(
        \UART_IF_CTS/n7 ) );
  notech_or2 \UART_IF_CTS/U9  ( .A(\UART_IF_RI/n3 ), .B(\UART_IF_CTS/n7 ), .Z(
        \UART_IF_CTS/n6 ) );
  notech_mux2 \UART_IF_CTS/U8  ( .A(\UART_IF_CTS/n5 ), .B(\UART_IF_CTS/n6 ), 
        .S(\UART_IF_CTS/iCount[1] ), .Z(\UART_IF_CTS/n17 ) );
  notech_xor2 \UART_IF_CTS/U7  ( .A(\UART_IF_CTS/iCount[1] ), .B(iCTSNs), .Z(
        \UART_IF_CTS/n4 ) );
  notech_nor2 \UART_IF_CTS/U6  ( .A(\UART_IF_CTS/iCount[0] ), .B(
        \UART_IF_CTS/n4 ), .Z(\UART_IF_CTS/n2 ) );
  notech_nor2 \UART_IF_CTS/U5  ( .A(\UART_IF_CTS/n2 ), .B(\UART_IF_RI/n3 ), 
        .Z(\UART_IF_CTS/n1 ) );
  notech_xor2 \UART_IF_CTS/U4  ( .A(\UART_IF_CTS/iCount[0] ), .B(
        \UART_IF_CTS/n1 ), .Z(\UART_IF_CTS/n18 ) );
  notech_inv \UART_IF_CTS/U3  ( .A(RST), .Z(\UART_IF_CTS/n8 ) );
  notech_reg \UART_IF_CTS/Q_reg  ( .D(\UART_IF_CTS/n16 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(iCTSn) );
  notech_reg \UART_IF_CTS/iCount_reg[1]  ( .D(\UART_IF_CTS/n17 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_IF_CTS/iCount[1] ) );
  notech_reg \UART_IF_CTS/iCount_reg[0]  ( .D(\UART_IF_CTS/n18 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_IF_CTS/iCount[0] ) );
  notech_mux2 \UART_IF_DSR/U13  ( .A(\UART_IF_DSR/iCount[1] ), .B(iDSRn), .S(
        \UART_IF_DSR/iCount[0] ), .Z(\UART_IF_DSR/n11 ) );
  notech_and3 \UART_IF_DSR/U12  ( .A(\UART_IF_DSR/iCount[0] ), .B(iDSRNs), .C(
        iBaudtick2x), .Z(\UART_IF_DSR/n5 ) );
  notech_xor2 \UART_IF_DSR/U10  ( .A(\UART_IF_DSR/iCount[0] ), .B(iDSRNs), .Z(
        \UART_IF_DSR/n7 ) );
  notech_or2 \UART_IF_DSR/U9  ( .A(\UART_IF_RI/n3 ), .B(\UART_IF_DSR/n7 ), .Z(
        \UART_IF_DSR/n6 ) );
  notech_mux2 \UART_IF_DSR/U8  ( .A(\UART_IF_DSR/n5 ), .B(\UART_IF_DSR/n6 ), 
        .S(\UART_IF_DSR/iCount[1] ), .Z(\UART_IF_DSR/n10 ) );
  notech_xor2 \UART_IF_DSR/U7  ( .A(\UART_IF_DSR/iCount[1] ), .B(iDSRNs), .Z(
        \UART_IF_DSR/n4 ) );
  notech_nor2 \UART_IF_DSR/U6  ( .A(\UART_IF_DSR/iCount[0] ), .B(
        \UART_IF_DSR/n4 ), .Z(\UART_IF_DSR/n2 ) );
  notech_nor2 \UART_IF_DSR/U5  ( .A(\UART_IF_DSR/n2 ), .B(\UART_IF_RI/n3 ), 
        .Z(\UART_IF_DSR/n1 ) );
  notech_xor2 \UART_IF_DSR/U4  ( .A(\UART_IF_DSR/iCount[0] ), .B(
        \UART_IF_DSR/n1 ), .Z(\UART_IF_DSR/n9 ) );
  notech_inv \UART_IF_DSR/U3  ( .A(RST), .Z(\UART_IF_DSR/n8 ) );
  notech_reg \UART_IF_DSR/Q_reg  ( .D(\UART_IF_DSR/n11 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(iDSRn) );
  notech_reg \UART_IF_DSR/iCount_reg[1]  ( .D(\UART_IF_DSR/n10 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_IF_DSR/iCount[1] ) );
  notech_reg \UART_IF_DSR/iCount_reg[0]  ( .D(\UART_IF_DSR/n9 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_IF_DSR/iCount[0] ) );
  notech_mux2 \UART_IF_DCD/U13  ( .A(\UART_IF_DCD/iCount[1] ), .B(iDCDn), .S(
        \UART_IF_DCD/iCount[0] ), .Z(\UART_IF_DCD/n11 ) );
  notech_and3 \UART_IF_DCD/U12  ( .A(\UART_IF_DCD/iCount[0] ), .B(iDCDNs), .C(
        iBaudtick2x), .Z(\UART_IF_DCD/n5 ) );
  notech_xor2 \UART_IF_DCD/U10  ( .A(\UART_IF_DCD/iCount[0] ), .B(iDCDNs), .Z(
        \UART_IF_DCD/n7 ) );
  notech_or2 \UART_IF_DCD/U9  ( .A(\UART_IF_RI/n3 ), .B(\UART_IF_DCD/n7 ), .Z(
        \UART_IF_DCD/n6 ) );
  notech_mux2 \UART_IF_DCD/U8  ( .A(\UART_IF_DCD/n5 ), .B(\UART_IF_DCD/n6 ), 
        .S(\UART_IF_DCD/iCount[1] ), .Z(\UART_IF_DCD/n10 ) );
  notech_xor2 \UART_IF_DCD/U7  ( .A(\UART_IF_DCD/iCount[1] ), .B(iDCDNs), .Z(
        \UART_IF_DCD/n4 ) );
  notech_nor2 \UART_IF_DCD/U6  ( .A(\UART_IF_DCD/iCount[0] ), .B(
        \UART_IF_DCD/n4 ), .Z(\UART_IF_DCD/n2 ) );
  notech_nor2 \UART_IF_DCD/U5  ( .A(\UART_IF_DCD/n2 ), .B(\UART_IF_RI/n3 ), 
        .Z(\UART_IF_DCD/n1 ) );
  notech_xor2 \UART_IF_DCD/U4  ( .A(\UART_IF_DCD/iCount[0] ), .B(
        \UART_IF_DCD/n1 ), .Z(\UART_IF_DCD/n9 ) );
  notech_reg \UART_IF_DCD/Q_reg  ( .D(\UART_IF_DCD/n11 ), .CP(CLK), .CD(n419), 
        .Q(iDCDn) );
  notech_reg \UART_IF_DCD/iCount_reg[1]  ( .D(\UART_IF_DCD/n10 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_IF_DCD/iCount[1] ) );
  notech_reg \UART_IF_DCD/iCount_reg[0]  ( .D(\UART_IF_DCD/n9 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_IF_DCD/iCount[0] ) );
  notech_mux2 \UART_IF_RI/U13  ( .A(\UART_IF_RI/iCount[1] ), .B(iRIn), .S(
        \UART_IF_RI/iCount[0] ), .Z(\UART_IF_RI/n11 ) );
  notech_and3 \UART_IF_RI/U12  ( .A(\UART_IF_RI/iCount[0] ), .B(iRINs), .C(
        iBaudtick2x), .Z(\UART_IF_RI/n5 ) );
  notech_inv \UART_IF_RI/U11  ( .A(iBaudtick2x), .Z(\UART_IF_RI/n3 ) );
  notech_xor2 \UART_IF_RI/U10  ( .A(\UART_IF_RI/iCount[0] ), .B(iRINs), .Z(
        \UART_IF_RI/n7 ) );
  notech_or2 \UART_IF_RI/U9  ( .A(\UART_IF_RI/n3 ), .B(\UART_IF_RI/n7 ), .Z(
        \UART_IF_RI/n6 ) );
  notech_mux2 \UART_IF_RI/U8  ( .A(\UART_IF_RI/n5 ), .B(\UART_IF_RI/n6 ), .S(
        \UART_IF_RI/iCount[1] ), .Z(\UART_IF_RI/n10 ) );
  notech_xor2 \UART_IF_RI/U7  ( .A(\UART_IF_RI/iCount[1] ), .B(iRINs), .Z(
        \UART_IF_RI/n4 ) );
  notech_nor2 \UART_IF_RI/U6  ( .A(\UART_IF_RI/iCount[0] ), .B(\UART_IF_RI/n4 ), .Z(\UART_IF_RI/n2 ) );
  notech_nor2 \UART_IF_RI/U5  ( .A(\UART_IF_RI/n2 ), .B(\UART_IF_RI/n3 ), .Z(
        \UART_IF_RI/n1 ) );
  notech_xor2 \UART_IF_RI/U4  ( .A(\UART_IF_RI/iCount[0] ), .B(\UART_IF_RI/n1 ), .Z(\UART_IF_RI/n9 ) );
  notech_reg \UART_IF_RI/Q_reg  ( .D(\UART_IF_RI/n11 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(iRIn) );
  notech_reg \UART_IF_RI/iCount_reg[1]  ( .D(\UART_IF_RI/n10 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_IF_RI/iCount[1] ) );
  notech_reg \UART_IF_RI/iCount_reg[0]  ( .D(\UART_IF_RI/n9 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_IF_RI/iCount[0] ) );
  notech_nand2 \UART_IIC/U18  ( .A(iTHRInterrupt), .B(iIER[1]), .Z(
        \UART_IIC/n5 ) );
  notech_and2 \UART_IIC/U16  ( .A(iMSR[0]), .B(n434), .Z(\UART_IIC/n9 ) );
  notech_or4 \UART_IIC/U15  ( .A(iMSR[1]), .B(\UART_IIC/n9 ), .C(iMSR[3]), .D(
        iMSR[2]), .Z(\UART_IIC/n8 ) );
  notech_nand2 \UART_IIC/U14  ( .A(iIER[3]), .B(\UART_IIC/n8 ), .Z(
        \UART_IIC/n6 ) );
  notech_or4 \UART_IIC/U13  ( .A(iLSR[2]), .B(iLSR[1]), .C(iLSR[4]), .D(
        iLSR[3]), .Z(\UART_IIC/n7 ) );
  notech_and2 \UART_IIC/U12  ( .A(iIER[2]), .B(\UART_IIC/n7 ), .Z(
        \UART_IIC/n1 ) );
  notech_nand2 \UART_IIC/U11  ( .A(iIER[0]), .B(iCharTimeout), .Z(
        \UART_IIC/n2 ) );
  notech_nand2 \UART_IIC/U10  ( .A(N66), .B(iIER[0]), .Z(\UART_IIC/n4 ) );
  notech_nao3 \UART_IIC/U9  ( .C(\UART_IIC/n1 ), .A(\UART_IIC/n2 ), .B(
        \UART_IIC/n4 ), .Z(\UART_IIC/N21 ) );
  notech_ao3 \UART_IIC/U8  ( .A(\UART_IIC/n5 ), .B(\UART_IIC/n6 ), .C(
        \UART_IIC/N21 ), .Z(\UART_IIC/N19 ) );
  notech_ao3 \UART_IIC/U7  ( .A(\UART_IIC/n4 ), .B(\UART_IIC/n2 ), .C(
        \UART_IIC/n5 ), .Z(\UART_IIC/n3 ) );
  notech_or2 \UART_IIC/U6  ( .A(\UART_IIC/n3 ), .B(\UART_IIC/n1 ), .Z(
        \UART_IIC/N20 ) );
  notech_nor2 \UART_IIC/U5  ( .A(\UART_IIC/n1 ), .B(\UART_IIC/n2 ), .Z(
        \UART_IIC/N22 ) );
  notech_inv \UART_IIC/U3  ( .A(\UART_IIC/IIR[0] ), .Z(INT) );
  notech_reg_set \UART_IIC/iIIR_reg[0]  ( .D(\UART_IIC/N19 ), .CP(CLK), .SD(
        \UART_IS_DSR/n1 ), .Q(\UART_IIC/IIR[0] ) );
  notech_reg \UART_IIC/iIIR_reg[1]  ( .D(\UART_IIC/N20 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(iIIR[1]) );
  notech_reg \UART_IIC/iIIR_reg[2]  ( .D(\UART_IIC/N21 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(iIIR[2]) );
  notech_reg \UART_IIC/iIIR_reg[3]  ( .D(\UART_IIC/N22 ), .CP(CLK), .CD(n420), 
        .Q(iIIR[3]) );
  notech_inv \UART_IIC_THRE_ED/U6  ( .A(\UART_IIC_THRE_ED/iDd ), .Z(
        \UART_IIC_THRE_ED/n1 ) );
  notech_and2 \UART_IIC_THRE_ED/U5  ( .A(iTXFIFOEmpty), .B(
        \UART_IIC_THRE_ED/n1 ), .Z(iLSR_THRERE) );
  notech_reg \UART_IIC_THRE_ED/iDd_reg  ( .D(iTXFIFOEmpty), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(\UART_IIC_THRE_ED/iDd ) );
  notech_inv \UART_PEDET/U6  ( .A(\UART_PEDET/iDd ), .Z(\UART_PEDET/n1 ) );
  notech_and2 \UART_PEDET/U5  ( .A(N146), .B(\UART_PEDET/n1 ), .Z(iPERE) );
  notech_reg \UART_PEDET/iDd_reg  ( .D(N146), .CP(CLK), .CD(\UART_IS_CTS/n1 ), 
        .Q(\UART_PEDET/iDd ) );
  notech_inv \UART_FEDET/U6  ( .A(\UART_FEDET/iDd ), .Z(\UART_FEDET/n1 ) );
  notech_and2 \UART_FEDET/U5  ( .A(n675), .B(\UART_FEDET/n1 ), .Z(iFERE) );
  notech_reg \UART_FEDET/iDd_reg  ( .D(n675), .CP(CLK), .CD(\UART_IS_RI/n1 ), 
        .Q(\UART_FEDET/iDd ) );
  notech_inv \UART_BIDET/U6  ( .A(\UART_BIDET/iDd ), .Z(\UART_BIDET/n1 ) );
  notech_and2 \UART_BIDET/U5  ( .A(n674), .B(\UART_BIDET/n1 ), .Z(iBIRE) );
  notech_reg \UART_BIDET/iDd_reg  ( .D(n674), .CP(CLK), .CD(\UART_IF_CTS/n8 ), 
        .Q(\UART_BIDET/iDd ) );
  notech_inv \UART_ED_CTS/U6  ( .A(\UART_ED_CTS/iDd ), .Z(\UART_ED_CTS/n1 ) );
  notech_nor2 \UART_ED_CTS/U4  ( .A(\UART_ED_CTS/n1 ), .B(N154), .Z(iCTSnFE)
         );
  notech_reg \UART_ED_CTS/iDd_reg  ( .D(N154), .CP(CLK), .CD(\UART_IS_RI/n1 ), 
        .Q(\UART_ED_CTS/iDd ) );
  notech_inv \UART_ED_DSR/U6  ( .A(\UART_ED_DSR/iDd ), .Z(\UART_ED_DSR/n1 ) );
  notech_nor2 \UART_ED_DSR/U4  ( .A(\UART_ED_DSR/n1 ), .B(N155), .Z(iDSRnFE)
         );
  notech_reg \UART_ED_DSR/iDd_reg  ( .D(N155), .CP(CLK), .CD(\UART_IS_SIN/n1 ), 
        .Q(\UART_ED_DSR/iDd ) );
  notech_inv \UART_ED_RI/U6  ( .A(\UART_ED_RI/iDd ), .Z(\UART_ED_RI/n1 ) );
  notech_nor2 \UART_ED_RI/U4  ( .A(\UART_ED_RI/n1 ), .B(N156), .Z(iRInFE) );
  notech_reg \UART_ED_RI/iDd_reg  ( .D(N156), .CP(CLK), .CD(\UART_IF_DSR/n8 ), 
        .Q(\UART_ED_RI/iDd ) );
  notech_inv \UART_ED_DCD/U6  ( .A(\UART_ED_DCD/iDd ), .Z(\UART_ED_DCD/n1 ) );
  notech_nor2 \UART_ED_DCD/U4  ( .A(\UART_ED_DCD/n1 ), .B(N157), .Z(iDCDnFE)
         );
  notech_reg \UART_ED_DCD/iDd_reg  ( .D(N157), .CP(CLK), .CD(\UART_IS_CTS/n1 ), 
        .Q(\UART_ED_DCD/iDd ) );
  notech_xor2 \UART_BG16/U76  ( .A(\UART_BG16/iCounter[4] ), .B(iDLL[4]), .Z(
        \UART_BG16/n69 ) );
  notech_xor2 \UART_BG16/U75  ( .A(\UART_BG16/iCounter[5] ), .B(iDLL[5]), .Z(
        \UART_BG16/n70 ) );
  notech_xor2 \UART_BG16/U74  ( .A(\UART_BG16/iCounter[9] ), .B(iDLM[1]), .Z(
        \UART_BG16/n71 ) );
  notech_xor2 \UART_BG16/U73  ( .A(\UART_BG16/iCounter[10] ), .B(iDLM[2]), .Z(
        \UART_BG16/n72 ) );
  notech_or4 \UART_BG16/U72  ( .A(\UART_BG16/n69 ), .B(\UART_BG16/n70 ), .C(
        \UART_BG16/n71 ), .D(\UART_BG16/n72 ), .Z(\UART_BG16/n37 ) );
  notech_xor2 \UART_BG16/U71  ( .A(\UART_BG16/iCounter[1] ), .B(iDLL[1]), .Z(
        \UART_BG16/n65 ) );
  notech_xor2 \UART_BG16/U70  ( .A(\UART_BG16/iCounter[2] ), .B(iDLL[2]), .Z(
        \UART_BG16/n66 ) );
  notech_xor2 \UART_BG16/U69  ( .A(\UART_BG16/iCounter[6] ), .B(iDLL[6]), .Z(
        \UART_BG16/n67 ) );
  notech_xor2 \UART_BG16/U68  ( .A(\UART_BG16/iCounter[0] ), .B(iDLL[0]), .Z(
        \UART_BG16/n68 ) );
  notech_or4 \UART_BG16/U67  ( .A(\UART_BG16/n65 ), .B(\UART_BG16/n66 ), .C(
        \UART_BG16/n67 ), .D(\UART_BG16/n68 ), .Z(\UART_BG16/n38 ) );
  notech_xor2 \UART_BG16/U66  ( .A(\UART_BG16/iCounter[3] ), .B(iDLL[3]), .Z(
        \UART_BG16/n61 ) );
  notech_xor2 \UART_BG16/U65  ( .A(\UART_BG16/iCounter[15] ), .B(iDLM[7]), .Z(
        \UART_BG16/n62 ) );
  notech_xor2 \UART_BG16/U64  ( .A(\UART_BG16/iCounter[11] ), .B(iDLM[3]), .Z(
        \UART_BG16/n63 ) );
  notech_xor2 \UART_BG16/U63  ( .A(\UART_BG16/iCounter[7] ), .B(iDLL[7]), .Z(
        \UART_BG16/n64 ) );
  notech_or4 \UART_BG16/U62  ( .A(\UART_BG16/n61 ), .B(\UART_BG16/n62 ), .C(
        \UART_BG16/n63 ), .D(\UART_BG16/n64 ), .Z(\UART_BG16/n39 ) );
  notech_xor2 \UART_BG16/U61  ( .A(\UART_BG16/iCounter[14] ), .B(iDLM[6]), .Z(
        \UART_BG16/n57 ) );
  notech_xor2 \UART_BG16/U60  ( .A(\UART_BG16/iCounter[8] ), .B(iDLM[0]), .Z(
        \UART_BG16/n58 ) );
  notech_xor2 \UART_BG16/U59  ( .A(\UART_BG16/iCounter[12] ), .B(iDLM[4]), .Z(
        \UART_BG16/n59 ) );
  notech_xor2 \UART_BG16/U58  ( .A(\UART_BG16/iCounter[13] ), .B(iDLM[5]), .Z(
        \UART_BG16/n60 ) );
  notech_or4 \UART_BG16/U57  ( .A(\UART_BG16/n57 ), .B(\UART_BG16/n58 ), .C(
        \UART_BG16/n59 ), .D(\UART_BG16/n60 ), .Z(\UART_BG16/n56 ) );
  notech_nor4 \UART_BG16/U56  ( .A(\UART_BG16/n37 ), .B(\UART_BG16/n38 ), .C(
        \UART_BG16/n39 ), .D(\UART_BG16/n56 ), .Z(\UART_BG16/N40 ) );
  notech_inv \UART_BG16/U55  ( .A(\UART_BG16/N40 ), .Z(\UART_BG16/n35 ) );
  notech_inv \UART_BG16/U53  ( .A(\UART_BG16/N22 ), .Z(\UART_BG16/n32 ) );
  notech_inv \UART_BG16/U52  ( .A(\UART_BG16/iCounter[15] ), .Z(
        \UART_BG16/n33 ) );
  notech_nao4 \UART_BG16/U48  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n32 ), .C(
        \UART_BG16/n33 ), .D(n682), .Z(\UART_BG16/n40 ) );
  notech_inv \UART_BG16/U47  ( .A(\UART_BG16/N21 ), .Z(\UART_BG16/n30 ) );
  notech_inv \UART_BG16/U46  ( .A(\UART_BG16/iCounter[14] ), .Z(
        \UART_BG16/n31 ) );
  notech_nao4 \UART_BG16/U45  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n30 ), .C(
        \UART_BG16/n31 ), .D(n682), .Z(\UART_BG16/n41 ) );
  notech_inv \UART_BG16/U44  ( .A(\UART_BG16/N20 ), .Z(\UART_BG16/n28 ) );
  notech_inv \UART_BG16/U43  ( .A(\UART_BG16/iCounter[13] ), .Z(
        \UART_BG16/n29 ) );
  notech_nao4 \UART_BG16/U42  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n28 ), .C(
        \UART_BG16/n29 ), .D(n682), .Z(\UART_BG16/n42 ) );
  notech_inv \UART_BG16/U41  ( .A(\UART_BG16/N19 ), .Z(\UART_BG16/n26 ) );
  notech_inv \UART_BG16/U40  ( .A(\UART_BG16/iCounter[12] ), .Z(
        \UART_BG16/n27 ) );
  notech_nao4 \UART_BG16/U39  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n26 ), .C(
        \UART_BG16/n27 ), .D(n682), .Z(\UART_BG16/n43 ) );
  notech_inv \UART_BG16/U38  ( .A(\UART_BG16/N18 ), .Z(\UART_BG16/n24 ) );
  notech_inv \UART_BG16/U37  ( .A(\UART_BG16/iCounter[11] ), .Z(
        \UART_BG16/n25 ) );
  notech_nao4 \UART_BG16/U36  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n24 ), .C(
        \UART_BG16/n25 ), .D(n682), .Z(\UART_BG16/n44 ) );
  notech_inv \UART_BG16/U35  ( .A(\UART_BG16/N17 ), .Z(\UART_BG16/n22 ) );
  notech_inv \UART_BG16/U34  ( .A(\UART_BG16/iCounter[10] ), .Z(
        \UART_BG16/n23 ) );
  notech_nao4 \UART_BG16/U33  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n22 ), .C(
        \UART_BG16/n23 ), .D(n682), .Z(\UART_BG16/n45 ) );
  notech_inv \UART_BG16/U32  ( .A(\UART_BG16/N16 ), .Z(\UART_BG16/n20 ) );
  notech_inv \UART_BG16/U31  ( .A(\UART_BG16/iCounter[9] ), .Z(\UART_BG16/n21 ) );
  notech_nao4 \UART_BG16/U30  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n20 ), .C(
        \UART_BG16/n21 ), .D(n682), .Z(\UART_BG16/n46 ) );
  notech_inv \UART_BG16/U29  ( .A(\UART_BG16/N15 ), .Z(\UART_BG16/n18 ) );
  notech_inv \UART_BG16/U28  ( .A(\UART_BG16/iCounter[8] ), .Z(\UART_BG16/n19 ) );
  notech_nao4 \UART_BG16/U27  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n18 ), .C(
        \UART_BG16/n19 ), .D(n682), .Z(\UART_BG16/n47 ) );
  notech_inv \UART_BG16/U26  ( .A(\UART_BG16/N14 ), .Z(\UART_BG16/n16 ) );
  notech_inv \UART_BG16/U25  ( .A(\UART_BG16/iCounter[7] ), .Z(\UART_BG16/n17 ) );
  notech_nao4 \UART_BG16/U24  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n16 ), .C(
        \UART_BG16/n17 ), .D(n682), .Z(\UART_BG16/n48 ) );
  notech_inv \UART_BG16/U23  ( .A(\UART_BG16/N13 ), .Z(\UART_BG16/n14 ) );
  notech_inv \UART_BG16/U22  ( .A(\UART_BG16/iCounter[6] ), .Z(\UART_BG16/n15 ) );
  notech_nao4 \UART_BG16/U21  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n14 ), .C(
        \UART_BG16/n15 ), .D(n682), .Z(\UART_BG16/n49 ) );
  notech_inv \UART_BG16/U20  ( .A(\UART_BG16/N12 ), .Z(\UART_BG16/n12 ) );
  notech_inv \UART_BG16/U19  ( .A(\UART_BG16/iCounter[5] ), .Z(\UART_BG16/n13 ) );
  notech_nao4 \UART_BG16/U18  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n12 ), .C(
        \UART_BG16/n13 ), .D(n682), .Z(\UART_BG16/n50 ) );
  notech_inv \UART_BG16/U17  ( .A(\UART_BG16/N11 ), .Z(\UART_BG16/n10 ) );
  notech_inv \UART_BG16/U16  ( .A(\UART_BG16/iCounter[4] ), .Z(\UART_BG16/n11 ) );
  notech_nao4 \UART_BG16/U15  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n10 ), .C(
        \UART_BG16/n11 ), .D(n682), .Z(\UART_BG16/n51 ) );
  notech_inv \UART_BG16/U14  ( .A(\UART_BG16/N10 ), .Z(\UART_BG16/n8 ) );
  notech_inv \UART_BG16/U13  ( .A(\UART_BG16/iCounter[3] ), .Z(\UART_BG16/n9 )
         );
  notech_nao4 \UART_BG16/U12  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n8 ), .C(
        \UART_BG16/n9 ), .D(n682), .Z(\UART_BG16/n52 ) );
  notech_inv \UART_BG16/U11  ( .A(\UART_BG16/N9 ), .Z(\UART_BG16/n6 ) );
  notech_inv \UART_BG16/U10  ( .A(\UART_BG16/iCounter[2] ), .Z(\UART_BG16/n7 )
         );
  notech_nao4 \UART_BG16/U9  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n6 ), .C(
        \UART_BG16/n7 ), .D(n682), .Z(\UART_BG16/n53 ) );
  notech_inv \UART_BG16/U8  ( .A(\UART_BG16/N8 ), .Z(\UART_BG16/n4 ) );
  notech_inv \UART_BG16/U7  ( .A(\UART_BG16/iCounter[1] ), .Z(\UART_BG16/n5 )
         );
  notech_nao4 \UART_BG16/U6  ( .A(\UART_BG16/n2 ), .B(\UART_BG16/n4 ), .C(
        \UART_BG16/n5 ), .D(n682), .Z(\UART_BG16/n54 ) );
  notech_mux2 \UART_BG16/U5  ( .A(\UART_BG16/n2 ), .B(n682), .S(
        \UART_BG16/iCounter[0] ), .Z(\UART_BG16/n1 ) );
  notech_inv \UART_BG16/U4  ( .A(\UART_BG16/n1 ), .Z(\UART_BG16/n55 ) );
  notech_reg \UART_BG16/iCounter_reg[15]  ( .D(\UART_BG16/n40 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_BG16/iCounter[15] ) );
  notech_reg \UART_BG16/iCounter_reg[14]  ( .D(\UART_BG16/n41 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_BG16/iCounter[14] ) );
  notech_reg \UART_BG16/iCounter_reg[13]  ( .D(\UART_BG16/n42 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_BG16/iCounter[13] ) );
  notech_reg \UART_BG16/iCounter_reg[12]  ( .D(\UART_BG16/n43 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_BG16/iCounter[12] ) );
  notech_reg \UART_BG16/iCounter_reg[11]  ( .D(\UART_BG16/n44 ), .CP(CLK), 
        .CD(\UART_IS_SIN/n1 ), .Q(\UART_BG16/iCounter[11] ) );
  notech_reg \UART_BG16/iCounter_reg[10]  ( .D(\UART_BG16/n45 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_BG16/iCounter[10] ) );
  notech_reg \UART_BG16/iCounter_reg[9]  ( .D(\UART_BG16/n46 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_BG16/iCounter[9] ) );
  notech_reg \UART_BG16/iCounter_reg[8]  ( .D(\UART_BG16/n47 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_BG16/iCounter[8] ) );
  notech_reg \UART_BG16/iCounter_reg[7]  ( .D(\UART_BG16/n48 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(\UART_BG16/iCounter[7] ) );
  notech_reg \UART_BG16/iCounter_reg[6]  ( .D(\UART_BG16/n49 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(\UART_BG16/iCounter[6] ) );
  notech_reg \UART_BG16/iCounter_reg[5]  ( .D(\UART_BG16/n50 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(\UART_BG16/iCounter[5] ) );
  notech_reg \UART_BG16/iCounter_reg[4]  ( .D(\UART_BG16/n51 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(\UART_BG16/iCounter[4] ) );
  notech_reg \UART_BG16/iCounter_reg[3]  ( .D(\UART_BG16/n52 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(\UART_BG16/iCounter[3] ) );
  notech_reg \UART_BG16/iCounter_reg[2]  ( .D(\UART_BG16/n53 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_BG16/iCounter[2] ) );
  notech_reg \UART_BG16/iCounter_reg[1]  ( .D(\UART_BG16/n54 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_BG16/iCounter[1] ) );
  notech_reg \UART_BG16/BAUDTICK_reg  ( .D(\UART_BG16/N40 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(iBaudtick16x) );
  notech_reg \UART_BG16/iCounter_reg[0]  ( .D(\UART_BG16/n55 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_BG16/iCounter[0] ) );
  notech_xor2 \UART_BG16/add_54/U1  ( .A(\UART_BG16/add_54/carry [15]), .B(
        \UART_BG16/iCounter[15] ), .Z(\UART_BG16/N22 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_1  ( .A(\UART_BG16/iCounter[1] ), .B(
        \UART_BG16/iCounter[0] ), .CO(\UART_BG16/add_54/carry [2]), .Z(
        \UART_BG16/N8 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_2  ( .A(\UART_BG16/iCounter[2] ), .B(
        \UART_BG16/add_54/carry [2]), .CO(\UART_BG16/add_54/carry [3]), .Z(
        \UART_BG16/N9 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_3  ( .A(\UART_BG16/iCounter[3] ), .B(
        \UART_BG16/add_54/carry [3]), .CO(\UART_BG16/add_54/carry [4]), .Z(
        \UART_BG16/N10 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_4  ( .A(\UART_BG16/iCounter[4] ), .B(
        \UART_BG16/add_54/carry [4]), .CO(\UART_BG16/add_54/carry [5]), .Z(
        \UART_BG16/N11 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_5  ( .A(\UART_BG16/iCounter[5] ), .B(
        \UART_BG16/add_54/carry [5]), .CO(\UART_BG16/add_54/carry [6]), .Z(
        \UART_BG16/N12 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_6  ( .A(\UART_BG16/iCounter[6] ), .B(
        \UART_BG16/add_54/carry [6]), .CO(\UART_BG16/add_54/carry [7]), .Z(
        \UART_BG16/N13 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_7  ( .A(\UART_BG16/iCounter[7] ), .B(
        \UART_BG16/add_54/carry [7]), .CO(\UART_BG16/add_54/carry [8]), .Z(
        \UART_BG16/N14 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_8  ( .A(\UART_BG16/iCounter[8] ), .B(
        \UART_BG16/add_54/carry [8]), .CO(\UART_BG16/add_54/carry [9]), .Z(
        \UART_BG16/N15 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_9  ( .A(\UART_BG16/iCounter[9] ), .B(
        \UART_BG16/add_54/carry [9]), .CO(\UART_BG16/add_54/carry [10]), .Z(
        \UART_BG16/N16 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_10  ( .A(\UART_BG16/iCounter[10] ), .B(
        \UART_BG16/add_54/carry [10]), .CO(\UART_BG16/add_54/carry [11]), .Z(
        \UART_BG16/N17 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_11  ( .A(\UART_BG16/iCounter[11] ), .B(
        \UART_BG16/add_54/carry [11]), .CO(\UART_BG16/add_54/carry [12]), .Z(
        \UART_BG16/N18 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_12  ( .A(\UART_BG16/iCounter[12] ), .B(
        \UART_BG16/add_54/carry [12]), .CO(\UART_BG16/add_54/carry [13]), .Z(
        \UART_BG16/N19 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_13  ( .A(\UART_BG16/iCounter[13] ), .B(
        \UART_BG16/add_54/carry [13]), .CO(\UART_BG16/add_54/carry [14]), .Z(
        \UART_BG16/N20 ) );
  notech_ha2 \UART_BG16/add_54/U1_1_14  ( .A(\UART_BG16/iCounter[14] ), .B(
        \UART_BG16/add_54/carry [14]), .CO(\UART_BG16/add_54/carry [15]), .Z(
        \UART_BG16/N21 ) );
  notech_and2 \UART_BG2/U9  ( .A(iBaudtick16x), .B(\UART_BG2/iCounter[0] ), 
        .Z(\UART_BG2/n1 ) );
  notech_and3 \UART_BG2/U8  ( .A(\UART_BG2/n1 ), .B(\UART_BG2/iCounter[1] ), 
        .C(\UART_BG2/iCounter[2] ), .Z(\UART_BG2/N14 ) );
  notech_and2 \UART_BG2/U7  ( .A(\UART_BG2/n1 ), .B(\UART_BG2/iCounter[1] ), 
        .Z(\UART_BG2/n2 ) );
  notech_xor2 \UART_BG2/U6  ( .A(\UART_BG2/iCounter[2] ), .B(\UART_BG2/n2 ), 
        .Z(\UART_BG2/n3 ) );
  notech_xor2 \UART_BG2/U5  ( .A(\UART_BG2/iCounter[1] ), .B(\UART_BG2/n1 ), 
        .Z(\UART_BG2/n4 ) );
  notech_xor2 \UART_BG2/U4  ( .A(\UART_BG2/iCounter[0] ), .B(iBaudtick16x), 
        .Z(\UART_BG2/n6 ) );
  notech_reg \UART_BG2/iQ_reg  ( .D(\UART_BG2/N14 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(iBaudtick2x) );
  notech_reg \UART_BG2/iCounter_reg[2]  ( .D(\UART_BG2/n3 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_BG2/iCounter[2] ) );
  notech_reg \UART_BG2/iCounter_reg[1]  ( .D(\UART_BG2/n4 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_BG2/iCounter[1] ) );
  notech_reg \UART_BG2/iCounter_reg[0]  ( .D(\UART_BG2/n6 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_BG2/iCounter[0] ) );
  notech_inv \UART_RCLK/U6  ( .A(\UART_RCLK/iDd ), .Z(\UART_RCLK/n1 ) );
  notech_and2 \UART_RCLK/U5  ( .A(RCLK), .B(\UART_RCLK/n1 ), .Z(iRCLK) );
  notech_reg \UART_RCLK/iDd_reg  ( .D(RCLK), .CP(CLK), .CD(\UART_IS_DSR/n1 ), 
        .Q(\UART_RCLK/iDd ) );
  notech_xor2 \UART_TXFF/U926  ( .A(\UART_TXFF/iWRAddr[1] ), .B(
        \UART_TXFF/N13 ), .Z(\UART_TXFF/n367 ) );
  notech_xor2 \UART_TXFF/U925  ( .A(\UART_TXFF/iWRAddr[5] ), .B(
        \UART_TXFF/N17 ), .Z(\UART_TXFF/n368 ) );
  notech_xor2 \UART_TXFF/U924  ( .A(\UART_TXFF/iWRAddr[0] ), .B(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n369 ) );
  notech_inv \UART_TXFF/U923  ( .A(\UART_TXFF/N14 ), .Z(\UART_TXFF/n232 ) );
  notech_xor2 \UART_TXFF/U922  ( .A(\UART_TXFF/n232 ), .B(
        \UART_TXFF/iWRAddr[2] ), .Z(\UART_TXFF/n371 ) );
  notech_inv \UART_TXFF/U921  ( .A(\UART_TXFF/N15 ), .Z(\UART_TXFF/n234 ) );
  notech_xor2 \UART_TXFF/U920  ( .A(\UART_TXFF/n234 ), .B(
        \UART_TXFF/iWRAddr[3] ), .Z(\UART_TXFF/n372 ) );
  notech_inv \UART_TXFF/U919  ( .A(\UART_TXFF/N16 ), .Z(\UART_TXFF/n236 ) );
  notech_xor2 \UART_TXFF/U918  ( .A(\UART_TXFF/n236 ), .B(
        \UART_TXFF/iWRAddr[4] ), .Z(\UART_TXFF/n373 ) );
  notech_nand3 \UART_TXFF/U917  ( .A(\UART_TXFF/n371 ), .B(\UART_TXFF/n372 ), 
        .C(\UART_TXFF/n373 ), .Z(\UART_TXFF/n370 ) );
  notech_nor4 \UART_TXFF/U916  ( .A(\UART_TXFF/n367 ), .B(\UART_TXFF/n368 ), 
        .C(\UART_TXFF/n369 ), .D(\UART_TXFF/n370 ), .Z(\UART_TXFF/n364 ) );
  notech_inv \UART_TXFF/U915  ( .A(\UART_TXFF/n364 ), .Z(\UART_TXFF/n366 ) );
  notech_inv \UART_TXFF/U914  ( .A(\UART_TXFF/iWRAddr[6] ), .Z(
        \UART_TXFF/n213 ) );
  notech_xor2 \UART_TXFF/U913  ( .A(\UART_TXFF/iRDAddr[6] ), .B(
        \UART_TXFF/n213 ), .Z(\UART_TXFF/n365 ) );
  notech_nor2 \UART_TXFF/U912  ( .A(\UART_TXFF/n366 ), .B(\UART_TXFF/n365 ), 
        .Z(iTXFIFO64Full) );
  notech_and2 \UART_TXFF/U911  ( .A(\UART_TXFF/n364 ), .B(\UART_TXFF/n365 ), 
        .Z(\UART_TXFF/N56 ) );
  notech_and3 \UART_TXFF/U910  ( .A(\UART_TXFF/USAGE[2] ), .B(
        \UART_TXFF/USAGE[0] ), .C(\UART_TXFF/USAGE[1] ), .Z(\UART_TXFF/n346 )
         );
  notech_inv \UART_TXFF/U909  ( .A(N169), .Z(\UART_TXFF/n363 ) );
  notech_nand3 \UART_TXFF/U907  ( .A(\UART_TXFF/n363 ), .B(iTXFIFORead), .C(
        n520), .Z(\UART_TXFF/n358 ) );
  notech_nor2 \UART_TXFF/U906  ( .A(iTXFIFO64Full), .B(\UART_TXFF/n363 ), .Z(
        \UART_TXFF/n287 ) );
  notech_or2 \UART_TXFF/U905  ( .A(\UART_TXFF/n287 ), .B(iFCR[2]), .Z(
        \UART_TXFF/n214 ) );
  notech_inv \UART_TXFF/U904  ( .A(iFCR[2]), .Z(\UART_TXFF/n228 ) );
  notech_nand2 \UART_TXFF/U903  ( .A(\UART_TXFF/n228 ), .B(iTXFIFORead), .Z(
        \UART_TXFF/n362 ) );
  notech_nand2 \UART_TXFF/U902  ( .A(\UART_TXFF/n214 ), .B(\UART_TXFF/n362 ), 
        .Z(\UART_TXFF/n361 ) );
  notech_nand2 \UART_TXFF/U901  ( .A(\UART_TXFF/n361 ), .B(\UART_TXFF/n358 ), 
        .Z(\UART_TXFF/n328 ) );
  notech_ao3 \UART_TXFF/U900  ( .A(\UART_TXFF/n358 ), .B(\UART_TXFF/n328 ), 
        .C(iFCR[2]), .Z(\UART_TXFF/n334 ) );
  notech_and3 \UART_TXFF/U899  ( .A(\UART_TXFF/n346 ), .B(\UART_TXFF/USAGE[3] ), .C(\UART_TXFF/n334 ), .Z(\UART_TXFF/n349 ) );
  notech_inv \UART_TXFF/U897  ( .A(\UART_TXFF/USAGE[1] ), .Z(\UART_TXFF/n359 )
         );
  notech_inv \UART_TXFF/U896  ( .A(\UART_TXFF/USAGE[0] ), .Z(\UART_TXFF/n360 )
         );
  notech_ao3 \UART_TXFF/U895  ( .A(\UART_TXFF/n359 ), .B(\UART_TXFF/n360 ), 
        .C(\UART_TXFF/USAGE[2] ), .Z(\UART_TXFF/n337 ) );
  notech_or2 \UART_TXFF/U894  ( .A(\UART_TXFF/n358 ), .B(iFCR[2]), .Z(
        \UART_TXFF/n330 ) );
  notech_inv \UART_TXFF/U893  ( .A(\UART_TXFF/n330 ), .Z(\UART_TXFF/n333 ) );
  notech_nao3 \UART_TXFF/U892  ( .C(\UART_TXFF/USAGE[3] ), .A(\UART_TXFF/n337 ), .B(\UART_TXFF/n333 ), .Z(\UART_TXFF/n343 ) );
  notech_nor2 \UART_TXFF/U891  ( .A(\UART_TXFF/n343 ), .B(\iTXFIFOUsage[4] ), 
        .Z(\UART_TXFF/n348 ) );
  notech_or2 \UART_TXFF/U889  ( .A(\UART_TXFF/n330 ), .B(\UART_TXFF/n337 ), 
        .Z(\UART_TXFF/n355 ) );
  notech_inv \UART_TXFF/U888  ( .A(\UART_TXFF/n334 ), .Z(\UART_TXFF/n329 ) );
  notech_or2 \UART_TXFF/U887  ( .A(\UART_TXFF/n329 ), .B(\UART_TXFF/n346 ), 
        .Z(\UART_TXFF/n356 ) );
  notech_and3 \UART_TXFF/U886  ( .A(\UART_TXFF/n355 ), .B(\UART_TXFF/n356 ), 
        .C(\UART_TXFF/n328 ), .Z(\UART_TXFF/n345 ) );
  notech_mux2 \UART_TXFF/U885  ( .A(\UART_TXFF/n329 ), .B(\UART_TXFF/n330 ), 
        .S(\UART_TXFF/USAGE[3] ), .Z(\UART_TXFF/n354 ) );
  notech_nand2 \UART_TXFF/U884  ( .A(\UART_TXFF/n345 ), .B(\UART_TXFF/n354 ), 
        .Z(\UART_TXFF/n350 ) );
  notech_mux2 \UART_TXFF/U880  ( .A(\UART_TXFF/n349 ), .B(\UART_TXFF/n350 ), 
        .S(\iTXFIFOUsage[4] ), .Z(\UART_TXFF/n347 ) );
  notech_or2 \UART_TXFF/U879  ( .A(\UART_TXFF/n347 ), .B(\UART_TXFF/n348 ), 
        .Z(\UART_TXFF/n1287 ) );
  notech_nand2 \UART_TXFF/U878  ( .A(\UART_TXFF/n334 ), .B(\UART_TXFF/n346 ), 
        .Z(\UART_TXFF/n344 ) );
  notech_mux2 \UART_TXFF/U877  ( .A(\UART_TXFF/n344 ), .B(\UART_TXFF/n345 ), 
        .S(\UART_TXFF/USAGE[3] ), .Z(\UART_TXFF/n342 ) );
  notech_nand2 \UART_TXFF/U876  ( .A(\UART_TXFF/n342 ), .B(\UART_TXFF/n343 ), 
        .Z(\UART_TXFF/n1288 ) );
  notech_nand3 \UART_TXFF/U875  ( .A(\UART_TXFF/n334 ), .B(
        \UART_TXFF/USAGE[0] ), .C(\UART_TXFF/USAGE[1] ), .Z(\UART_TXFF/n338 )
         );
  notech_mux2 \UART_TXFF/U874  ( .A(\UART_TXFF/n329 ), .B(\UART_TXFF/n330 ), 
        .S(\UART_TXFF/USAGE[0] ), .Z(\UART_TXFF/n341 ) );
  notech_nand2 \UART_TXFF/U873  ( .A(\UART_TXFF/n341 ), .B(\UART_TXFF/n328 ), 
        .Z(\UART_TXFF/n332 ) );
  notech_mux2 \UART_TXFF/U872  ( .A(\UART_TXFF/n334 ), .B(\UART_TXFF/n333 ), 
        .S(\UART_TXFF/USAGE[1] ), .Z(\UART_TXFF/n340 ) );
  notech_nor2 \UART_TXFF/U871  ( .A(\UART_TXFF/n332 ), .B(\UART_TXFF/n340 ), 
        .Z(\UART_TXFF/n339 ) );
  notech_mux2 \UART_TXFF/U870  ( .A(\UART_TXFF/n338 ), .B(\UART_TXFF/n339 ), 
        .S(\UART_TXFF/USAGE[2] ), .Z(\UART_TXFF/n335 ) );
  notech_nand2 \UART_TXFF/U869  ( .A(\UART_TXFF/n333 ), .B(\UART_TXFF/n337 ), 
        .Z(\UART_TXFF/n336 ) );
  notech_nand2 \UART_TXFF/U868  ( .A(\UART_TXFF/n335 ), .B(\UART_TXFF/n336 ), 
        .Z(\UART_TXFF/n1289 ) );
  notech_mux2 \UART_TXFF/U867  ( .A(\UART_TXFF/n333 ), .B(\UART_TXFF/n334 ), 
        .S(\UART_TXFF/USAGE[0] ), .Z(\UART_TXFF/n331 ) );
  notech_mux2 \UART_TXFF/U866  ( .A(\UART_TXFF/n331 ), .B(\UART_TXFF/n332 ), 
        .S(\UART_TXFF/USAGE[1] ), .Z(\UART_TXFF/n1290 ) );
  notech_nand2 \UART_TXFF/U865  ( .A(\UART_TXFF/n329 ), .B(\UART_TXFF/n330 ), 
        .Z(\UART_TXFF/n326 ) );
  notech_inv \UART_TXFF/U864  ( .A(\UART_TXFF/n328 ), .Z(\UART_TXFF/n327 ) );
  notech_mux2 \UART_TXFF/U863  ( .A(\UART_TXFF/n326 ), .B(\UART_TXFF/n327 ), 
        .S(\UART_TXFF/USAGE[0] ), .Z(\UART_TXFF/n1291 ) );
  notech_inv \UART_TXFF/U862  ( .A(\UART_TXFF/iWRAddr[3] ), .Z(
        \UART_TXFF/n222 ) );
  notech_ao3 \UART_TXFF/U860  ( .A(\UART_IF_CTS/n8 ), .B(\UART_TXFF/n287 ), 
        .C(\UART_TXFF/iWRAddr[5] ), .Z(\UART_TXFF/n297 ) );
  notech_ao3 \UART_TXFF/U859  ( .A(\UART_TXFF/n222 ), .B(\UART_TXFF/n297 ), 
        .C(\UART_TXFF/iWRAddr[4] ), .Z(\UART_TXFF/n317 ) );
  notech_inv \UART_TXFF/U858  ( .A(\UART_TXFF/iWRAddr[0] ), .Z(
        \UART_TXFF/n319 ) );
  notech_inv \UART_TXFF/U857  ( .A(\UART_TXFF/iWRAddr[2] ), .Z(
        \UART_TXFF/n220 ) );
  notech_inv \UART_TXFF/U856  ( .A(\UART_TXFF/iWRAddr[1] ), .Z(
        \UART_TXFF/n218 ) );
  notech_and3 \UART_TXFF/U855  ( .A(\UART_TXFF/n319 ), .B(\UART_TXFF/n220 ), 
        .C(\UART_TXFF/n218 ), .Z(\UART_TXFF/n258 ) );
  notech_and2 \UART_TXFF/U854  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n325 ) );
  notech_mux2 \UART_TXFF/U853  ( .A(\UART_TXFF/iFIFOMem[0][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1292 ) );
  notech_mux2 \UART_TXFF/U852  ( .A(\UART_TXFF/iFIFOMem[0][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1293 ) );
  notech_mux2 \UART_TXFF/U851  ( .A(\UART_TXFF/iFIFOMem[0][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1294 ) );
  notech_mux2 \UART_TXFF/U850  ( .A(\UART_TXFF/iFIFOMem[0][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1295 ) );
  notech_mux2 \UART_TXFF/U849  ( .A(\UART_TXFF/iFIFOMem[0][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1296 ) );
  notech_mux2 \UART_TXFF/U848  ( .A(\UART_TXFF/iFIFOMem[0][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1297 ) );
  notech_mux2 \UART_TXFF/U847  ( .A(\UART_TXFF/iFIFOMem[0][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1298 ) );
  notech_mux2 \UART_TXFF/U846  ( .A(\UART_TXFF/iFIFOMem[0][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n325 ), .Z(\UART_TXFF/n1299 ) );
  notech_and3 \UART_TXFF/U845  ( .A(\UART_TXFF/iWRAddr[0] ), .B(
        \UART_TXFF/n220 ), .C(\UART_TXFF/n218 ), .Z(\UART_TXFF/n256 ) );
  notech_and2 \UART_TXFF/U844  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n324 ) );
  notech_mux2 \UART_TXFF/U843  ( .A(\UART_TXFF/iFIFOMem[1][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1300 ) );
  notech_mux2 \UART_TXFF/U842  ( .A(\UART_TXFF/iFIFOMem[1][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1301 ) );
  notech_mux2 \UART_TXFF/U841  ( .A(\UART_TXFF/iFIFOMem[1][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1302 ) );
  notech_mux2 \UART_TXFF/U840  ( .A(\UART_TXFF/iFIFOMem[1][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1303 ) );
  notech_mux2 \UART_TXFF/U839  ( .A(\UART_TXFF/iFIFOMem[1][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1304 ) );
  notech_mux2 \UART_TXFF/U838  ( .A(\UART_TXFF/iFIFOMem[1][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1305 ) );
  notech_mux2 \UART_TXFF/U837  ( .A(\UART_TXFF/iFIFOMem[1][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1306 ) );
  notech_mux2 \UART_TXFF/U836  ( .A(\UART_TXFF/iFIFOMem[1][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n324 ), .Z(\UART_TXFF/n1307 ) );
  notech_and3 \UART_TXFF/U835  ( .A(\UART_TXFF/iWRAddr[1] ), .B(
        \UART_TXFF/n220 ), .C(\UART_TXFF/n319 ), .Z(\UART_TXFF/n254 ) );
  notech_and2 \UART_TXFF/U834  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n323 ) );
  notech_mux2 \UART_TXFF/U833  ( .A(\UART_TXFF/iFIFOMem[2][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1308 ) );
  notech_mux2 \UART_TXFF/U832  ( .A(\UART_TXFF/iFIFOMem[2][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1309 ) );
  notech_mux2 \UART_TXFF/U831  ( .A(\UART_TXFF/iFIFOMem[2][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1310 ) );
  notech_mux2 \UART_TXFF/U830  ( .A(\UART_TXFF/iFIFOMem[2][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1311 ) );
  notech_mux2 \UART_TXFF/U829  ( .A(\UART_TXFF/iFIFOMem[2][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1312 ) );
  notech_mux2 \UART_TXFF/U828  ( .A(\UART_TXFF/iFIFOMem[2][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1313 ) );
  notech_mux2 \UART_TXFF/U827  ( .A(\UART_TXFF/iFIFOMem[2][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1314 ) );
  notech_mux2 \UART_TXFF/U826  ( .A(\UART_TXFF/iFIFOMem[2][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n323 ), .Z(\UART_TXFF/n1315 ) );
  notech_and3 \UART_TXFF/U825  ( .A(\UART_TXFF/iWRAddr[0] ), .B(
        \UART_TXFF/iWRAddr[1] ), .C(\UART_TXFF/n220 ), .Z(\UART_TXFF/n252 ) );
  notech_and2 \UART_TXFF/U824  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n322 ) );
  notech_mux2 \UART_TXFF/U823  ( .A(\UART_TXFF/iFIFOMem[3][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1316 ) );
  notech_mux2 \UART_TXFF/U822  ( .A(\UART_TXFF/iFIFOMem[3][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1317 ) );
  notech_mux2 \UART_TXFF/U821  ( .A(\UART_TXFF/iFIFOMem[3][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1318 ) );
  notech_mux2 \UART_TXFF/U820  ( .A(\UART_TXFF/iFIFOMem[3][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1319 ) );
  notech_mux2 \UART_TXFF/U819  ( .A(\UART_TXFF/iFIFOMem[3][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1320 ) );
  notech_mux2 \UART_TXFF/U818  ( .A(\UART_TXFF/iFIFOMem[3][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1321 ) );
  notech_mux2 \UART_TXFF/U817  ( .A(\UART_TXFF/iFIFOMem[3][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1322 ) );
  notech_mux2 \UART_TXFF/U816  ( .A(\UART_TXFF/iFIFOMem[3][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n322 ), .Z(\UART_TXFF/n1323 ) );
  notech_and3 \UART_TXFF/U815  ( .A(\UART_TXFF/iWRAddr[2] ), .B(
        \UART_TXFF/n218 ), .C(\UART_TXFF/n319 ), .Z(\UART_TXFF/n250 ) );
  notech_and2 \UART_TXFF/U814  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n321 ) );
  notech_mux2 \UART_TXFF/U813  ( .A(\UART_TXFF/iFIFOMem[4][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1324 ) );
  notech_mux2 \UART_TXFF/U812  ( .A(\UART_TXFF/iFIFOMem[4][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1325 ) );
  notech_mux2 \UART_TXFF/U811  ( .A(\UART_TXFF/iFIFOMem[4][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1326 ) );
  notech_mux2 \UART_TXFF/U810  ( .A(\UART_TXFF/iFIFOMem[4][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1327 ) );
  notech_mux2 \UART_TXFF/U809  ( .A(\UART_TXFF/iFIFOMem[4][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1328 ) );
  notech_mux2 \UART_TXFF/U808  ( .A(\UART_TXFF/iFIFOMem[4][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1329 ) );
  notech_mux2 \UART_TXFF/U807  ( .A(\UART_TXFF/iFIFOMem[4][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1330 ) );
  notech_mux2 \UART_TXFF/U806  ( .A(\UART_TXFF/iFIFOMem[4][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n321 ), .Z(\UART_TXFF/n1331 ) );
  notech_and3 \UART_TXFF/U805  ( .A(\UART_TXFF/iWRAddr[0] ), .B(
        \UART_TXFF/iWRAddr[2] ), .C(\UART_TXFF/n218 ), .Z(\UART_TXFF/n248 ) );
  notech_and2 \UART_TXFF/U804  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n320 ) );
  notech_mux2 \UART_TXFF/U803  ( .A(\UART_TXFF/iFIFOMem[5][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1332 ) );
  notech_mux2 \UART_TXFF/U802  ( .A(\UART_TXFF/iFIFOMem[5][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1333 ) );
  notech_mux2 \UART_TXFF/U801  ( .A(\UART_TXFF/iFIFOMem[5][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1334 ) );
  notech_mux2 \UART_TXFF/U800  ( .A(\UART_TXFF/iFIFOMem[5][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1335 ) );
  notech_mux2 \UART_TXFF/U799  ( .A(\UART_TXFF/iFIFOMem[5][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1336 ) );
  notech_mux2 \UART_TXFF/U798  ( .A(\UART_TXFF/iFIFOMem[5][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1337 ) );
  notech_mux2 \UART_TXFF/U797  ( .A(\UART_TXFF/iFIFOMem[5][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1338 ) );
  notech_mux2 \UART_TXFF/U796  ( .A(\UART_TXFF/iFIFOMem[5][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n320 ), .Z(\UART_TXFF/n1339 ) );
  notech_and3 \UART_TXFF/U795  ( .A(\UART_TXFF/iWRAddr[1] ), .B(
        \UART_TXFF/iWRAddr[2] ), .C(\UART_TXFF/n319 ), .Z(\UART_TXFF/n246 ) );
  notech_and2 \UART_TXFF/U794  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n318 ) );
  notech_mux2 \UART_TXFF/U793  ( .A(\UART_TXFF/iFIFOMem[6][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1340 ) );
  notech_mux2 \UART_TXFF/U792  ( .A(\UART_TXFF/iFIFOMem[6][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1341 ) );
  notech_mux2 \UART_TXFF/U791  ( .A(\UART_TXFF/iFIFOMem[6][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1342 ) );
  notech_mux2 \UART_TXFF/U790  ( .A(\UART_TXFF/iFIFOMem[6][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1343 ) );
  notech_mux2 \UART_TXFF/U789  ( .A(\UART_TXFF/iFIFOMem[6][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1344 ) );
  notech_mux2 \UART_TXFF/U788  ( .A(\UART_TXFF/iFIFOMem[6][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1345 ) );
  notech_mux2 \UART_TXFF/U787  ( .A(\UART_TXFF/iFIFOMem[6][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1346 ) );
  notech_mux2 \UART_TXFF/U786  ( .A(\UART_TXFF/iFIFOMem[6][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n318 ), .Z(\UART_TXFF/n1347 ) );
  notech_and3 \UART_TXFF/U785  ( .A(\UART_TXFF/iWRAddr[0] ), .B(
        \UART_TXFF/iWRAddr[2] ), .C(\UART_TXFF/iWRAddr[1] ), .Z(
        \UART_TXFF/n244 ) );
  notech_and2 \UART_TXFF/U784  ( .A(\UART_TXFF/n317 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n316 ) );
  notech_mux2 \UART_TXFF/U783  ( .A(\UART_TXFF/iFIFOMem[7][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1348 ) );
  notech_mux2 \UART_TXFF/U782  ( .A(\UART_TXFF/iFIFOMem[7][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1349 ) );
  notech_mux2 \UART_TXFF/U781  ( .A(\UART_TXFF/iFIFOMem[7][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1350 ) );
  notech_mux2 \UART_TXFF/U780  ( .A(\UART_TXFF/iFIFOMem[7][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1351 ) );
  notech_mux2 \UART_TXFF/U779  ( .A(\UART_TXFF/iFIFOMem[7][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1352 ) );
  notech_mux2 \UART_TXFF/U778  ( .A(\UART_TXFF/iFIFOMem[7][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1353 ) );
  notech_mux2 \UART_TXFF/U777  ( .A(\UART_TXFF/iFIFOMem[7][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1354 ) );
  notech_mux2 \UART_TXFF/U776  ( .A(\UART_TXFF/iFIFOMem[7][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n316 ), .Z(\UART_TXFF/n1355 ) );
  notech_ao3 \UART_TXFF/U775  ( .A(\UART_TXFF/iWRAddr[3] ), .B(
        \UART_TXFF/n297 ), .C(\UART_TXFF/iWRAddr[4] ), .Z(\UART_TXFF/n308 ) );
  notech_and2 \UART_TXFF/U774  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n315 ) );
  notech_mux2 \UART_TXFF/U773  ( .A(\UART_TXFF/iFIFOMem[8][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1356 ) );
  notech_mux2 \UART_TXFF/U772  ( .A(\UART_TXFF/iFIFOMem[8][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1357 ) );
  notech_mux2 \UART_TXFF/U771  ( .A(\UART_TXFF/iFIFOMem[8][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1358 ) );
  notech_mux2 \UART_TXFF/U770  ( .A(\UART_TXFF/iFIFOMem[8][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1359 ) );
  notech_mux2 \UART_TXFF/U769  ( .A(\UART_TXFF/iFIFOMem[8][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1360 ) );
  notech_mux2 \UART_TXFF/U768  ( .A(\UART_TXFF/iFIFOMem[8][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1361 ) );
  notech_mux2 \UART_TXFF/U767  ( .A(\UART_TXFF/iFIFOMem[8][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1362 ) );
  notech_mux2 \UART_TXFF/U766  ( .A(\UART_TXFF/iFIFOMem[8][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n315 ), .Z(\UART_TXFF/n1363 ) );
  notech_and2 \UART_TXFF/U765  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n314 ) );
  notech_mux2 \UART_TXFF/U764  ( .A(\UART_TXFF/iFIFOMem[9][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1364 ) );
  notech_mux2 \UART_TXFF/U763  ( .A(\UART_TXFF/iFIFOMem[9][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1365 ) );
  notech_mux2 \UART_TXFF/U762  ( .A(\UART_TXFF/iFIFOMem[9][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1366 ) );
  notech_mux2 \UART_TXFF/U761  ( .A(\UART_TXFF/iFIFOMem[9][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1367 ) );
  notech_mux2 \UART_TXFF/U760  ( .A(\UART_TXFF/iFIFOMem[9][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1368 ) );
  notech_mux2 \UART_TXFF/U759  ( .A(\UART_TXFF/iFIFOMem[9][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1369 ) );
  notech_mux2 \UART_TXFF/U758  ( .A(\UART_TXFF/iFIFOMem[9][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1370 ) );
  notech_mux2 \UART_TXFF/U757  ( .A(\UART_TXFF/iFIFOMem[9][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n314 ), .Z(\UART_TXFF/n1371 ) );
  notech_and2 \UART_TXFF/U756  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n313 ) );
  notech_mux2 \UART_TXFF/U755  ( .A(\UART_TXFF/iFIFOMem[10][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1372 ) );
  notech_mux2 \UART_TXFF/U754  ( .A(\UART_TXFF/iFIFOMem[10][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1373 ) );
  notech_mux2 \UART_TXFF/U753  ( .A(\UART_TXFF/iFIFOMem[10][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1374 ) );
  notech_mux2 \UART_TXFF/U752  ( .A(\UART_TXFF/iFIFOMem[10][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1375 ) );
  notech_mux2 \UART_TXFF/U751  ( .A(\UART_TXFF/iFIFOMem[10][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1376 ) );
  notech_mux2 \UART_TXFF/U750  ( .A(\UART_TXFF/iFIFOMem[10][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1377 ) );
  notech_mux2 \UART_TXFF/U749  ( .A(\UART_TXFF/iFIFOMem[10][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1378 ) );
  notech_mux2 \UART_TXFF/U748  ( .A(\UART_TXFF/iFIFOMem[10][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n313 ), .Z(\UART_TXFF/n1379 ) );
  notech_and2 \UART_TXFF/U747  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n312 ) );
  notech_mux2 \UART_TXFF/U746  ( .A(\UART_TXFF/iFIFOMem[11][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1380 ) );
  notech_mux2 \UART_TXFF/U745  ( .A(\UART_TXFF/iFIFOMem[11][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1381 ) );
  notech_mux2 \UART_TXFF/U744  ( .A(\UART_TXFF/iFIFOMem[11][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1382 ) );
  notech_mux2 \UART_TXFF/U743  ( .A(\UART_TXFF/iFIFOMem[11][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1383 ) );
  notech_mux2 \UART_TXFF/U742  ( .A(\UART_TXFF/iFIFOMem[11][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1384 ) );
  notech_mux2 \UART_TXFF/U741  ( .A(\UART_TXFF/iFIFOMem[11][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1385 ) );
  notech_mux2 \UART_TXFF/U740  ( .A(\UART_TXFF/iFIFOMem[11][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1386 ) );
  notech_mux2 \UART_TXFF/U739  ( .A(\UART_TXFF/iFIFOMem[11][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n312 ), .Z(\UART_TXFF/n1387 ) );
  notech_and2 \UART_TXFF/U738  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n311 ) );
  notech_mux2 \UART_TXFF/U737  ( .A(\UART_TXFF/iFIFOMem[12][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1388 ) );
  notech_mux2 \UART_TXFF/U736  ( .A(\UART_TXFF/iFIFOMem[12][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1389 ) );
  notech_mux2 \UART_TXFF/U735  ( .A(\UART_TXFF/iFIFOMem[12][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1390 ) );
  notech_mux2 \UART_TXFF/U734  ( .A(\UART_TXFF/iFIFOMem[12][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1391 ) );
  notech_mux2 \UART_TXFF/U733  ( .A(\UART_TXFF/iFIFOMem[12][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1392 ) );
  notech_mux2 \UART_TXFF/U732  ( .A(\UART_TXFF/iFIFOMem[12][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1393 ) );
  notech_mux2 \UART_TXFF/U731  ( .A(\UART_TXFF/iFIFOMem[12][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1394 ) );
  notech_mux2 \UART_TXFF/U730  ( .A(\UART_TXFF/iFIFOMem[12][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n311 ), .Z(\UART_TXFF/n1395 ) );
  notech_and2 \UART_TXFF/U729  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n310 ) );
  notech_mux2 \UART_TXFF/U728  ( .A(\UART_TXFF/iFIFOMem[13][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1396 ) );
  notech_mux2 \UART_TXFF/U727  ( .A(\UART_TXFF/iFIFOMem[13][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1397 ) );
  notech_mux2 \UART_TXFF/U726  ( .A(\UART_TXFF/iFIFOMem[13][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1398 ) );
  notech_mux2 \UART_TXFF/U725  ( .A(\UART_TXFF/iFIFOMem[13][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1399 ) );
  notech_mux2 \UART_TXFF/U724  ( .A(\UART_TXFF/iFIFOMem[13][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1400 ) );
  notech_mux2 \UART_TXFF/U723  ( .A(\UART_TXFF/iFIFOMem[13][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1401 ) );
  notech_mux2 \UART_TXFF/U722  ( .A(\UART_TXFF/iFIFOMem[13][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1402 ) );
  notech_mux2 \UART_TXFF/U721  ( .A(\UART_TXFF/iFIFOMem[13][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n310 ), .Z(\UART_TXFF/n1403 ) );
  notech_and2 \UART_TXFF/U720  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n309 ) );
  notech_mux2 \UART_TXFF/U719  ( .A(\UART_TXFF/iFIFOMem[14][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1404 ) );
  notech_mux2 \UART_TXFF/U718  ( .A(\UART_TXFF/iFIFOMem[14][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1405 ) );
  notech_mux2 \UART_TXFF/U717  ( .A(\UART_TXFF/iFIFOMem[14][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1406 ) );
  notech_mux2 \UART_TXFF/U716  ( .A(\UART_TXFF/iFIFOMem[14][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1407 ) );
  notech_mux2 \UART_TXFF/U715  ( .A(\UART_TXFF/iFIFOMem[14][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1408 ) );
  notech_mux2 \UART_TXFF/U714  ( .A(\UART_TXFF/iFIFOMem[14][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1409 ) );
  notech_mux2 \UART_TXFF/U713  ( .A(\UART_TXFF/iFIFOMem[14][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1410 ) );
  notech_mux2 \UART_TXFF/U712  ( .A(\UART_TXFF/iFIFOMem[14][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n309 ), .Z(\UART_TXFF/n1411 ) );
  notech_and2 \UART_TXFF/U711  ( .A(\UART_TXFF/n308 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n307 ) );
  notech_mux2 \UART_TXFF/U710  ( .A(\UART_TXFF/iFIFOMem[15][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1412 ) );
  notech_mux2 \UART_TXFF/U709  ( .A(\UART_TXFF/iFIFOMem[15][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1413 ) );
  notech_mux2 \UART_TXFF/U708  ( .A(\UART_TXFF/iFIFOMem[15][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1414 ) );
  notech_mux2 \UART_TXFF/U707  ( .A(\UART_TXFF/iFIFOMem[15][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1415 ) );
  notech_mux2 \UART_TXFF/U706  ( .A(\UART_TXFF/iFIFOMem[15][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1416 ) );
  notech_mux2 \UART_TXFF/U705  ( .A(\UART_TXFF/iFIFOMem[15][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1417 ) );
  notech_mux2 \UART_TXFF/U704  ( .A(\UART_TXFF/iFIFOMem[15][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1418 ) );
  notech_mux2 \UART_TXFF/U703  ( .A(\UART_TXFF/iFIFOMem[15][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n307 ), .Z(\UART_TXFF/n1419 ) );
  notech_ao3 \UART_TXFF/U702  ( .A(\UART_TXFF/iWRAddr[4] ), .B(
        \UART_TXFF/n297 ), .C(\UART_TXFF/iWRAddr[3] ), .Z(\UART_TXFF/n299 ) );
  notech_and2 \UART_TXFF/U701  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n306 ) );
  notech_mux2 \UART_TXFF/U700  ( .A(\UART_TXFF/iFIFOMem[16][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1420 ) );
  notech_mux2 \UART_TXFF/U699  ( .A(\UART_TXFF/iFIFOMem[16][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1421 ) );
  notech_mux2 \UART_TXFF/U698  ( .A(\UART_TXFF/iFIFOMem[16][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1422 ) );
  notech_mux2 \UART_TXFF/U697  ( .A(\UART_TXFF/iFIFOMem[16][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1423 ) );
  notech_mux2 \UART_TXFF/U696  ( .A(\UART_TXFF/iFIFOMem[16][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1424 ) );
  notech_mux2 \UART_TXFF/U695  ( .A(\UART_TXFF/iFIFOMem[16][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1425 ) );
  notech_mux2 \UART_TXFF/U694  ( .A(\UART_TXFF/iFIFOMem[16][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1426 ) );
  notech_mux2 \UART_TXFF/U693  ( .A(\UART_TXFF/iFIFOMem[16][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n306 ), .Z(\UART_TXFF/n1427 ) );
  notech_and2 \UART_TXFF/U692  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n305 ) );
  notech_mux2 \UART_TXFF/U691  ( .A(\UART_TXFF/iFIFOMem[17][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1428 ) );
  notech_mux2 \UART_TXFF/U690  ( .A(\UART_TXFF/iFIFOMem[17][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1429 ) );
  notech_mux2 \UART_TXFF/U689  ( .A(\UART_TXFF/iFIFOMem[17][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1430 ) );
  notech_mux2 \UART_TXFF/U688  ( .A(\UART_TXFF/iFIFOMem[17][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1431 ) );
  notech_mux2 \UART_TXFF/U687  ( .A(\UART_TXFF/iFIFOMem[17][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1432 ) );
  notech_mux2 \UART_TXFF/U686  ( .A(\UART_TXFF/iFIFOMem[17][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1433 ) );
  notech_mux2 \UART_TXFF/U685  ( .A(\UART_TXFF/iFIFOMem[17][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1434 ) );
  notech_mux2 \UART_TXFF/U684  ( .A(\UART_TXFF/iFIFOMem[17][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n305 ), .Z(\UART_TXFF/n1435 ) );
  notech_and2 \UART_TXFF/U683  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n304 ) );
  notech_mux2 \UART_TXFF/U682  ( .A(\UART_TXFF/iFIFOMem[18][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1436 ) );
  notech_mux2 \UART_TXFF/U681  ( .A(\UART_TXFF/iFIFOMem[18][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1437 ) );
  notech_mux2 \UART_TXFF/U680  ( .A(\UART_TXFF/iFIFOMem[18][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1438 ) );
  notech_mux2 \UART_TXFF/U679  ( .A(\UART_TXFF/iFIFOMem[18][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1439 ) );
  notech_mux2 \UART_TXFF/U678  ( .A(\UART_TXFF/iFIFOMem[18][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1440 ) );
  notech_mux2 \UART_TXFF/U677  ( .A(\UART_TXFF/iFIFOMem[18][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1441 ) );
  notech_mux2 \UART_TXFF/U676  ( .A(\UART_TXFF/iFIFOMem[18][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1442 ) );
  notech_mux2 \UART_TXFF/U675  ( .A(\UART_TXFF/iFIFOMem[18][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n304 ), .Z(\UART_TXFF/n1443 ) );
  notech_and2 \UART_TXFF/U674  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n303 ) );
  notech_mux2 \UART_TXFF/U673  ( .A(\UART_TXFF/iFIFOMem[19][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1444 ) );
  notech_mux2 \UART_TXFF/U672  ( .A(\UART_TXFF/iFIFOMem[19][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1445 ) );
  notech_mux2 \UART_TXFF/U671  ( .A(\UART_TXFF/iFIFOMem[19][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1446 ) );
  notech_mux2 \UART_TXFF/U670  ( .A(\UART_TXFF/iFIFOMem[19][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1447 ) );
  notech_mux2 \UART_TXFF/U669  ( .A(\UART_TXFF/iFIFOMem[19][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1448 ) );
  notech_mux2 \UART_TXFF/U668  ( .A(\UART_TXFF/iFIFOMem[19][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1449 ) );
  notech_mux2 \UART_TXFF/U667  ( .A(\UART_TXFF/iFIFOMem[19][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1450 ) );
  notech_mux2 \UART_TXFF/U666  ( .A(\UART_TXFF/iFIFOMem[19][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n303 ), .Z(\UART_TXFF/n1451 ) );
  notech_and2 \UART_TXFF/U665  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n302 ) );
  notech_mux2 \UART_TXFF/U664  ( .A(\UART_TXFF/iFIFOMem[20][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1452 ) );
  notech_mux2 \UART_TXFF/U663  ( .A(\UART_TXFF/iFIFOMem[20][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1453 ) );
  notech_mux2 \UART_TXFF/U662  ( .A(\UART_TXFF/iFIFOMem[20][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1454 ) );
  notech_mux2 \UART_TXFF/U661  ( .A(\UART_TXFF/iFIFOMem[20][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1455 ) );
  notech_mux2 \UART_TXFF/U660  ( .A(\UART_TXFF/iFIFOMem[20][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1456 ) );
  notech_mux2 \UART_TXFF/U659  ( .A(\UART_TXFF/iFIFOMem[20][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1457 ) );
  notech_mux2 \UART_TXFF/U658  ( .A(\UART_TXFF/iFIFOMem[20][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1458 ) );
  notech_mux2 \UART_TXFF/U657  ( .A(\UART_TXFF/iFIFOMem[20][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n302 ), .Z(\UART_TXFF/n1459 ) );
  notech_and2 \UART_TXFF/U656  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n301 ) );
  notech_mux2 \UART_TXFF/U655  ( .A(\UART_TXFF/iFIFOMem[21][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1460 ) );
  notech_mux2 \UART_TXFF/U654  ( .A(\UART_TXFF/iFIFOMem[21][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1461 ) );
  notech_mux2 \UART_TXFF/U653  ( .A(\UART_TXFF/iFIFOMem[21][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1462 ) );
  notech_mux2 \UART_TXFF/U652  ( .A(\UART_TXFF/iFIFOMem[21][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1463 ) );
  notech_mux2 \UART_TXFF/U651  ( .A(\UART_TXFF/iFIFOMem[21][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1464 ) );
  notech_mux2 \UART_TXFF/U650  ( .A(\UART_TXFF/iFIFOMem[21][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1465 ) );
  notech_mux2 \UART_TXFF/U649  ( .A(\UART_TXFF/iFIFOMem[21][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1466 ) );
  notech_mux2 \UART_TXFF/U648  ( .A(\UART_TXFF/iFIFOMem[21][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n301 ), .Z(\UART_TXFF/n1467 ) );
  notech_and2 \UART_TXFF/U647  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n300 ) );
  notech_mux2 \UART_TXFF/U646  ( .A(\UART_TXFF/iFIFOMem[22][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1468 ) );
  notech_mux2 \UART_TXFF/U645  ( .A(\UART_TXFF/iFIFOMem[22][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1469 ) );
  notech_mux2 \UART_TXFF/U644  ( .A(\UART_TXFF/iFIFOMem[22][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1470 ) );
  notech_mux2 \UART_TXFF/U643  ( .A(\UART_TXFF/iFIFOMem[22][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1471 ) );
  notech_mux2 \UART_TXFF/U642  ( .A(\UART_TXFF/iFIFOMem[22][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1472 ) );
  notech_mux2 \UART_TXFF/U641  ( .A(\UART_TXFF/iFIFOMem[22][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1473 ) );
  notech_mux2 \UART_TXFF/U640  ( .A(\UART_TXFF/iFIFOMem[22][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1474 ) );
  notech_mux2 \UART_TXFF/U639  ( .A(\UART_TXFF/iFIFOMem[22][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n300 ), .Z(\UART_TXFF/n1475 ) );
  notech_and2 \UART_TXFF/U638  ( .A(\UART_TXFF/n299 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n298 ) );
  notech_mux2 \UART_TXFF/U637  ( .A(\UART_TXFF/iFIFOMem[23][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1476 ) );
  notech_mux2 \UART_TXFF/U636  ( .A(\UART_TXFF/iFIFOMem[23][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1477 ) );
  notech_mux2 \UART_TXFF/U635  ( .A(\UART_TXFF/iFIFOMem[23][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1478 ) );
  notech_mux2 \UART_TXFF/U634  ( .A(\UART_TXFF/iFIFOMem[23][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1479 ) );
  notech_mux2 \UART_TXFF/U633  ( .A(\UART_TXFF/iFIFOMem[23][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1480 ) );
  notech_mux2 \UART_TXFF/U632  ( .A(\UART_TXFF/iFIFOMem[23][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1481 ) );
  notech_mux2 \UART_TXFF/U631  ( .A(\UART_TXFF/iFIFOMem[23][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1482 ) );
  notech_mux2 \UART_TXFF/U630  ( .A(\UART_TXFF/iFIFOMem[23][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n298 ), .Z(\UART_TXFF/n1483 ) );
  notech_ao3 \UART_TXFF/U629  ( .A(\UART_TXFF/iWRAddr[4] ), .B(
        \UART_TXFF/n297 ), .C(\UART_TXFF/n222 ), .Z(\UART_TXFF/n289 ) );
  notech_and2 \UART_TXFF/U628  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n296 ) );
  notech_mux2 \UART_TXFF/U627  ( .A(\UART_TXFF/iFIFOMem[24][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1484 ) );
  notech_mux2 \UART_TXFF/U626  ( .A(\UART_TXFF/iFIFOMem[24][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1485 ) );
  notech_mux2 \UART_TXFF/U625  ( .A(\UART_TXFF/iFIFOMem[24][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1486 ) );
  notech_mux2 \UART_TXFF/U624  ( .A(\UART_TXFF/iFIFOMem[24][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1487 ) );
  notech_mux2 \UART_TXFF/U623  ( .A(\UART_TXFF/iFIFOMem[24][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1488 ) );
  notech_mux2 \UART_TXFF/U622  ( .A(\UART_TXFF/iFIFOMem[24][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1489 ) );
  notech_mux2 \UART_TXFF/U621  ( .A(\UART_TXFF/iFIFOMem[24][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1490 ) );
  notech_mux2 \UART_TXFF/U620  ( .A(\UART_TXFF/iFIFOMem[24][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n296 ), .Z(\UART_TXFF/n1491 ) );
  notech_and2 \UART_TXFF/U619  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n295 ) );
  notech_mux2 \UART_TXFF/U618  ( .A(\UART_TXFF/iFIFOMem[25][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1492 ) );
  notech_mux2 \UART_TXFF/U617  ( .A(\UART_TXFF/iFIFOMem[25][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1493 ) );
  notech_mux2 \UART_TXFF/U616  ( .A(\UART_TXFF/iFIFOMem[25][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1494 ) );
  notech_mux2 \UART_TXFF/U615  ( .A(\UART_TXFF/iFIFOMem[25][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1495 ) );
  notech_mux2 \UART_TXFF/U614  ( .A(\UART_TXFF/iFIFOMem[25][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1496 ) );
  notech_mux2 \UART_TXFF/U613  ( .A(\UART_TXFF/iFIFOMem[25][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1497 ) );
  notech_mux2 \UART_TXFF/U612  ( .A(\UART_TXFF/iFIFOMem[25][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1498 ) );
  notech_mux2 \UART_TXFF/U611  ( .A(\UART_TXFF/iFIFOMem[25][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n295 ), .Z(\UART_TXFF/n1499 ) );
  notech_and2 \UART_TXFF/U610  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n294 ) );
  notech_mux2 \UART_TXFF/U609  ( .A(\UART_TXFF/iFIFOMem[26][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1500 ) );
  notech_mux2 \UART_TXFF/U608  ( .A(\UART_TXFF/iFIFOMem[26][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1501 ) );
  notech_mux2 \UART_TXFF/U607  ( .A(\UART_TXFF/iFIFOMem[26][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1502 ) );
  notech_mux2 \UART_TXFF/U606  ( .A(\UART_TXFF/iFIFOMem[26][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1503 ) );
  notech_mux2 \UART_TXFF/U605  ( .A(\UART_TXFF/iFIFOMem[26][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1504 ) );
  notech_mux2 \UART_TXFF/U604  ( .A(\UART_TXFF/iFIFOMem[26][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1505 ) );
  notech_mux2 \UART_TXFF/U603  ( .A(\UART_TXFF/iFIFOMem[26][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1506 ) );
  notech_mux2 \UART_TXFF/U602  ( .A(\UART_TXFF/iFIFOMem[26][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n294 ), .Z(\UART_TXFF/n1507 ) );
  notech_and2 \UART_TXFF/U601  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n293 ) );
  notech_mux2 \UART_TXFF/U600  ( .A(\UART_TXFF/iFIFOMem[27][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1508 ) );
  notech_mux2 \UART_TXFF/U599  ( .A(\UART_TXFF/iFIFOMem[27][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1509 ) );
  notech_mux2 \UART_TXFF/U598  ( .A(\UART_TXFF/iFIFOMem[27][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1510 ) );
  notech_mux2 \UART_TXFF/U597  ( .A(\UART_TXFF/iFIFOMem[27][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1511 ) );
  notech_mux2 \UART_TXFF/U596  ( .A(\UART_TXFF/iFIFOMem[27][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1512 ) );
  notech_mux2 \UART_TXFF/U595  ( .A(\UART_TXFF/iFIFOMem[27][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1513 ) );
  notech_mux2 \UART_TXFF/U594  ( .A(\UART_TXFF/iFIFOMem[27][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1514 ) );
  notech_mux2 \UART_TXFF/U593  ( .A(\UART_TXFF/iFIFOMem[27][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n293 ), .Z(\UART_TXFF/n1515 ) );
  notech_and2 \UART_TXFF/U592  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n292 ) );
  notech_mux2 \UART_TXFF/U591  ( .A(\UART_TXFF/iFIFOMem[28][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1516 ) );
  notech_mux2 \UART_TXFF/U590  ( .A(\UART_TXFF/iFIFOMem[28][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1517 ) );
  notech_mux2 \UART_TXFF/U589  ( .A(\UART_TXFF/iFIFOMem[28][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1518 ) );
  notech_mux2 \UART_TXFF/U588  ( .A(\UART_TXFF/iFIFOMem[28][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1519 ) );
  notech_mux2 \UART_TXFF/U587  ( .A(\UART_TXFF/iFIFOMem[28][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1520 ) );
  notech_mux2 \UART_TXFF/U586  ( .A(\UART_TXFF/iFIFOMem[28][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1521 ) );
  notech_mux2 \UART_TXFF/U585  ( .A(\UART_TXFF/iFIFOMem[28][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1522 ) );
  notech_mux2 \UART_TXFF/U584  ( .A(\UART_TXFF/iFIFOMem[28][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n292 ), .Z(\UART_TXFF/n1523 ) );
  notech_and2 \UART_TXFF/U583  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n291 ) );
  notech_mux2 \UART_TXFF/U582  ( .A(\UART_TXFF/iFIFOMem[29][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1524 ) );
  notech_mux2 \UART_TXFF/U581  ( .A(\UART_TXFF/iFIFOMem[29][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1525 ) );
  notech_mux2 \UART_TXFF/U580  ( .A(\UART_TXFF/iFIFOMem[29][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1526 ) );
  notech_mux2 \UART_TXFF/U579  ( .A(\UART_TXFF/iFIFOMem[29][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1527 ) );
  notech_mux2 \UART_TXFF/U578  ( .A(\UART_TXFF/iFIFOMem[29][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1528 ) );
  notech_mux2 \UART_TXFF/U577  ( .A(\UART_TXFF/iFIFOMem[29][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1529 ) );
  notech_mux2 \UART_TXFF/U576  ( .A(\UART_TXFF/iFIFOMem[29][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1530 ) );
  notech_mux2 \UART_TXFF/U575  ( .A(\UART_TXFF/iFIFOMem[29][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n291 ), .Z(\UART_TXFF/n1531 ) );
  notech_and2 \UART_TXFF/U574  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n290 ) );
  notech_mux2 \UART_TXFF/U573  ( .A(\UART_TXFF/iFIFOMem[30][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1532 ) );
  notech_mux2 \UART_TXFF/U572  ( .A(\UART_TXFF/iFIFOMem[30][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1533 ) );
  notech_mux2 \UART_TXFF/U571  ( .A(\UART_TXFF/iFIFOMem[30][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1534 ) );
  notech_mux2 \UART_TXFF/U570  ( .A(\UART_TXFF/iFIFOMem[30][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1535 ) );
  notech_mux2 \UART_TXFF/U569  ( .A(\UART_TXFF/iFIFOMem[30][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1536 ) );
  notech_mux2 \UART_TXFF/U568  ( .A(\UART_TXFF/iFIFOMem[30][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1537 ) );
  notech_mux2 \UART_TXFF/U567  ( .A(\UART_TXFF/iFIFOMem[30][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1538 ) );
  notech_mux2 \UART_TXFF/U566  ( .A(\UART_TXFF/iFIFOMem[30][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n290 ), .Z(\UART_TXFF/n1539 ) );
  notech_and2 \UART_TXFF/U565  ( .A(\UART_TXFF/n289 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n288 ) );
  notech_mux2 \UART_TXFF/U564  ( .A(\UART_TXFF/iFIFOMem[31][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1540 ) );
  notech_mux2 \UART_TXFF/U563  ( .A(\UART_TXFF/iFIFOMem[31][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1541 ) );
  notech_mux2 \UART_TXFF/U562  ( .A(\UART_TXFF/iFIFOMem[31][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1542 ) );
  notech_mux2 \UART_TXFF/U561  ( .A(\UART_TXFF/iFIFOMem[31][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1543 ) );
  notech_mux2 \UART_TXFF/U560  ( .A(\UART_TXFF/iFIFOMem[31][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1544 ) );
  notech_mux2 \UART_TXFF/U559  ( .A(\UART_TXFF/iFIFOMem[31][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1545 ) );
  notech_mux2 \UART_TXFF/U558  ( .A(\UART_TXFF/iFIFOMem[31][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1546 ) );
  notech_mux2 \UART_TXFF/U557  ( .A(\UART_TXFF/iFIFOMem[31][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n288 ), .Z(\UART_TXFF/n1547 ) );
  notech_ao3 \UART_TXFF/U556  ( .A(\UART_TXFF/iWRAddr[5] ), .B(
        \UART_TXFF/n287 ), .C(RST), .Z(\UART_TXFF/n259 ) );
  notech_ao3 \UART_TXFF/U555  ( .A(\UART_TXFF/n222 ), .B(\UART_TXFF/n259 ), 
        .C(\UART_TXFF/iWRAddr[4] ), .Z(\UART_TXFF/n279 ) );
  notech_and2 \UART_TXFF/U554  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n286 ) );
  notech_mux2 \UART_TXFF/U553  ( .A(\UART_TXFF/iFIFOMem[32][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1548 ) );
  notech_mux2 \UART_TXFF/U552  ( .A(\UART_TXFF/iFIFOMem[32][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1549 ) );
  notech_mux2 \UART_TXFF/U551  ( .A(\UART_TXFF/iFIFOMem[32][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1550 ) );
  notech_mux2 \UART_TXFF/U550  ( .A(\UART_TXFF/iFIFOMem[32][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1551 ) );
  notech_mux2 \UART_TXFF/U549  ( .A(\UART_TXFF/iFIFOMem[32][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1552 ) );
  notech_mux2 \UART_TXFF/U548  ( .A(\UART_TXFF/iFIFOMem[32][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1553 ) );
  notech_mux2 \UART_TXFF/U547  ( .A(\UART_TXFF/iFIFOMem[32][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1554 ) );
  notech_mux2 \UART_TXFF/U546  ( .A(\UART_TXFF/iFIFOMem[32][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n286 ), .Z(\UART_TXFF/n1555 ) );
  notech_and2 \UART_TXFF/U545  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n285 ) );
  notech_mux2 \UART_TXFF/U544  ( .A(\UART_TXFF/iFIFOMem[33][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1556 ) );
  notech_mux2 \UART_TXFF/U543  ( .A(\UART_TXFF/iFIFOMem[33][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1557 ) );
  notech_mux2 \UART_TXFF/U542  ( .A(\UART_TXFF/iFIFOMem[33][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1558 ) );
  notech_mux2 \UART_TXFF/U541  ( .A(\UART_TXFF/iFIFOMem[33][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1559 ) );
  notech_mux2 \UART_TXFF/U540  ( .A(\UART_TXFF/iFIFOMem[33][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1560 ) );
  notech_mux2 \UART_TXFF/U539  ( .A(\UART_TXFF/iFIFOMem[33][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1561 ) );
  notech_mux2 \UART_TXFF/U538  ( .A(\UART_TXFF/iFIFOMem[33][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1562 ) );
  notech_mux2 \UART_TXFF/U537  ( .A(\UART_TXFF/iFIFOMem[33][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n285 ), .Z(\UART_TXFF/n1563 ) );
  notech_and2 \UART_TXFF/U536  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n284 ) );
  notech_mux2 \UART_TXFF/U535  ( .A(\UART_TXFF/iFIFOMem[34][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1564 ) );
  notech_mux2 \UART_TXFF/U534  ( .A(\UART_TXFF/iFIFOMem[34][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1565 ) );
  notech_mux2 \UART_TXFF/U533  ( .A(\UART_TXFF/iFIFOMem[34][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1566 ) );
  notech_mux2 \UART_TXFF/U532  ( .A(\UART_TXFF/iFIFOMem[34][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1567 ) );
  notech_mux2 \UART_TXFF/U531  ( .A(\UART_TXFF/iFIFOMem[34][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1568 ) );
  notech_mux2 \UART_TXFF/U530  ( .A(\UART_TXFF/iFIFOMem[34][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1569 ) );
  notech_mux2 \UART_TXFF/U529  ( .A(\UART_TXFF/iFIFOMem[34][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1570 ) );
  notech_mux2 \UART_TXFF/U528  ( .A(\UART_TXFF/iFIFOMem[34][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n284 ), .Z(\UART_TXFF/n1571 ) );
  notech_and2 \UART_TXFF/U527  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n283 ) );
  notech_mux2 \UART_TXFF/U526  ( .A(\UART_TXFF/iFIFOMem[35][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1572 ) );
  notech_mux2 \UART_TXFF/U525  ( .A(\UART_TXFF/iFIFOMem[35][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1573 ) );
  notech_mux2 \UART_TXFF/U524  ( .A(\UART_TXFF/iFIFOMem[35][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1574 ) );
  notech_mux2 \UART_TXFF/U523  ( .A(\UART_TXFF/iFIFOMem[35][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1575 ) );
  notech_mux2 \UART_TXFF/U522  ( .A(\UART_TXFF/iFIFOMem[35][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1576 ) );
  notech_mux2 \UART_TXFF/U521  ( .A(\UART_TXFF/iFIFOMem[35][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1577 ) );
  notech_mux2 \UART_TXFF/U520  ( .A(\UART_TXFF/iFIFOMem[35][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1578 ) );
  notech_mux2 \UART_TXFF/U519  ( .A(\UART_TXFF/iFIFOMem[35][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n283 ), .Z(\UART_TXFF/n1579 ) );
  notech_and2 \UART_TXFF/U518  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n282 ) );
  notech_mux2 \UART_TXFF/U517  ( .A(\UART_TXFF/iFIFOMem[36][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1580 ) );
  notech_mux2 \UART_TXFF/U516  ( .A(\UART_TXFF/iFIFOMem[36][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1581 ) );
  notech_mux2 \UART_TXFF/U515  ( .A(\UART_TXFF/iFIFOMem[36][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1582 ) );
  notech_mux2 \UART_TXFF/U514  ( .A(\UART_TXFF/iFIFOMem[36][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1583 ) );
  notech_mux2 \UART_TXFF/U513  ( .A(\UART_TXFF/iFIFOMem[36][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1584 ) );
  notech_mux2 \UART_TXFF/U512  ( .A(\UART_TXFF/iFIFOMem[36][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1585 ) );
  notech_mux2 \UART_TXFF/U511  ( .A(\UART_TXFF/iFIFOMem[36][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1586 ) );
  notech_mux2 \UART_TXFF/U510  ( .A(\UART_TXFF/iFIFOMem[36][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n282 ), .Z(\UART_TXFF/n1587 ) );
  notech_and2 \UART_TXFF/U509  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n281 ) );
  notech_mux2 \UART_TXFF/U508  ( .A(\UART_TXFF/iFIFOMem[37][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1588 ) );
  notech_mux2 \UART_TXFF/U507  ( .A(\UART_TXFF/iFIFOMem[37][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1589 ) );
  notech_mux2 \UART_TXFF/U506  ( .A(\UART_TXFF/iFIFOMem[37][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1590 ) );
  notech_mux2 \UART_TXFF/U505  ( .A(\UART_TXFF/iFIFOMem[37][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1591 ) );
  notech_mux2 \UART_TXFF/U504  ( .A(\UART_TXFF/iFIFOMem[37][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1592 ) );
  notech_mux2 \UART_TXFF/U503  ( .A(\UART_TXFF/iFIFOMem[37][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1593 ) );
  notech_mux2 \UART_TXFF/U502  ( .A(\UART_TXFF/iFIFOMem[37][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1594 ) );
  notech_mux2 \UART_TXFF/U501  ( .A(\UART_TXFF/iFIFOMem[37][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n281 ), .Z(\UART_TXFF/n1595 ) );
  notech_and2 \UART_TXFF/U500  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n280 ) );
  notech_mux2 \UART_TXFF/U499  ( .A(\UART_TXFF/iFIFOMem[38][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1596 ) );
  notech_mux2 \UART_TXFF/U498  ( .A(\UART_TXFF/iFIFOMem[38][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1597 ) );
  notech_mux2 \UART_TXFF/U497  ( .A(\UART_TXFF/iFIFOMem[38][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1598 ) );
  notech_mux2 \UART_TXFF/U496  ( .A(\UART_TXFF/iFIFOMem[38][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1599 ) );
  notech_mux2 \UART_TXFF/U495  ( .A(\UART_TXFF/iFIFOMem[38][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1600 ) );
  notech_mux2 \UART_TXFF/U494  ( .A(\UART_TXFF/iFIFOMem[38][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1601 ) );
  notech_mux2 \UART_TXFF/U493  ( .A(\UART_TXFF/iFIFOMem[38][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1602 ) );
  notech_mux2 \UART_TXFF/U492  ( .A(\UART_TXFF/iFIFOMem[38][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n280 ), .Z(\UART_TXFF/n1603 ) );
  notech_and2 \UART_TXFF/U491  ( .A(\UART_TXFF/n279 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n278 ) );
  notech_mux2 \UART_TXFF/U490  ( .A(\UART_TXFF/iFIFOMem[39][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1604 ) );
  notech_mux2 \UART_TXFF/U489  ( .A(\UART_TXFF/iFIFOMem[39][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1605 ) );
  notech_mux2 \UART_TXFF/U488  ( .A(\UART_TXFF/iFIFOMem[39][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1606 ) );
  notech_mux2 \UART_TXFF/U487  ( .A(\UART_TXFF/iFIFOMem[39][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1607 ) );
  notech_mux2 \UART_TXFF/U486  ( .A(\UART_TXFF/iFIFOMem[39][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1608 ) );
  notech_mux2 \UART_TXFF/U485  ( .A(\UART_TXFF/iFIFOMem[39][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1609 ) );
  notech_mux2 \UART_TXFF/U484  ( .A(\UART_TXFF/iFIFOMem[39][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1610 ) );
  notech_mux2 \UART_TXFF/U483  ( .A(\UART_TXFF/iFIFOMem[39][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n278 ), .Z(\UART_TXFF/n1611 ) );
  notech_ao3 \UART_TXFF/U482  ( .A(\UART_TXFF/iWRAddr[3] ), .B(
        \UART_TXFF/n259 ), .C(\UART_TXFF/iWRAddr[4] ), .Z(\UART_TXFF/n270 ) );
  notech_and2 \UART_TXFF/U481  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n277 ) );
  notech_mux2 \UART_TXFF/U480  ( .A(\UART_TXFF/iFIFOMem[40][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1612 ) );
  notech_mux2 \UART_TXFF/U479  ( .A(\UART_TXFF/iFIFOMem[40][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1613 ) );
  notech_mux2 \UART_TXFF/U478  ( .A(\UART_TXFF/iFIFOMem[40][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1614 ) );
  notech_mux2 \UART_TXFF/U477  ( .A(\UART_TXFF/iFIFOMem[40][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1615 ) );
  notech_mux2 \UART_TXFF/U476  ( .A(\UART_TXFF/iFIFOMem[40][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1616 ) );
  notech_mux2 \UART_TXFF/U475  ( .A(\UART_TXFF/iFIFOMem[40][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1617 ) );
  notech_mux2 \UART_TXFF/U474  ( .A(\UART_TXFF/iFIFOMem[40][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1618 ) );
  notech_mux2 \UART_TXFF/U473  ( .A(\UART_TXFF/iFIFOMem[40][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n277 ), .Z(\UART_TXFF/n1619 ) );
  notech_and2 \UART_TXFF/U472  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n276 ) );
  notech_mux2 \UART_TXFF/U471  ( .A(\UART_TXFF/iFIFOMem[41][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1620 ) );
  notech_mux2 \UART_TXFF/U470  ( .A(\UART_TXFF/iFIFOMem[41][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1621 ) );
  notech_mux2 \UART_TXFF/U469  ( .A(\UART_TXFF/iFIFOMem[41][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1622 ) );
  notech_mux2 \UART_TXFF/U468  ( .A(\UART_TXFF/iFIFOMem[41][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1623 ) );
  notech_mux2 \UART_TXFF/U467  ( .A(\UART_TXFF/iFIFOMem[41][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1624 ) );
  notech_mux2 \UART_TXFF/U466  ( .A(\UART_TXFF/iFIFOMem[41][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1625 ) );
  notech_mux2 \UART_TXFF/U465  ( .A(\UART_TXFF/iFIFOMem[41][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1626 ) );
  notech_mux2 \UART_TXFF/U464  ( .A(\UART_TXFF/iFIFOMem[41][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n276 ), .Z(\UART_TXFF/n1627 ) );
  notech_and2 \UART_TXFF/U463  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n275 ) );
  notech_mux2 \UART_TXFF/U462  ( .A(\UART_TXFF/iFIFOMem[42][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1628 ) );
  notech_mux2 \UART_TXFF/U461  ( .A(\UART_TXFF/iFIFOMem[42][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1629 ) );
  notech_mux2 \UART_TXFF/U460  ( .A(\UART_TXFF/iFIFOMem[42][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1630 ) );
  notech_mux2 \UART_TXFF/U459  ( .A(\UART_TXFF/iFIFOMem[42][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1631 ) );
  notech_mux2 \UART_TXFF/U458  ( .A(\UART_TXFF/iFIFOMem[42][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1632 ) );
  notech_mux2 \UART_TXFF/U457  ( .A(\UART_TXFF/iFIFOMem[42][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1633 ) );
  notech_mux2 \UART_TXFF/U456  ( .A(\UART_TXFF/iFIFOMem[42][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1634 ) );
  notech_mux2 \UART_TXFF/U455  ( .A(\UART_TXFF/iFIFOMem[42][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n275 ), .Z(\UART_TXFF/n1635 ) );
  notech_and2 \UART_TXFF/U454  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n274 ) );
  notech_mux2 \UART_TXFF/U453  ( .A(\UART_TXFF/iFIFOMem[43][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1636 ) );
  notech_mux2 \UART_TXFF/U452  ( .A(\UART_TXFF/iFIFOMem[43][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1637 ) );
  notech_mux2 \UART_TXFF/U451  ( .A(\UART_TXFF/iFIFOMem[43][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1638 ) );
  notech_mux2 \UART_TXFF/U450  ( .A(\UART_TXFF/iFIFOMem[43][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1639 ) );
  notech_mux2 \UART_TXFF/U449  ( .A(\UART_TXFF/iFIFOMem[43][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1640 ) );
  notech_mux2 \UART_TXFF/U448  ( .A(\UART_TXFF/iFIFOMem[43][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1641 ) );
  notech_mux2 \UART_TXFF/U447  ( .A(\UART_TXFF/iFIFOMem[43][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1642 ) );
  notech_mux2 \UART_TXFF/U446  ( .A(\UART_TXFF/iFIFOMem[43][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n274 ), .Z(\UART_TXFF/n1643 ) );
  notech_and2 \UART_TXFF/U445  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n273 ) );
  notech_mux2 \UART_TXFF/U444  ( .A(\UART_TXFF/iFIFOMem[44][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1644 ) );
  notech_mux2 \UART_TXFF/U443  ( .A(\UART_TXFF/iFIFOMem[44][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1645 ) );
  notech_mux2 \UART_TXFF/U442  ( .A(\UART_TXFF/iFIFOMem[44][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1646 ) );
  notech_mux2 \UART_TXFF/U441  ( .A(\UART_TXFF/iFIFOMem[44][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1647 ) );
  notech_mux2 \UART_TXFF/U440  ( .A(\UART_TXFF/iFIFOMem[44][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1648 ) );
  notech_mux2 \UART_TXFF/U439  ( .A(\UART_TXFF/iFIFOMem[44][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1649 ) );
  notech_mux2 \UART_TXFF/U438  ( .A(\UART_TXFF/iFIFOMem[44][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1650 ) );
  notech_mux2 \UART_TXFF/U437  ( .A(\UART_TXFF/iFIFOMem[44][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n273 ), .Z(\UART_TXFF/n1651 ) );
  notech_and2 \UART_TXFF/U436  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n272 ) );
  notech_mux2 \UART_TXFF/U435  ( .A(\UART_TXFF/iFIFOMem[45][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1652 ) );
  notech_mux2 \UART_TXFF/U434  ( .A(\UART_TXFF/iFIFOMem[45][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1653 ) );
  notech_mux2 \UART_TXFF/U433  ( .A(\UART_TXFF/iFIFOMem[45][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1654 ) );
  notech_mux2 \UART_TXFF/U432  ( .A(\UART_TXFF/iFIFOMem[45][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1655 ) );
  notech_mux2 \UART_TXFF/U431  ( .A(\UART_TXFF/iFIFOMem[45][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1656 ) );
  notech_mux2 \UART_TXFF/U430  ( .A(\UART_TXFF/iFIFOMem[45][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1657 ) );
  notech_mux2 \UART_TXFF/U429  ( .A(\UART_TXFF/iFIFOMem[45][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1658 ) );
  notech_mux2 \UART_TXFF/U428  ( .A(\UART_TXFF/iFIFOMem[45][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n272 ), .Z(\UART_TXFF/n1659 ) );
  notech_and2 \UART_TXFF/U427  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n271 ) );
  notech_mux2 \UART_TXFF/U426  ( .A(\UART_TXFF/iFIFOMem[46][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1660 ) );
  notech_mux2 \UART_TXFF/U425  ( .A(\UART_TXFF/iFIFOMem[46][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1661 ) );
  notech_mux2 \UART_TXFF/U424  ( .A(\UART_TXFF/iFIFOMem[46][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1662 ) );
  notech_mux2 \UART_TXFF/U423  ( .A(\UART_TXFF/iFIFOMem[46][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1663 ) );
  notech_mux2 \UART_TXFF/U422  ( .A(\UART_TXFF/iFIFOMem[46][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1664 ) );
  notech_mux2 \UART_TXFF/U421  ( .A(\UART_TXFF/iFIFOMem[46][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1665 ) );
  notech_mux2 \UART_TXFF/U420  ( .A(\UART_TXFF/iFIFOMem[46][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1666 ) );
  notech_mux2 \UART_TXFF/U419  ( .A(\UART_TXFF/iFIFOMem[46][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n271 ), .Z(\UART_TXFF/n1667 ) );
  notech_and2 \UART_TXFF/U418  ( .A(\UART_TXFF/n270 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n269 ) );
  notech_mux2 \UART_TXFF/U417  ( .A(\UART_TXFF/iFIFOMem[47][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1668 ) );
  notech_mux2 \UART_TXFF/U416  ( .A(\UART_TXFF/iFIFOMem[47][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1669 ) );
  notech_mux2 \UART_TXFF/U415  ( .A(\UART_TXFF/iFIFOMem[47][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1670 ) );
  notech_mux2 \UART_TXFF/U414  ( .A(\UART_TXFF/iFIFOMem[47][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1671 ) );
  notech_mux2 \UART_TXFF/U413  ( .A(\UART_TXFF/iFIFOMem[47][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1672 ) );
  notech_mux2 \UART_TXFF/U412  ( .A(\UART_TXFF/iFIFOMem[47][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1673 ) );
  notech_mux2 \UART_TXFF/U411  ( .A(\UART_TXFF/iFIFOMem[47][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1674 ) );
  notech_mux2 \UART_TXFF/U410  ( .A(\UART_TXFF/iFIFOMem[47][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n269 ), .Z(\UART_TXFF/n1675 ) );
  notech_ao3 \UART_TXFF/U409  ( .A(\UART_TXFF/iWRAddr[4] ), .B(
        \UART_TXFF/n259 ), .C(\UART_TXFF/iWRAddr[3] ), .Z(\UART_TXFF/n261 ) );
  notech_and2 \UART_TXFF/U408  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n268 ) );
  notech_mux2 \UART_TXFF/U407  ( .A(\UART_TXFF/iFIFOMem[48][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1676 ) );
  notech_mux2 \UART_TXFF/U406  ( .A(\UART_TXFF/iFIFOMem[48][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1677 ) );
  notech_mux2 \UART_TXFF/U405  ( .A(\UART_TXFF/iFIFOMem[48][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1678 ) );
  notech_mux2 \UART_TXFF/U404  ( .A(\UART_TXFF/iFIFOMem[48][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1679 ) );
  notech_mux2 \UART_TXFF/U403  ( .A(\UART_TXFF/iFIFOMem[48][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1680 ) );
  notech_mux2 \UART_TXFF/U402  ( .A(\UART_TXFF/iFIFOMem[48][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1681 ) );
  notech_mux2 \UART_TXFF/U401  ( .A(\UART_TXFF/iFIFOMem[48][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1682 ) );
  notech_mux2 \UART_TXFF/U400  ( .A(\UART_TXFF/iFIFOMem[48][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n268 ), .Z(\UART_TXFF/n1683 ) );
  notech_and2 \UART_TXFF/U399  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n267 ) );
  notech_mux2 \UART_TXFF/U398  ( .A(\UART_TXFF/iFIFOMem[49][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1684 ) );
  notech_mux2 \UART_TXFF/U397  ( .A(\UART_TXFF/iFIFOMem[49][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1685 ) );
  notech_mux2 \UART_TXFF/U396  ( .A(\UART_TXFF/iFIFOMem[49][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1686 ) );
  notech_mux2 \UART_TXFF/U395  ( .A(\UART_TXFF/iFIFOMem[49][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1687 ) );
  notech_mux2 \UART_TXFF/U394  ( .A(\UART_TXFF/iFIFOMem[49][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1688 ) );
  notech_mux2 \UART_TXFF/U393  ( .A(\UART_TXFF/iFIFOMem[49][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1689 ) );
  notech_mux2 \UART_TXFF/U392  ( .A(\UART_TXFF/iFIFOMem[49][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1690 ) );
  notech_mux2 \UART_TXFF/U391  ( .A(\UART_TXFF/iFIFOMem[49][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n267 ), .Z(\UART_TXFF/n1691 ) );
  notech_and2 \UART_TXFF/U390  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n266 ) );
  notech_mux2 \UART_TXFF/U389  ( .A(\UART_TXFF/iFIFOMem[50][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1692 ) );
  notech_mux2 \UART_TXFF/U388  ( .A(\UART_TXFF/iFIFOMem[50][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1693 ) );
  notech_mux2 \UART_TXFF/U387  ( .A(\UART_TXFF/iFIFOMem[50][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1694 ) );
  notech_mux2 \UART_TXFF/U386  ( .A(\UART_TXFF/iFIFOMem[50][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1695 ) );
  notech_mux2 \UART_TXFF/U385  ( .A(\UART_TXFF/iFIFOMem[50][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1696 ) );
  notech_mux2 \UART_TXFF/U384  ( .A(\UART_TXFF/iFIFOMem[50][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1697 ) );
  notech_mux2 \UART_TXFF/U383  ( .A(\UART_TXFF/iFIFOMem[50][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1698 ) );
  notech_mux2 \UART_TXFF/U382  ( .A(\UART_TXFF/iFIFOMem[50][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n266 ), .Z(\UART_TXFF/n1699 ) );
  notech_and2 \UART_TXFF/U381  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n265 ) );
  notech_mux2 \UART_TXFF/U380  ( .A(\UART_TXFF/iFIFOMem[51][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1700 ) );
  notech_mux2 \UART_TXFF/U379  ( .A(\UART_TXFF/iFIFOMem[51][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1701 ) );
  notech_mux2 \UART_TXFF/U378  ( .A(\UART_TXFF/iFIFOMem[51][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1702 ) );
  notech_mux2 \UART_TXFF/U377  ( .A(\UART_TXFF/iFIFOMem[51][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1703 ) );
  notech_mux2 \UART_TXFF/U376  ( .A(\UART_TXFF/iFIFOMem[51][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1704 ) );
  notech_mux2 \UART_TXFF/U375  ( .A(\UART_TXFF/iFIFOMem[51][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1705 ) );
  notech_mux2 \UART_TXFF/U374  ( .A(\UART_TXFF/iFIFOMem[51][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1706 ) );
  notech_mux2 \UART_TXFF/U373  ( .A(\UART_TXFF/iFIFOMem[51][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n265 ), .Z(\UART_TXFF/n1707 ) );
  notech_and2 \UART_TXFF/U372  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n264 ) );
  notech_mux2 \UART_TXFF/U371  ( .A(\UART_TXFF/iFIFOMem[52][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1708 ) );
  notech_mux2 \UART_TXFF/U370  ( .A(\UART_TXFF/iFIFOMem[52][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1709 ) );
  notech_mux2 \UART_TXFF/U369  ( .A(\UART_TXFF/iFIFOMem[52][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1710 ) );
  notech_mux2 \UART_TXFF/U368  ( .A(\UART_TXFF/iFIFOMem[52][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1711 ) );
  notech_mux2 \UART_TXFF/U367  ( .A(\UART_TXFF/iFIFOMem[52][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1712 ) );
  notech_mux2 \UART_TXFF/U366  ( .A(\UART_TXFF/iFIFOMem[52][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1713 ) );
  notech_mux2 \UART_TXFF/U365  ( .A(\UART_TXFF/iFIFOMem[52][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1714 ) );
  notech_mux2 \UART_TXFF/U364  ( .A(\UART_TXFF/iFIFOMem[52][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n264 ), .Z(\UART_TXFF/n1715 ) );
  notech_and2 \UART_TXFF/U363  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n263 ) );
  notech_mux2 \UART_TXFF/U362  ( .A(\UART_TXFF/iFIFOMem[53][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1716 ) );
  notech_mux2 \UART_TXFF/U361  ( .A(\UART_TXFF/iFIFOMem[53][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1717 ) );
  notech_mux2 \UART_TXFF/U360  ( .A(\UART_TXFF/iFIFOMem[53][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1718 ) );
  notech_mux2 \UART_TXFF/U359  ( .A(\UART_TXFF/iFIFOMem[53][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1719 ) );
  notech_mux2 \UART_TXFF/U358  ( .A(\UART_TXFF/iFIFOMem[53][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1720 ) );
  notech_mux2 \UART_TXFF/U357  ( .A(\UART_TXFF/iFIFOMem[53][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1721 ) );
  notech_mux2 \UART_TXFF/U356  ( .A(\UART_TXFF/iFIFOMem[53][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1722 ) );
  notech_mux2 \UART_TXFF/U355  ( .A(\UART_TXFF/iFIFOMem[53][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n263 ), .Z(\UART_TXFF/n1723 ) );
  notech_and2 \UART_TXFF/U354  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n262 ) );
  notech_mux2 \UART_TXFF/U353  ( .A(\UART_TXFF/iFIFOMem[54][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1724 ) );
  notech_mux2 \UART_TXFF/U352  ( .A(\UART_TXFF/iFIFOMem[54][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1725 ) );
  notech_mux2 \UART_TXFF/U351  ( .A(\UART_TXFF/iFIFOMem[54][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1726 ) );
  notech_mux2 \UART_TXFF/U350  ( .A(\UART_TXFF/iFIFOMem[54][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1727 ) );
  notech_mux2 \UART_TXFF/U349  ( .A(\UART_TXFF/iFIFOMem[54][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1728 ) );
  notech_mux2 \UART_TXFF/U348  ( .A(\UART_TXFF/iFIFOMem[54][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1729 ) );
  notech_mux2 \UART_TXFF/U347  ( .A(\UART_TXFF/iFIFOMem[54][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1730 ) );
  notech_mux2 \UART_TXFF/U346  ( .A(\UART_TXFF/iFIFOMem[54][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n262 ), .Z(\UART_TXFF/n1731 ) );
  notech_and2 \UART_TXFF/U345  ( .A(\UART_TXFF/n261 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n260 ) );
  notech_mux2 \UART_TXFF/U344  ( .A(\UART_TXFF/iFIFOMem[55][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1732 ) );
  notech_mux2 \UART_TXFF/U343  ( .A(\UART_TXFF/iFIFOMem[55][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1733 ) );
  notech_mux2 \UART_TXFF/U342  ( .A(\UART_TXFF/iFIFOMem[55][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1734 ) );
  notech_mux2 \UART_TXFF/U341  ( .A(\UART_TXFF/iFIFOMem[55][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1735 ) );
  notech_mux2 \UART_TXFF/U340  ( .A(\UART_TXFF/iFIFOMem[55][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1736 ) );
  notech_mux2 \UART_TXFF/U339  ( .A(\UART_TXFF/iFIFOMem[55][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1737 ) );
  notech_mux2 \UART_TXFF/U338  ( .A(\UART_TXFF/iFIFOMem[55][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1738 ) );
  notech_mux2 \UART_TXFF/U337  ( .A(\UART_TXFF/iFIFOMem[55][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n260 ), .Z(\UART_TXFF/n1739 ) );
  notech_and3 \UART_TXFF/U336  ( .A(\UART_TXFF/iWRAddr[4] ), .B(
        \UART_TXFF/n259 ), .C(\UART_TXFF/iWRAddr[3] ), .Z(\UART_TXFF/n243 ) );
  notech_and2 \UART_TXFF/U335  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n258 ), 
        .Z(\UART_TXFF/n257 ) );
  notech_mux2 \UART_TXFF/U334  ( .A(\UART_TXFF/iFIFOMem[56][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1740 ) );
  notech_mux2 \UART_TXFF/U333  ( .A(\UART_TXFF/iFIFOMem[56][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1741 ) );
  notech_mux2 \UART_TXFF/U332  ( .A(\UART_TXFF/iFIFOMem[56][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1742 ) );
  notech_mux2 \UART_TXFF/U331  ( .A(\UART_TXFF/iFIFOMem[56][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1743 ) );
  notech_mux2 \UART_TXFF/U330  ( .A(\UART_TXFF/iFIFOMem[56][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1744 ) );
  notech_mux2 \UART_TXFF/U329  ( .A(\UART_TXFF/iFIFOMem[56][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1745 ) );
  notech_mux2 \UART_TXFF/U328  ( .A(\UART_TXFF/iFIFOMem[56][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1746 ) );
  notech_mux2 \UART_TXFF/U327  ( .A(\UART_TXFF/iFIFOMem[56][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n257 ), .Z(\UART_TXFF/n1747 ) );
  notech_and2 \UART_TXFF/U326  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n256 ), 
        .Z(\UART_TXFF/n255 ) );
  notech_mux2 \UART_TXFF/U325  ( .A(\UART_TXFF/iFIFOMem[57][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1748 ) );
  notech_mux2 \UART_TXFF/U324  ( .A(\UART_TXFF/iFIFOMem[57][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1749 ) );
  notech_mux2 \UART_TXFF/U323  ( .A(\UART_TXFF/iFIFOMem[57][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1750 ) );
  notech_mux2 \UART_TXFF/U322  ( .A(\UART_TXFF/iFIFOMem[57][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1751 ) );
  notech_mux2 \UART_TXFF/U321  ( .A(\UART_TXFF/iFIFOMem[57][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1752 ) );
  notech_mux2 \UART_TXFF/U320  ( .A(\UART_TXFF/iFIFOMem[57][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1753 ) );
  notech_mux2 \UART_TXFF/U319  ( .A(\UART_TXFF/iFIFOMem[57][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1754 ) );
  notech_mux2 \UART_TXFF/U318  ( .A(\UART_TXFF/iFIFOMem[57][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n255 ), .Z(\UART_TXFF/n1755 ) );
  notech_and2 \UART_TXFF/U317  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n254 ), 
        .Z(\UART_TXFF/n253 ) );
  notech_mux2 \UART_TXFF/U316  ( .A(\UART_TXFF/iFIFOMem[58][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1756 ) );
  notech_mux2 \UART_TXFF/U315  ( .A(\UART_TXFF/iFIFOMem[58][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1757 ) );
  notech_mux2 \UART_TXFF/U314  ( .A(\UART_TXFF/iFIFOMem[58][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1758 ) );
  notech_mux2 \UART_TXFF/U313  ( .A(\UART_TXFF/iFIFOMem[58][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1759 ) );
  notech_mux2 \UART_TXFF/U312  ( .A(\UART_TXFF/iFIFOMem[58][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1760 ) );
  notech_mux2 \UART_TXFF/U311  ( .A(\UART_TXFF/iFIFOMem[58][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1761 ) );
  notech_mux2 \UART_TXFF/U310  ( .A(\UART_TXFF/iFIFOMem[58][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1762 ) );
  notech_mux2 \UART_TXFF/U309  ( .A(\UART_TXFF/iFIFOMem[58][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n253 ), .Z(\UART_TXFF/n1763 ) );
  notech_and2 \UART_TXFF/U308  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n252 ), 
        .Z(\UART_TXFF/n251 ) );
  notech_mux2 \UART_TXFF/U307  ( .A(\UART_TXFF/iFIFOMem[59][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1764 ) );
  notech_mux2 \UART_TXFF/U306  ( .A(\UART_TXFF/iFIFOMem[59][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1765 ) );
  notech_mux2 \UART_TXFF/U305  ( .A(\UART_TXFF/iFIFOMem[59][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1766 ) );
  notech_mux2 \UART_TXFF/U304  ( .A(\UART_TXFF/iFIFOMem[59][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1767 ) );
  notech_mux2 \UART_TXFF/U303  ( .A(\UART_TXFF/iFIFOMem[59][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1768 ) );
  notech_mux2 \UART_TXFF/U302  ( .A(\UART_TXFF/iFIFOMem[59][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1769 ) );
  notech_mux2 \UART_TXFF/U301  ( .A(\UART_TXFF/iFIFOMem[59][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1770 ) );
  notech_mux2 \UART_TXFF/U300  ( .A(\UART_TXFF/iFIFOMem[59][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n251 ), .Z(\UART_TXFF/n1771 ) );
  notech_and2 \UART_TXFF/U299  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n250 ), 
        .Z(\UART_TXFF/n249 ) );
  notech_mux2 \UART_TXFF/U298  ( .A(\UART_TXFF/iFIFOMem[60][0] ), .B(iDIN[0]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1772 ) );
  notech_mux2 \UART_TXFF/U297  ( .A(\UART_TXFF/iFIFOMem[60][1] ), .B(iDIN[1]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1773 ) );
  notech_mux2 \UART_TXFF/U296  ( .A(\UART_TXFF/iFIFOMem[60][2] ), .B(iDIN[2]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1774 ) );
  notech_mux2 \UART_TXFF/U295  ( .A(\UART_TXFF/iFIFOMem[60][3] ), .B(iDIN[3]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1775 ) );
  notech_mux2 \UART_TXFF/U294  ( .A(\UART_TXFF/iFIFOMem[60][4] ), .B(iDIN[4]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1776 ) );
  notech_mux2 \UART_TXFF/U293  ( .A(\UART_TXFF/iFIFOMem[60][5] ), .B(iDIN[5]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1777 ) );
  notech_mux2 \UART_TXFF/U292  ( .A(\UART_TXFF/iFIFOMem[60][6] ), .B(iDIN[6]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1778 ) );
  notech_mux2 \UART_TXFF/U291  ( .A(\UART_TXFF/iFIFOMem[60][7] ), .B(iDIN[7]), 
        .S(\UART_TXFF/n249 ), .Z(\UART_TXFF/n1779 ) );
  notech_and2 \UART_TXFF/U290  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n248 ), 
        .Z(\UART_TXFF/n247 ) );
  notech_mux2 \UART_TXFF/U289  ( .A(\UART_TXFF/iFIFOMem[61][0] ), .B(
        \UART_TXFF/n4 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1780 ) );
  notech_mux2 \UART_TXFF/U288  ( .A(\UART_TXFF/iFIFOMem[61][1] ), .B(
        \UART_TXFF/n8 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1781 ) );
  notech_mux2 \UART_TXFF/U287  ( .A(\UART_TXFF/iFIFOMem[61][2] ), .B(
        \UART_TXFF/n12 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1782 ) );
  notech_mux2 \UART_TXFF/U286  ( .A(\UART_TXFF/iFIFOMem[61][3] ), .B(
        \UART_TXFF/n16 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1783 ) );
  notech_mux2 \UART_TXFF/U285  ( .A(\UART_TXFF/iFIFOMem[61][4] ), .B(
        \UART_TXFF/n20 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1784 ) );
  notech_mux2 \UART_TXFF/U284  ( .A(\UART_TXFF/iFIFOMem[61][5] ), .B(
        \UART_TXFF/n24 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1785 ) );
  notech_mux2 \UART_TXFF/U283  ( .A(\UART_TXFF/iFIFOMem[61][6] ), .B(
        \UART_TXFF/n28 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1786 ) );
  notech_mux2 \UART_TXFF/U282  ( .A(\UART_TXFF/iFIFOMem[61][7] ), .B(
        \UART_TXFF/n32 ), .S(\UART_TXFF/n247 ), .Z(\UART_TXFF/n1787 ) );
  notech_and2 \UART_TXFF/U281  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n246 ), 
        .Z(\UART_TXFF/n245 ) );
  notech_mux2 \UART_TXFF/U280  ( .A(\UART_TXFF/iFIFOMem[62][0] ), .B(
        \UART_TXFF/n3 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1788 ) );
  notech_mux2 \UART_TXFF/U279  ( .A(\UART_TXFF/iFIFOMem[62][1] ), .B(
        \UART_TXFF/n7 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1789 ) );
  notech_mux2 \UART_TXFF/U278  ( .A(\UART_TXFF/iFIFOMem[62][2] ), .B(
        \UART_TXFF/n11 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1790 ) );
  notech_mux2 \UART_TXFF/U277  ( .A(\UART_TXFF/iFIFOMem[62][3] ), .B(
        \UART_TXFF/n15 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1791 ) );
  notech_mux2 \UART_TXFF/U276  ( .A(\UART_TXFF/iFIFOMem[62][4] ), .B(
        \UART_TXFF/n19 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1792 ) );
  notech_mux2 \UART_TXFF/U275  ( .A(\UART_TXFF/iFIFOMem[62][5] ), .B(
        \UART_TXFF/n23 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1793 ) );
  notech_mux2 \UART_TXFF/U274  ( .A(\UART_TXFF/iFIFOMem[62][6] ), .B(
        \UART_TXFF/n27 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1794 ) );
  notech_mux2 \UART_TXFF/U273  ( .A(\UART_TXFF/iFIFOMem[62][7] ), .B(
        \UART_TXFF/n31 ), .S(\UART_TXFF/n245 ), .Z(\UART_TXFF/n1795 ) );
  notech_and2 \UART_TXFF/U272  ( .A(\UART_TXFF/n243 ), .B(\UART_TXFF/n244 ), 
        .Z(\UART_TXFF/n242 ) );
  notech_mux2 \UART_TXFF/U271  ( .A(\UART_TXFF/iFIFOMem[63][0] ), .B(
        \UART_TXFF/n2 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1796 ) );
  notech_mux2 \UART_TXFF/U270  ( .A(\UART_TXFF/iFIFOMem[63][1] ), .B(
        \UART_TXFF/n6 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1797 ) );
  notech_mux2 \UART_TXFF/U269  ( .A(\UART_TXFF/iFIFOMem[63][2] ), .B(
        \UART_TXFF/n10 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1798 ) );
  notech_mux2 \UART_TXFF/U268  ( .A(\UART_TXFF/iFIFOMem[63][3] ), .B(
        \UART_TXFF/n14 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1799 ) );
  notech_mux2 \UART_TXFF/U267  ( .A(\UART_TXFF/iFIFOMem[63][4] ), .B(
        \UART_TXFF/n18 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1800 ) );
  notech_mux2 \UART_TXFF/U266  ( .A(\UART_TXFF/iFIFOMem[63][5] ), .B(
        \UART_TXFF/n22 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1801 ) );
  notech_mux2 \UART_TXFF/U265  ( .A(\UART_TXFF/iFIFOMem[63][6] ), .B(
        \UART_TXFF/n26 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1802 ) );
  notech_mux2 \UART_TXFF/U264  ( .A(\UART_TXFF/iFIFOMem[63][7] ), .B(
        \UART_TXFF/n30 ), .S(\UART_TXFF/n242 ), .Z(\UART_TXFF/n1803 ) );
  notech_and2 \UART_TXFF/U263  ( .A(iTXFIFORead), .B(n520), .Z(
        \UART_TXFF/n240 ) );
  notech_or2 \UART_TXFF/U262  ( .A(\UART_TXFF/n240 ), .B(iFCR[2]), .Z(
        \UART_TXFF/n212 ) );
  notech_inv \UART_TXFF/U261  ( .A(\UART_TXFF/N17 ), .Z(\UART_TXFF/n238 ) );
  notech_nand2 \UART_TXFF/U260  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n228 ), 
        .Z(\UART_TXFF/n211 ) );
  notech_inv \UART_TXFF/U259  ( .A(\UART_TXFF/N37 ), .Z(\UART_TXFF/n239 ) );
  notech_nao4 \UART_TXFF/U258  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n238 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n239 ), .Z(\UART_TXFF/n1804 ) );
  notech_inv \UART_TXFF/U257  ( .A(\UART_TXFF/N36 ), .Z(\UART_TXFF/n237 ) );
  notech_nao4 \UART_TXFF/U256  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n236 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n237 ), .Z(\UART_TXFF/n1805 ) );
  notech_inv \UART_TXFF/U255  ( .A(\UART_TXFF/N35 ), .Z(\UART_TXFF/n235 ) );
  notech_nao4 \UART_TXFF/U254  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n234 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n235 ), .Z(\UART_TXFF/n1806 ) );
  notech_inv \UART_TXFF/U253  ( .A(\UART_TXFF/N34 ), .Z(\UART_TXFF/n233 ) );
  notech_nao4 \UART_TXFF/U252  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n232 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n233 ), .Z(\UART_TXFF/n1807 ) );
  notech_inv \UART_TXFF/U251  ( .A(\UART_TXFF/N33 ), .Z(\UART_TXFF/n231 ) );
  notech_nao4 \UART_TXFF/U250  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n42 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n231 ), .Z(\UART_TXFF/n1808 ) );
  notech_inv \UART_TXFF/U249  ( .A(\UART_TXFF/iRDAddr[6] ), .Z(
        \UART_TXFF/n229 ) );
  notech_inv \UART_TXFF/U248  ( .A(\UART_TXFF/N38 ), .Z(\UART_TXFF/n230 ) );
  notech_nao4 \UART_TXFF/U247  ( .A(\UART_TXFF/n212 ), .B(\UART_TXFF/n229 ), 
        .C(\UART_TXFF/n211 ), .D(\UART_TXFF/n230 ), .Z(\UART_TXFF/n1809 ) );
  notech_inv \UART_TXFF/U246  ( .A(\UART_TXFF/iWRAddr[5] ), .Z(
        \UART_TXFF/n226 ) );
  notech_nand2 \UART_TXFF/U245  ( .A(\UART_TXFF/n214 ), .B(\UART_TXFF/n228 ), 
        .Z(\UART_TXFF/n215 ) );
  notech_inv \UART_TXFF/U244  ( .A(\UART_TXFF/N29 ), .Z(\UART_TXFF/n227 ) );
  notech_nao4 \UART_TXFF/U243  ( .A(\UART_TXFF/n226 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n227 ), .Z(\UART_TXFF/n1810 ) );
  notech_inv \UART_TXFF/U242  ( .A(\UART_TXFF/iWRAddr[4] ), .Z(
        \UART_TXFF/n224 ) );
  notech_inv \UART_TXFF/U241  ( .A(\UART_TXFF/N28 ), .Z(\UART_TXFF/n225 ) );
  notech_nao4 \UART_TXFF/U240  ( .A(\UART_TXFF/n224 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n225 ), .Z(\UART_TXFF/n1811 ) );
  notech_inv \UART_TXFF/U239  ( .A(\UART_TXFF/N27 ), .Z(\UART_TXFF/n223 ) );
  notech_nao4 \UART_TXFF/U238  ( .A(\UART_TXFF/n222 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n223 ), .Z(\UART_TXFF/n1812 ) );
  notech_inv \UART_TXFF/U237  ( .A(\UART_TXFF/N26 ), .Z(\UART_TXFF/n221 ) );
  notech_nao4 \UART_TXFF/U236  ( .A(\UART_TXFF/n220 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n221 ), .Z(\UART_TXFF/n1813 ) );
  notech_inv \UART_TXFF/U235  ( .A(\UART_TXFF/N25 ), .Z(\UART_TXFF/n219 ) );
  notech_nao4 \UART_TXFF/U234  ( .A(\UART_TXFF/n218 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n219 ), .Z(\UART_TXFF/n1814 ) );
  notech_mux2 \UART_TXFF/U233  ( .A(\UART_TXFF/n215 ), .B(\UART_TXFF/n214 ), 
        .S(\UART_TXFF/iWRAddr[0] ), .Z(\UART_TXFF/n217 ) );
  notech_inv \UART_TXFF/U232  ( .A(\UART_TXFF/n217 ), .Z(\UART_TXFF/n1815 ) );
  notech_inv \UART_TXFF/U231  ( .A(\UART_TXFF/N30 ), .Z(\UART_TXFF/n216 ) );
  notech_nao4 \UART_TXFF/U230  ( .A(\UART_TXFF/n213 ), .B(\UART_TXFF/n214 ), 
        .C(\UART_TXFF/n215 ), .D(\UART_TXFF/n216 ), .Z(\UART_TXFF/n1816 ) );
  notech_mux2 \UART_TXFF/U229  ( .A(\UART_TXFF/n211 ), .B(\UART_TXFF/n212 ), 
        .S(\UART_TXFF/N12 ), .Z(\UART_TXFF/n210 ) );
  notech_inv \UART_TXFF/U228  ( .A(\UART_TXFF/n210 ), .Z(\UART_TXFF/n1817 ) );
  notech_mux2 \UART_TXFF/U227  ( .A(\UART_TXFF/N130 ), .B(iTXFIFOQ[0]), .S(RST), .Z(\UART_TXFF/n758 ) );
  notech_mux2 \UART_TXFF/U226  ( .A(\UART_TXFF/N129 ), .B(iTXFIFOQ[1]), .S(RST), .Z(\UART_TXFF/n760 ) );
  notech_mux2 \UART_TXFF/U225  ( .A(\UART_TXFF/N128 ), .B(iTXFIFOQ[2]), .S(RST), .Z(\UART_TXFF/n762 ) );
  notech_mux2 \UART_TXFF/U224  ( .A(\UART_TXFF/N127 ), .B(iTXFIFOQ[3]), .S(RST), .Z(\UART_TXFF/n764 ) );
  notech_mux2 \UART_TXFF/U223  ( .A(\UART_TXFF/N126 ), .B(iTXFIFOQ[4]), .S(RST), .Z(\UART_TXFF/n766 ) );
  notech_mux2 \UART_TXFF/U222  ( .A(\UART_TXFF/N125 ), .B(iTXFIFOQ[5]), .S(RST), .Z(\UART_TXFF/n768 ) );
  notech_mux2 \UART_TXFF/U221  ( .A(\UART_TXFF/N124 ), .B(iTXFIFOQ[6]), .S(RST), .Z(\UART_TXFF/n770 ) );
  notech_mux2 \UART_TXFF/U220  ( .A(\UART_TXFF/N123 ), .B(iTXFIFOQ[7]), .S(RST), .Z(\UART_TXFF/n772 ) );
  notech_mux4 \UART_TXFF/U219  ( .A(\UART_TXFF/n209 ), .B(\UART_TXFF/n199 ), 
        .C(\UART_TXFF/n204 ), .D(\UART_TXFF/n194 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N123 ) );
  notech_mux4 \UART_TXFF/U218  ( .A(\UART_TXFF/n208 ), .B(\UART_TXFF/n206 ), 
        .C(\UART_TXFF/n207 ), .D(\UART_TXFF/n205 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n209 ) );
  notech_mux4 \UART_TXFF/U217  ( .A(\UART_TXFF/iFIFOMem[0][7] ), .B(
        \UART_TXFF/iFIFOMem[2][7] ), .C(\UART_TXFF/iFIFOMem[1][7] ), .D(
        \UART_TXFF/iFIFOMem[3][7] ), .S0(\UART_TXFF/N13 ), .S1(\UART_TXFF/N12 ), .Z(\UART_TXFF/n208 ) );
  notech_mux4 \UART_TXFF/U216  ( .A(\UART_TXFF/iFIFOMem[4][7] ), .B(
        \UART_TXFF/iFIFOMem[6][7] ), .C(\UART_TXFF/iFIFOMem[5][7] ), .D(
        \UART_TXFF/iFIFOMem[7][7] ), .S0(\UART_TXFF/N13 ), .S1(\UART_TXFF/N12 ), .Z(\UART_TXFF/n207 ) );
  notech_mux4 \UART_TXFF/U215  ( .A(\UART_TXFF/iFIFOMem[8][7] ), .B(
        \UART_TXFF/iFIFOMem[10][7] ), .C(\UART_TXFF/iFIFOMem[9][7] ), .D(
        \UART_TXFF/iFIFOMem[11][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n206 ) );
  notech_mux4 \UART_TXFF/U214  ( .A(\UART_TXFF/iFIFOMem[12][7] ), .B(
        \UART_TXFF/iFIFOMem[14][7] ), .C(\UART_TXFF/iFIFOMem[13][7] ), .D(
        \UART_TXFF/iFIFOMem[15][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n205 ) );
  notech_mux4 \UART_TXFF/U213  ( .A(\UART_TXFF/n203 ), .B(\UART_TXFF/n201 ), 
        .C(\UART_TXFF/n202 ), .D(\UART_TXFF/n200 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n204 ) );
  notech_mux4 \UART_TXFF/U212  ( .A(\UART_TXFF/iFIFOMem[16][7] ), .B(
        \UART_TXFF/iFIFOMem[18][7] ), .C(\UART_TXFF/iFIFOMem[17][7] ), .D(
        \UART_TXFF/iFIFOMem[19][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n203 ) );
  notech_mux4 \UART_TXFF/U211  ( .A(\UART_TXFF/iFIFOMem[20][7] ), .B(
        \UART_TXFF/iFIFOMem[22][7] ), .C(\UART_TXFF/iFIFOMem[21][7] ), .D(
        \UART_TXFF/iFIFOMem[23][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n202 ) );
  notech_mux4 \UART_TXFF/U210  ( .A(\UART_TXFF/iFIFOMem[24][7] ), .B(
        \UART_TXFF/iFIFOMem[26][7] ), .C(\UART_TXFF/iFIFOMem[25][7] ), .D(
        \UART_TXFF/iFIFOMem[27][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n201 ) );
  notech_mux4 \UART_TXFF/U209  ( .A(\UART_TXFF/iFIFOMem[28][7] ), .B(
        \UART_TXFF/iFIFOMem[30][7] ), .C(\UART_TXFF/iFIFOMem[29][7] ), .D(
        \UART_TXFF/iFIFOMem[31][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n200 ) );
  notech_mux4 \UART_TXFF/U208  ( .A(\UART_TXFF/n198 ), .B(\UART_TXFF/n196 ), 
        .C(\UART_TXFF/n197 ), .D(\UART_TXFF/n195 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n199 ) );
  notech_mux4 \UART_TXFF/U207  ( .A(\UART_TXFF/iFIFOMem[32][7] ), .B(
        \UART_TXFF/iFIFOMem[34][7] ), .C(\UART_TXFF/iFIFOMem[33][7] ), .D(
        \UART_TXFF/iFIFOMem[35][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n198 ) );
  notech_mux4 \UART_TXFF/U206  ( .A(\UART_TXFF/iFIFOMem[36][7] ), .B(
        \UART_TXFF/iFIFOMem[38][7] ), .C(\UART_TXFF/iFIFOMem[37][7] ), .D(
        \UART_TXFF/iFIFOMem[39][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n197 ) );
  notech_mux4 \UART_TXFF/U205  ( .A(\UART_TXFF/iFIFOMem[40][7] ), .B(
        \UART_TXFF/iFIFOMem[42][7] ), .C(\UART_TXFF/iFIFOMem[41][7] ), .D(
        \UART_TXFF/iFIFOMem[43][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n196 ) );
  notech_mux4 \UART_TXFF/U204  ( .A(\UART_TXFF/iFIFOMem[44][7] ), .B(
        \UART_TXFF/iFIFOMem[46][7] ), .C(\UART_TXFF/iFIFOMem[45][7] ), .D(
        \UART_TXFF/iFIFOMem[47][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n195 ) );
  notech_mux4 \UART_TXFF/U203  ( .A(\UART_TXFF/n193 ), .B(\UART_TXFF/n191 ), 
        .C(\UART_TXFF/n192 ), .D(\UART_TXFF/n190 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n194 ) );
  notech_mux4 \UART_TXFF/U202  ( .A(\UART_TXFF/iFIFOMem[48][7] ), .B(
        \UART_TXFF/iFIFOMem[50][7] ), .C(\UART_TXFF/iFIFOMem[49][7] ), .D(
        \UART_TXFF/iFIFOMem[51][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n193 ) );
  notech_mux4 \UART_TXFF/U201  ( .A(\UART_TXFF/iFIFOMem[52][7] ), .B(
        \UART_TXFF/iFIFOMem[54][7] ), .C(\UART_TXFF/iFIFOMem[53][7] ), .D(
        \UART_TXFF/iFIFOMem[55][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n192 ) );
  notech_mux4 \UART_TXFF/U200  ( .A(\UART_TXFF/iFIFOMem[56][7] ), .B(
        \UART_TXFF/iFIFOMem[58][7] ), .C(\UART_TXFF/iFIFOMem[57][7] ), .D(
        \UART_TXFF/iFIFOMem[59][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n191 ) );
  notech_mux4 \UART_TXFF/U199  ( .A(\UART_TXFF/iFIFOMem[60][7] ), .B(
        \UART_TXFF/iFIFOMem[62][7] ), .C(\UART_TXFF/iFIFOMem[61][7] ), .D(
        \UART_TXFF/iFIFOMem[63][7] ), .S0(\UART_TXFF/N13 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n190 ) );
  notech_mux4 \UART_TXFF/U198  ( .A(\UART_TXFF/n189 ), .B(\UART_TXFF/n179 ), 
        .C(\UART_TXFF/n184 ), .D(\UART_TXFF/n174 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N124 ) );
  notech_mux4 \UART_TXFF/U197  ( .A(\UART_TXFF/n188 ), .B(\UART_TXFF/n186 ), 
        .C(\UART_TXFF/n187 ), .D(\UART_TXFF/n185 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n189 ) );
  notech_mux4 \UART_TXFF/U196  ( .A(\UART_TXFF/iFIFOMem[0][6] ), .B(
        \UART_TXFF/iFIFOMem[2][6] ), .C(\UART_TXFF/iFIFOMem[1][6] ), .D(
        \UART_TXFF/iFIFOMem[3][6] ), .S0(\UART_TXFF/n41 ), .S1(\UART_TXFF/n48 ), .Z(\UART_TXFF/n188 ) );
  notech_mux4 \UART_TXFF/U195  ( .A(\UART_TXFF/iFIFOMem[4][6] ), .B(
        \UART_TXFF/iFIFOMem[6][6] ), .C(\UART_TXFF/iFIFOMem[5][6] ), .D(
        \UART_TXFF/iFIFOMem[7][6] ), .S0(\UART_TXFF/n36 ), .S1(\UART_TXFF/n48 ), .Z(\UART_TXFF/n187 ) );
  notech_mux4 \UART_TXFF/U194  ( .A(\UART_TXFF/iFIFOMem[8][6] ), .B(
        \UART_TXFF/iFIFOMem[10][6] ), .C(\UART_TXFF/iFIFOMem[9][6] ), .D(
        \UART_TXFF/iFIFOMem[11][6] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n186 ) );
  notech_mux4 \UART_TXFF/U193  ( .A(\UART_TXFF/iFIFOMem[12][6] ), .B(
        \UART_TXFF/iFIFOMem[14][6] ), .C(\UART_TXFF/iFIFOMem[13][6] ), .D(
        \UART_TXFF/iFIFOMem[15][6] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n185 ) );
  notech_mux4 \UART_TXFF/U192  ( .A(\UART_TXFF/n183 ), .B(\UART_TXFF/n181 ), 
        .C(\UART_TXFF/n182 ), .D(\UART_TXFF/n180 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n184 ) );
  notech_mux4 \UART_TXFF/U191  ( .A(\UART_TXFF/iFIFOMem[16][6] ), .B(
        \UART_TXFF/iFIFOMem[18][6] ), .C(\UART_TXFF/iFIFOMem[17][6] ), .D(
        \UART_TXFF/iFIFOMem[19][6] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n183 ) );
  notech_mux4 \UART_TXFF/U190  ( .A(\UART_TXFF/iFIFOMem[20][6] ), .B(
        \UART_TXFF/iFIFOMem[22][6] ), .C(\UART_TXFF/iFIFOMem[21][6] ), .D(
        \UART_TXFF/iFIFOMem[23][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n182 ) );
  notech_mux4 \UART_TXFF/U189  ( .A(\UART_TXFF/iFIFOMem[24][6] ), .B(
        \UART_TXFF/iFIFOMem[26][6] ), .C(\UART_TXFF/iFIFOMem[25][6] ), .D(
        \UART_TXFF/iFIFOMem[27][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n181 ) );
  notech_mux4 \UART_TXFF/U188  ( .A(\UART_TXFF/iFIFOMem[28][6] ), .B(
        \UART_TXFF/iFIFOMem[30][6] ), .C(\UART_TXFF/iFIFOMem[29][6] ), .D(
        \UART_TXFF/iFIFOMem[31][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n180 ) );
  notech_mux4 \UART_TXFF/U187  ( .A(\UART_TXFF/n178 ), .B(\UART_TXFF/n176 ), 
        .C(\UART_TXFF/n177 ), .D(\UART_TXFF/n175 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n179 ) );
  notech_mux4 \UART_TXFF/U186  ( .A(\UART_TXFF/iFIFOMem[32][6] ), .B(
        \UART_TXFF/iFIFOMem[34][6] ), .C(\UART_TXFF/iFIFOMem[33][6] ), .D(
        \UART_TXFF/iFIFOMem[35][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n178 ) );
  notech_mux4 \UART_TXFF/U185  ( .A(\UART_TXFF/iFIFOMem[36][6] ), .B(
        \UART_TXFF/iFIFOMem[38][6] ), .C(\UART_TXFF/iFIFOMem[37][6] ), .D(
        \UART_TXFF/iFIFOMem[39][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n177 ) );
  notech_mux4 \UART_TXFF/U184  ( .A(\UART_TXFF/iFIFOMem[40][6] ), .B(
        \UART_TXFF/iFIFOMem[42][6] ), .C(\UART_TXFF/iFIFOMem[41][6] ), .D(
        \UART_TXFF/iFIFOMem[43][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n176 ) );
  notech_mux4 \UART_TXFF/U183  ( .A(\UART_TXFF/iFIFOMem[44][6] ), .B(
        \UART_TXFF/iFIFOMem[46][6] ), .C(\UART_TXFF/iFIFOMem[45][6] ), .D(
        \UART_TXFF/iFIFOMem[47][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n175 ) );
  notech_mux4 \UART_TXFF/U182  ( .A(\UART_TXFF/n173 ), .B(\UART_TXFF/n171 ), 
        .C(\UART_TXFF/n172 ), .D(\UART_TXFF/n170 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n174 ) );
  notech_mux4 \UART_TXFF/U181  ( .A(\UART_TXFF/iFIFOMem[48][6] ), .B(
        \UART_TXFF/iFIFOMem[50][6] ), .C(\UART_TXFF/iFIFOMem[49][6] ), .D(
        \UART_TXFF/iFIFOMem[51][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n173 ) );
  notech_mux4 \UART_TXFF/U180  ( .A(\UART_TXFF/iFIFOMem[52][6] ), .B(
        \UART_TXFF/iFIFOMem[54][6] ), .C(\UART_TXFF/iFIFOMem[53][6] ), .D(
        \UART_TXFF/iFIFOMem[55][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n172 ) );
  notech_mux4 \UART_TXFF/U179  ( .A(\UART_TXFF/iFIFOMem[56][6] ), .B(
        \UART_TXFF/iFIFOMem[58][6] ), .C(\UART_TXFF/iFIFOMem[57][6] ), .D(
        \UART_TXFF/iFIFOMem[59][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n171 ) );
  notech_mux4 \UART_TXFF/U178  ( .A(\UART_TXFF/iFIFOMem[60][6] ), .B(
        \UART_TXFF/iFIFOMem[62][6] ), .C(\UART_TXFF/iFIFOMem[61][6] ), .D(
        \UART_TXFF/iFIFOMem[63][6] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n170 ) );
  notech_mux4 \UART_TXFF/U177  ( .A(\UART_TXFF/n169 ), .B(\UART_TXFF/n159 ), 
        .C(\UART_TXFF/n164 ), .D(\UART_TXFF/n154 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N125 ) );
  notech_mux4 \UART_TXFF/U176  ( .A(\UART_TXFF/n168 ), .B(\UART_TXFF/n166 ), 
        .C(\UART_TXFF/n167 ), .D(\UART_TXFF/n165 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n169 ) );
  notech_mux4 \UART_TXFF/U175  ( .A(\UART_TXFF/iFIFOMem[0][5] ), .B(
        \UART_TXFF/iFIFOMem[2][5] ), .C(\UART_TXFF/iFIFOMem[1][5] ), .D(
        \UART_TXFF/iFIFOMem[3][5] ), .S0(\UART_TXFF/n41 ), .S1(\UART_TXFF/n47 ), .Z(\UART_TXFF/n168 ) );
  notech_mux4 \UART_TXFF/U174  ( .A(\UART_TXFF/iFIFOMem[4][5] ), .B(
        \UART_TXFF/iFIFOMem[6][5] ), .C(\UART_TXFF/iFIFOMem[5][5] ), .D(
        \UART_TXFF/iFIFOMem[7][5] ), .S0(\UART_TXFF/n41 ), .S1(\UART_TXFF/n47 ), .Z(\UART_TXFF/n167 ) );
  notech_mux4 \UART_TXFF/U173  ( .A(\UART_TXFF/iFIFOMem[8][5] ), .B(
        \UART_TXFF/iFIFOMem[10][5] ), .C(\UART_TXFF/iFIFOMem[9][5] ), .D(
        \UART_TXFF/iFIFOMem[11][5] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n166 ) );
  notech_mux4 \UART_TXFF/U172  ( .A(\UART_TXFF/iFIFOMem[12][5] ), .B(
        \UART_TXFF/iFIFOMem[14][5] ), .C(\UART_TXFF/iFIFOMem[13][5] ), .D(
        \UART_TXFF/iFIFOMem[15][5] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n165 ) );
  notech_mux4 \UART_TXFF/U171  ( .A(\UART_TXFF/n163 ), .B(\UART_TXFF/n161 ), 
        .C(\UART_TXFF/n162 ), .D(\UART_TXFF/n160 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n164 ) );
  notech_mux4 \UART_TXFF/U170  ( .A(\UART_TXFF/iFIFOMem[16][5] ), .B(
        \UART_TXFF/iFIFOMem[18][5] ), .C(\UART_TXFF/iFIFOMem[17][5] ), .D(
        \UART_TXFF/iFIFOMem[19][5] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n163 ) );
  notech_mux4 \UART_TXFF/U169  ( .A(\UART_TXFF/iFIFOMem[20][5] ), .B(
        \UART_TXFF/iFIFOMem[22][5] ), .C(\UART_TXFF/iFIFOMem[21][5] ), .D(
        \UART_TXFF/iFIFOMem[23][5] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n162 ) );
  notech_mux4 \UART_TXFF/U168  ( .A(\UART_TXFF/iFIFOMem[24][5] ), .B(
        \UART_TXFF/iFIFOMem[26][5] ), .C(\UART_TXFF/iFIFOMem[25][5] ), .D(
        \UART_TXFF/iFIFOMem[27][5] ), .S0(\UART_TXFF/n41 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n161 ) );
  notech_mux4 \UART_TXFF/U167  ( .A(\UART_TXFF/iFIFOMem[28][5] ), .B(
        \UART_TXFF/iFIFOMem[30][5] ), .C(\UART_TXFF/iFIFOMem[29][5] ), .D(
        \UART_TXFF/iFIFOMem[31][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n160 ) );
  notech_mux4 \UART_TXFF/U166  ( .A(\UART_TXFF/n158 ), .B(\UART_TXFF/n156 ), 
        .C(\UART_TXFF/n157 ), .D(\UART_TXFF/n155 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n159 ) );
  notech_mux4 \UART_TXFF/U165  ( .A(\UART_TXFF/iFIFOMem[32][5] ), .B(
        \UART_TXFF/iFIFOMem[34][5] ), .C(\UART_TXFF/iFIFOMem[33][5] ), .D(
        \UART_TXFF/iFIFOMem[35][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n158 ) );
  notech_mux4 \UART_TXFF/U164  ( .A(\UART_TXFF/iFIFOMem[36][5] ), .B(
        \UART_TXFF/iFIFOMem[38][5] ), .C(\UART_TXFF/iFIFOMem[37][5] ), .D(
        \UART_TXFF/iFIFOMem[39][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n157 ) );
  notech_mux4 \UART_TXFF/U163  ( .A(\UART_TXFF/iFIFOMem[40][5] ), .B(
        \UART_TXFF/iFIFOMem[42][5] ), .C(\UART_TXFF/iFIFOMem[41][5] ), .D(
        \UART_TXFF/iFIFOMem[43][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n156 ) );
  notech_mux4 \UART_TXFF/U162  ( .A(\UART_TXFF/iFIFOMem[44][5] ), .B(
        \UART_TXFF/iFIFOMem[46][5] ), .C(\UART_TXFF/iFIFOMem[45][5] ), .D(
        \UART_TXFF/iFIFOMem[47][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n155 ) );
  notech_mux4 \UART_TXFF/U161  ( .A(\UART_TXFF/n153 ), .B(\UART_TXFF/n151 ), 
        .C(\UART_TXFF/n152 ), .D(\UART_TXFF/n150 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n154 ) );
  notech_mux4 \UART_TXFF/U160  ( .A(\UART_TXFF/iFIFOMem[48][5] ), .B(
        \UART_TXFF/iFIFOMem[50][5] ), .C(\UART_TXFF/iFIFOMem[49][5] ), .D(
        \UART_TXFF/iFIFOMem[51][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n153 ) );
  notech_mux4 \UART_TXFF/U159  ( .A(\UART_TXFF/iFIFOMem[52][5] ), .B(
        \UART_TXFF/iFIFOMem[54][5] ), .C(\UART_TXFF/iFIFOMem[53][5] ), .D(
        \UART_TXFF/iFIFOMem[55][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n152 ) );
  notech_mux4 \UART_TXFF/U158  ( .A(\UART_TXFF/iFIFOMem[56][5] ), .B(
        \UART_TXFF/iFIFOMem[58][5] ), .C(\UART_TXFF/iFIFOMem[57][5] ), .D(
        \UART_TXFF/iFIFOMem[59][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n151 ) );
  notech_mux4 \UART_TXFF/U157  ( .A(\UART_TXFF/iFIFOMem[60][5] ), .B(
        \UART_TXFF/iFIFOMem[62][5] ), .C(\UART_TXFF/iFIFOMem[61][5] ), .D(
        \UART_TXFF/iFIFOMem[63][5] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n150 ) );
  notech_mux4 \UART_TXFF/U156  ( .A(\UART_TXFF/n149 ), .B(\UART_TXFF/n139 ), 
        .C(\UART_TXFF/n144 ), .D(\UART_TXFF/n134 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N126 ) );
  notech_mux4 \UART_TXFF/U155  ( .A(\UART_TXFF/n148 ), .B(\UART_TXFF/n146 ), 
        .C(\UART_TXFF/n147 ), .D(\UART_TXFF/n145 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n149 ) );
  notech_mux4 \UART_TXFF/U154  ( .A(\UART_TXFF/iFIFOMem[0][4] ), .B(
        \UART_TXFF/iFIFOMem[2][4] ), .C(\UART_TXFF/iFIFOMem[1][4] ), .D(
        \UART_TXFF/iFIFOMem[3][4] ), .S0(\UART_TXFF/n40 ), .S1(\UART_TXFF/n46 ), .Z(\UART_TXFF/n148 ) );
  notech_mux4 \UART_TXFF/U153  ( .A(\UART_TXFF/iFIFOMem[4][4] ), .B(
        \UART_TXFF/iFIFOMem[6][4] ), .C(\UART_TXFF/iFIFOMem[5][4] ), .D(
        \UART_TXFF/iFIFOMem[7][4] ), .S0(\UART_TXFF/n40 ), .S1(\UART_TXFF/n46 ), .Z(\UART_TXFF/n147 ) );
  notech_mux4 \UART_TXFF/U152  ( .A(\UART_TXFF/iFIFOMem[8][4] ), .B(
        \UART_TXFF/iFIFOMem[10][4] ), .C(\UART_TXFF/iFIFOMem[9][4] ), .D(
        \UART_TXFF/iFIFOMem[11][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n146 ) );
  notech_mux4 \UART_TXFF/U151  ( .A(\UART_TXFF/iFIFOMem[12][4] ), .B(
        \UART_TXFF/iFIFOMem[14][4] ), .C(\UART_TXFF/iFIFOMem[13][4] ), .D(
        \UART_TXFF/iFIFOMem[15][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n145 ) );
  notech_mux4 \UART_TXFF/U150  ( .A(\UART_TXFF/n143 ), .B(\UART_TXFF/n141 ), 
        .C(\UART_TXFF/n142 ), .D(\UART_TXFF/n140 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n144 ) );
  notech_mux4 \UART_TXFF/U149  ( .A(\UART_TXFF/iFIFOMem[16][4] ), .B(
        \UART_TXFF/iFIFOMem[18][4] ), .C(\UART_TXFF/iFIFOMem[17][4] ), .D(
        \UART_TXFF/iFIFOMem[19][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n143 ) );
  notech_mux4 \UART_TXFF/U148  ( .A(\UART_TXFF/iFIFOMem[20][4] ), .B(
        \UART_TXFF/iFIFOMem[22][4] ), .C(\UART_TXFF/iFIFOMem[21][4] ), .D(
        \UART_TXFF/iFIFOMem[23][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n142 ) );
  notech_mux4 \UART_TXFF/U147  ( .A(\UART_TXFF/iFIFOMem[24][4] ), .B(
        \UART_TXFF/iFIFOMem[26][4] ), .C(\UART_TXFF/iFIFOMem[25][4] ), .D(
        \UART_TXFF/iFIFOMem[27][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n141 ) );
  notech_mux4 \UART_TXFF/U146  ( .A(\UART_TXFF/iFIFOMem[28][4] ), .B(
        \UART_TXFF/iFIFOMem[30][4] ), .C(\UART_TXFF/iFIFOMem[29][4] ), .D(
        \UART_TXFF/iFIFOMem[31][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n140 ) );
  notech_mux4 \UART_TXFF/U145  ( .A(\UART_TXFF/n138 ), .B(\UART_TXFF/n136 ), 
        .C(\UART_TXFF/n137 ), .D(\UART_TXFF/n135 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n139 ) );
  notech_mux4 \UART_TXFF/U144  ( .A(\UART_TXFF/iFIFOMem[32][4] ), .B(
        \UART_TXFF/iFIFOMem[34][4] ), .C(\UART_TXFF/iFIFOMem[33][4] ), .D(
        \UART_TXFF/iFIFOMem[35][4] ), .S0(\UART_TXFF/n40 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n138 ) );
  notech_mux4 \UART_TXFF/U143  ( .A(\UART_TXFF/iFIFOMem[36][4] ), .B(
        \UART_TXFF/iFIFOMem[38][4] ), .C(\UART_TXFF/iFIFOMem[37][4] ), .D(
        \UART_TXFF/iFIFOMem[39][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n46 ), .Z(\UART_TXFF/n137 ) );
  notech_mux4 \UART_TXFF/U142  ( .A(\UART_TXFF/iFIFOMem[40][4] ), .B(
        \UART_TXFF/iFIFOMem[42][4] ), .C(\UART_TXFF/iFIFOMem[41][4] ), .D(
        \UART_TXFF/iFIFOMem[43][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n136 ) );
  notech_mux4 \UART_TXFF/U141  ( .A(\UART_TXFF/iFIFOMem[44][4] ), .B(
        \UART_TXFF/iFIFOMem[46][4] ), .C(\UART_TXFF/iFIFOMem[45][4] ), .D(
        \UART_TXFF/iFIFOMem[47][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n135 ) );
  notech_mux4 \UART_TXFF/U140  ( .A(\UART_TXFF/n133 ), .B(\UART_TXFF/n131 ), 
        .C(\UART_TXFF/n132 ), .D(\UART_TXFF/n130 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n134 ) );
  notech_mux4 \UART_TXFF/U139  ( .A(\UART_TXFF/iFIFOMem[48][4] ), .B(
        \UART_TXFF/iFIFOMem[50][4] ), .C(\UART_TXFF/iFIFOMem[49][4] ), .D(
        \UART_TXFF/iFIFOMem[51][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n133 ) );
  notech_mux4 \UART_TXFF/U138  ( .A(\UART_TXFF/iFIFOMem[52][4] ), .B(
        \UART_TXFF/iFIFOMem[54][4] ), .C(\UART_TXFF/iFIFOMem[53][4] ), .D(
        \UART_TXFF/iFIFOMem[55][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n132 ) );
  notech_mux4 \UART_TXFF/U137  ( .A(\UART_TXFF/iFIFOMem[56][4] ), .B(
        \UART_TXFF/iFIFOMem[58][4] ), .C(\UART_TXFF/iFIFOMem[57][4] ), .D(
        \UART_TXFF/iFIFOMem[59][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n131 ) );
  notech_mux4 \UART_TXFF/U136  ( .A(\UART_TXFF/iFIFOMem[60][4] ), .B(
        \UART_TXFF/iFIFOMem[62][4] ), .C(\UART_TXFF/iFIFOMem[61][4] ), .D(
        \UART_TXFF/iFIFOMem[63][4] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n130 ) );
  notech_mux4 \UART_TXFF/U135  ( .A(\UART_TXFF/n129 ), .B(\UART_TXFF/n119 ), 
        .C(\UART_TXFF/n124 ), .D(\UART_TXFF/n114 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N127 ) );
  notech_mux4 \UART_TXFF/U134  ( .A(\UART_TXFF/n128 ), .B(\UART_TXFF/n126 ), 
        .C(\UART_TXFF/n127 ), .D(\UART_TXFF/n125 ), .S0(\UART_TXFF/n35 ), .S1(
        \UART_TXFF/n34 ), .Z(\UART_TXFF/n129 ) );
  notech_mux4 \UART_TXFF/U133  ( .A(\UART_TXFF/iFIFOMem[0][3] ), .B(
        \UART_TXFF/iFIFOMem[2][3] ), .C(\UART_TXFF/iFIFOMem[1][3] ), .D(
        \UART_TXFF/iFIFOMem[3][3] ), .S0(\UART_TXFF/n39 ), .S1(\UART_TXFF/n45 ), .Z(\UART_TXFF/n128 ) );
  notech_mux4 \UART_TXFF/U132  ( .A(\UART_TXFF/iFIFOMem[4][3] ), .B(
        \UART_TXFF/iFIFOMem[6][3] ), .C(\UART_TXFF/iFIFOMem[5][3] ), .D(
        \UART_TXFF/iFIFOMem[7][3] ), .S0(\UART_TXFF/n39 ), .S1(\UART_TXFF/n45 ), .Z(\UART_TXFF/n127 ) );
  notech_mux4 \UART_TXFF/U131  ( .A(\UART_TXFF/iFIFOMem[8][3] ), .B(
        \UART_TXFF/iFIFOMem[10][3] ), .C(\UART_TXFF/iFIFOMem[9][3] ), .D(
        \UART_TXFF/iFIFOMem[11][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n126 ) );
  notech_mux4 \UART_TXFF/U130  ( .A(\UART_TXFF/iFIFOMem[12][3] ), .B(
        \UART_TXFF/iFIFOMem[14][3] ), .C(\UART_TXFF/iFIFOMem[13][3] ), .D(
        \UART_TXFF/iFIFOMem[15][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n125 ) );
  notech_mux4 \UART_TXFF/U129  ( .A(\UART_TXFF/n123 ), .B(\UART_TXFF/n121 ), 
        .C(\UART_TXFF/n122 ), .D(\UART_TXFF/n120 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n124 ) );
  notech_mux4 \UART_TXFF/U128  ( .A(\UART_TXFF/iFIFOMem[16][3] ), .B(
        \UART_TXFF/iFIFOMem[18][3] ), .C(\UART_TXFF/iFIFOMem[17][3] ), .D(
        \UART_TXFF/iFIFOMem[19][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n123 ) );
  notech_mux4 \UART_TXFF/U127  ( .A(\UART_TXFF/iFIFOMem[20][3] ), .B(
        \UART_TXFF/iFIFOMem[22][3] ), .C(\UART_TXFF/iFIFOMem[21][3] ), .D(
        \UART_TXFF/iFIFOMem[23][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n122 ) );
  notech_mux4 \UART_TXFF/U126  ( .A(\UART_TXFF/iFIFOMem[24][3] ), .B(
        \UART_TXFF/iFIFOMem[26][3] ), .C(\UART_TXFF/iFIFOMem[25][3] ), .D(
        \UART_TXFF/iFIFOMem[27][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n121 ) );
  notech_mux4 \UART_TXFF/U125  ( .A(\UART_TXFF/iFIFOMem[28][3] ), .B(
        \UART_TXFF/iFIFOMem[30][3] ), .C(\UART_TXFF/iFIFOMem[29][3] ), .D(
        \UART_TXFF/iFIFOMem[31][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n120 ) );
  notech_mux4 \UART_TXFF/U124  ( .A(\UART_TXFF/n118 ), .B(\UART_TXFF/n116 ), 
        .C(\UART_TXFF/n117 ), .D(\UART_TXFF/n115 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n119 ) );
  notech_mux4 \UART_TXFF/U123  ( .A(\UART_TXFF/iFIFOMem[32][3] ), .B(
        \UART_TXFF/iFIFOMem[34][3] ), .C(\UART_TXFF/iFIFOMem[33][3] ), .D(
        \UART_TXFF/iFIFOMem[35][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n118 ) );
  notech_mux4 \UART_TXFF/U122  ( .A(\UART_TXFF/iFIFOMem[36][3] ), .B(
        \UART_TXFF/iFIFOMem[38][3] ), .C(\UART_TXFF/iFIFOMem[37][3] ), .D(
        \UART_TXFF/iFIFOMem[39][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n117 ) );
  notech_mux4 \UART_TXFF/U121  ( .A(\UART_TXFF/iFIFOMem[40][3] ), .B(
        \UART_TXFF/iFIFOMem[42][3] ), .C(\UART_TXFF/iFIFOMem[41][3] ), .D(
        \UART_TXFF/iFIFOMem[43][3] ), .S0(\UART_TXFF/n39 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n116 ) );
  notech_mux4 \UART_TXFF/U120  ( .A(\UART_TXFF/iFIFOMem[44][3] ), .B(
        \UART_TXFF/iFIFOMem[46][3] ), .C(\UART_TXFF/iFIFOMem[45][3] ), .D(
        \UART_TXFF/iFIFOMem[47][3] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n115 ) );
  notech_mux4 \UART_TXFF/U119  ( .A(\UART_TXFF/n113 ), .B(\UART_TXFF/n111 ), 
        .C(\UART_TXFF/n112 ), .D(\UART_TXFF/n110 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n114 ) );
  notech_mux4 \UART_TXFF/U118  ( .A(\UART_TXFF/iFIFOMem[48][3] ), .B(
        \UART_TXFF/iFIFOMem[50][3] ), .C(\UART_TXFF/iFIFOMem[49][3] ), .D(
        \UART_TXFF/iFIFOMem[51][3] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n113 ) );
  notech_mux4 \UART_TXFF/U117  ( .A(\UART_TXFF/iFIFOMem[52][3] ), .B(
        \UART_TXFF/iFIFOMem[54][3] ), .C(\UART_TXFF/iFIFOMem[53][3] ), .D(
        \UART_TXFF/iFIFOMem[55][3] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n112 ) );
  notech_mux4 \UART_TXFF/U116  ( .A(\UART_TXFF/iFIFOMem[56][3] ), .B(
        \UART_TXFF/iFIFOMem[58][3] ), .C(\UART_TXFF/iFIFOMem[57][3] ), .D(
        \UART_TXFF/iFIFOMem[59][3] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n111 ) );
  notech_mux4 \UART_TXFF/U115  ( .A(\UART_TXFF/iFIFOMem[60][3] ), .B(
        \UART_TXFF/iFIFOMem[62][3] ), .C(\UART_TXFF/iFIFOMem[61][3] ), .D(
        \UART_TXFF/iFIFOMem[63][3] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n110 ) );
  notech_mux4 \UART_TXFF/U114  ( .A(\UART_TXFF/n109 ), .B(\UART_TXFF/n99 ), 
        .C(\UART_TXFF/n104 ), .D(\UART_TXFF/n94 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N128 ) );
  notech_mux4 \UART_TXFF/U113  ( .A(\UART_TXFF/n108 ), .B(\UART_TXFF/n106 ), 
        .C(\UART_TXFF/n107 ), .D(\UART_TXFF/n105 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n109 ) );
  notech_mux4 \UART_TXFF/U112  ( .A(\UART_TXFF/iFIFOMem[0][2] ), .B(
        \UART_TXFF/iFIFOMem[2][2] ), .C(\UART_TXFF/iFIFOMem[1][2] ), .D(
        \UART_TXFF/iFIFOMem[3][2] ), .S0(\UART_TXFF/n38 ), .S1(\UART_TXFF/n44 ), .Z(\UART_TXFF/n108 ) );
  notech_mux4 \UART_TXFF/U111  ( .A(\UART_TXFF/iFIFOMem[4][2] ), .B(
        \UART_TXFF/iFIFOMem[6][2] ), .C(\UART_TXFF/iFIFOMem[5][2] ), .D(
        \UART_TXFF/iFIFOMem[7][2] ), .S0(\UART_TXFF/n38 ), .S1(\UART_TXFF/n44 ), .Z(\UART_TXFF/n107 ) );
  notech_mux4 \UART_TXFF/U110  ( .A(\UART_TXFF/iFIFOMem[8][2] ), .B(
        \UART_TXFF/iFIFOMem[10][2] ), .C(\UART_TXFF/iFIFOMem[9][2] ), .D(
        \UART_TXFF/iFIFOMem[11][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n106 ) );
  notech_mux4 \UART_TXFF/U109  ( .A(\UART_TXFF/iFIFOMem[12][2] ), .B(
        \UART_TXFF/iFIFOMem[14][2] ), .C(\UART_TXFF/iFIFOMem[13][2] ), .D(
        \UART_TXFF/iFIFOMem[15][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n105 ) );
  notech_mux4 \UART_TXFF/U108  ( .A(\UART_TXFF/n103 ), .B(\UART_TXFF/n101 ), 
        .C(\UART_TXFF/n102 ), .D(\UART_TXFF/n100 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n104 ) );
  notech_mux4 \UART_TXFF/U107  ( .A(\UART_TXFF/iFIFOMem[16][2] ), .B(
        \UART_TXFF/iFIFOMem[18][2] ), .C(\UART_TXFF/iFIFOMem[17][2] ), .D(
        \UART_TXFF/iFIFOMem[19][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n103 ) );
  notech_mux4 \UART_TXFF/U106  ( .A(\UART_TXFF/iFIFOMem[20][2] ), .B(
        \UART_TXFF/iFIFOMem[22][2] ), .C(\UART_TXFF/iFIFOMem[21][2] ), .D(
        \UART_TXFF/iFIFOMem[23][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n102 ) );
  notech_mux4 \UART_TXFF/U105  ( .A(\UART_TXFF/iFIFOMem[24][2] ), .B(
        \UART_TXFF/iFIFOMem[26][2] ), .C(\UART_TXFF/iFIFOMem[25][2] ), .D(
        \UART_TXFF/iFIFOMem[27][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n101 ) );
  notech_mux4 \UART_TXFF/U104  ( .A(\UART_TXFF/iFIFOMem[28][2] ), .B(
        \UART_TXFF/iFIFOMem[30][2] ), .C(\UART_TXFF/iFIFOMem[29][2] ), .D(
        \UART_TXFF/iFIFOMem[31][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n100 ) );
  notech_mux4 \UART_TXFF/U103  ( .A(\UART_TXFF/n98 ), .B(\UART_TXFF/n96 ), .C(
        \UART_TXFF/n97 ), .D(\UART_TXFF/n95 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n99 ) );
  notech_mux4 \UART_TXFF/U102  ( .A(\UART_TXFF/iFIFOMem[32][2] ), .B(
        \UART_TXFF/iFIFOMem[34][2] ), .C(\UART_TXFF/iFIFOMem[33][2] ), .D(
        \UART_TXFF/iFIFOMem[35][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n98 ) );
  notech_mux4 \UART_TXFF/U101  ( .A(\UART_TXFF/iFIFOMem[36][2] ), .B(
        \UART_TXFF/iFIFOMem[38][2] ), .C(\UART_TXFF/iFIFOMem[37][2] ), .D(
        \UART_TXFF/iFIFOMem[39][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n97 ) );
  notech_mux4 \UART_TXFF/U100  ( .A(\UART_TXFF/iFIFOMem[40][2] ), .B(
        \UART_TXFF/iFIFOMem[42][2] ), .C(\UART_TXFF/iFIFOMem[41][2] ), .D(
        \UART_TXFF/iFIFOMem[43][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n96 ) );
  notech_mux4 \UART_TXFF/U99  ( .A(\UART_TXFF/iFIFOMem[44][2] ), .B(
        \UART_TXFF/iFIFOMem[46][2] ), .C(\UART_TXFF/iFIFOMem[45][2] ), .D(
        \UART_TXFF/iFIFOMem[47][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n95 ) );
  notech_mux4 \UART_TXFF/U98  ( .A(\UART_TXFF/n93 ), .B(\UART_TXFF/n91 ), .C(
        \UART_TXFF/n92 ), .D(\UART_TXFF/n90 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n94 ) );
  notech_mux4 \UART_TXFF/U97  ( .A(\UART_TXFF/iFIFOMem[48][2] ), .B(
        \UART_TXFF/iFIFOMem[50][2] ), .C(\UART_TXFF/iFIFOMem[49][2] ), .D(
        \UART_TXFF/iFIFOMem[51][2] ), .S0(\UART_TXFF/n38 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n93 ) );
  notech_mux4 \UART_TXFF/U96  ( .A(\UART_TXFF/iFIFOMem[52][2] ), .B(
        \UART_TXFF/iFIFOMem[54][2] ), .C(\UART_TXFF/iFIFOMem[53][2] ), .D(
        \UART_TXFF/iFIFOMem[55][2] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n92 ) );
  notech_mux4 \UART_TXFF/U95  ( .A(\UART_TXFF/iFIFOMem[56][2] ), .B(
        \UART_TXFF/iFIFOMem[58][2] ), .C(\UART_TXFF/iFIFOMem[57][2] ), .D(
        \UART_TXFF/iFIFOMem[59][2] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n91 ) );
  notech_mux4 \UART_TXFF/U94  ( .A(\UART_TXFF/iFIFOMem[60][2] ), .B(
        \UART_TXFF/iFIFOMem[62][2] ), .C(\UART_TXFF/iFIFOMem[61][2] ), .D(
        \UART_TXFF/iFIFOMem[63][2] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n90 ) );
  notech_mux4 \UART_TXFF/U93  ( .A(\UART_TXFF/n89 ), .B(\UART_TXFF/n79 ), .C(
        \UART_TXFF/n84 ), .D(\UART_TXFF/n74 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N129 ) );
  notech_mux4 \UART_TXFF/U92  ( .A(\UART_TXFF/n88 ), .B(\UART_TXFF/n86 ), .C(
        \UART_TXFF/n87 ), .D(\UART_TXFF/n85 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n89 ) );
  notech_mux4 \UART_TXFF/U91  ( .A(\UART_TXFF/iFIFOMem[0][1] ), .B(
        \UART_TXFF/iFIFOMem[2][1] ), .C(\UART_TXFF/iFIFOMem[1][1] ), .D(
        \UART_TXFF/iFIFOMem[3][1] ), .S0(\UART_TXFF/n37 ), .S1(\UART_TXFF/n43 ), .Z(\UART_TXFF/n88 ) );
  notech_mux4 \UART_TXFF/U90  ( .A(\UART_TXFF/iFIFOMem[4][1] ), .B(
        \UART_TXFF/iFIFOMem[6][1] ), .C(\UART_TXFF/iFIFOMem[5][1] ), .D(
        \UART_TXFF/iFIFOMem[7][1] ), .S0(\UART_TXFF/n37 ), .S1(\UART_TXFF/n43 ), .Z(\UART_TXFF/n87 ) );
  notech_mux4 \UART_TXFF/U89  ( .A(\UART_TXFF/iFIFOMem[8][1] ), .B(
        \UART_TXFF/iFIFOMem[10][1] ), .C(\UART_TXFF/iFIFOMem[9][1] ), .D(
        \UART_TXFF/iFIFOMem[11][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n86 ) );
  notech_mux4 \UART_TXFF/U88  ( .A(\UART_TXFF/iFIFOMem[12][1] ), .B(
        \UART_TXFF/iFIFOMem[14][1] ), .C(\UART_TXFF/iFIFOMem[13][1] ), .D(
        \UART_TXFF/iFIFOMem[15][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n85 ) );
  notech_mux4 \UART_TXFF/U87  ( .A(\UART_TXFF/n83 ), .B(\UART_TXFF/n81 ), .C(
        \UART_TXFF/n82 ), .D(\UART_TXFF/n80 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n84 ) );
  notech_mux4 \UART_TXFF/U86  ( .A(\UART_TXFF/iFIFOMem[16][1] ), .B(
        \UART_TXFF/iFIFOMem[18][1] ), .C(\UART_TXFF/iFIFOMem[17][1] ), .D(
        \UART_TXFF/iFIFOMem[19][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n83 ) );
  notech_mux4 \UART_TXFF/U85  ( .A(\UART_TXFF/iFIFOMem[20][1] ), .B(
        \UART_TXFF/iFIFOMem[22][1] ), .C(\UART_TXFF/iFIFOMem[21][1] ), .D(
        \UART_TXFF/iFIFOMem[23][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n82 ) );
  notech_mux4 \UART_TXFF/U84  ( .A(\UART_TXFF/iFIFOMem[24][1] ), .B(
        \UART_TXFF/iFIFOMem[26][1] ), .C(\UART_TXFF/iFIFOMem[25][1] ), .D(
        \UART_TXFF/iFIFOMem[27][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n81 ) );
  notech_mux4 \UART_TXFF/U83  ( .A(\UART_TXFF/iFIFOMem[28][1] ), .B(
        \UART_TXFF/iFIFOMem[30][1] ), .C(\UART_TXFF/iFIFOMem[29][1] ), .D(
        \UART_TXFF/iFIFOMem[31][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n80 ) );
  notech_mux4 \UART_TXFF/U82  ( .A(\UART_TXFF/n78 ), .B(\UART_TXFF/n76 ), .C(
        \UART_TXFF/n77 ), .D(\UART_TXFF/n75 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n79 ) );
  notech_mux4 \UART_TXFF/U81  ( .A(\UART_TXFF/iFIFOMem[32][1] ), .B(
        \UART_TXFF/iFIFOMem[34][1] ), .C(\UART_TXFF/iFIFOMem[33][1] ), .D(
        \UART_TXFF/iFIFOMem[35][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n78 ) );
  notech_mux4 \UART_TXFF/U80  ( .A(\UART_TXFF/iFIFOMem[36][1] ), .B(
        \UART_TXFF/iFIFOMem[38][1] ), .C(\UART_TXFF/iFIFOMem[37][1] ), .D(
        \UART_TXFF/iFIFOMem[39][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n77 ) );
  notech_mux4 \UART_TXFF/U79  ( .A(\UART_TXFF/iFIFOMem[40][1] ), .B(
        \UART_TXFF/iFIFOMem[42][1] ), .C(\UART_TXFF/iFIFOMem[41][1] ), .D(
        \UART_TXFF/iFIFOMem[43][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n76 ) );
  notech_mux4 \UART_TXFF/U78  ( .A(\UART_TXFF/iFIFOMem[44][1] ), .B(
        \UART_TXFF/iFIFOMem[46][1] ), .C(\UART_TXFF/iFIFOMem[45][1] ), .D(
        \UART_TXFF/iFIFOMem[47][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n75 ) );
  notech_mux4 \UART_TXFF/U77  ( .A(\UART_TXFF/n73 ), .B(\UART_TXFF/n71 ), .C(
        \UART_TXFF/n72 ), .D(\UART_TXFF/n70 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n74 ) );
  notech_mux4 \UART_TXFF/U76  ( .A(\UART_TXFF/iFIFOMem[48][1] ), .B(
        \UART_TXFF/iFIFOMem[50][1] ), .C(\UART_TXFF/iFIFOMem[49][1] ), .D(
        \UART_TXFF/iFIFOMem[51][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n73 ) );
  notech_mux4 \UART_TXFF/U75  ( .A(\UART_TXFF/iFIFOMem[52][1] ), .B(
        \UART_TXFF/iFIFOMem[54][1] ), .C(\UART_TXFF/iFIFOMem[53][1] ), .D(
        \UART_TXFF/iFIFOMem[55][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n72 ) );
  notech_mux4 \UART_TXFF/U74  ( .A(\UART_TXFF/iFIFOMem[56][1] ), .B(
        \UART_TXFF/iFIFOMem[58][1] ), .C(\UART_TXFF/iFIFOMem[57][1] ), .D(
        \UART_TXFF/iFIFOMem[59][1] ), .S0(\UART_TXFF/n37 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n71 ) );
  notech_mux4 \UART_TXFF/U73  ( .A(\UART_TXFF/iFIFOMem[60][1] ), .B(
        \UART_TXFF/iFIFOMem[62][1] ), .C(\UART_TXFF/iFIFOMem[61][1] ), .D(
        \UART_TXFF/iFIFOMem[63][1] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n70 ) );
  notech_mux4 \UART_TXFF/U72  ( .A(\UART_TXFF/n69 ), .B(\UART_TXFF/n59 ), .C(
        \UART_TXFF/n64 ), .D(\UART_TXFF/n54 ), .S0(\UART_TXFF/N17 ), .S1(
        \UART_TXFF/N16 ), .Z(\UART_TXFF/N130 ) );
  notech_mux4 \UART_TXFF/U71  ( .A(\UART_TXFF/n68 ), .B(\UART_TXFF/n66 ), .C(
        \UART_TXFF/n67 ), .D(\UART_TXFF/n65 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n69 ) );
  notech_mux4 \UART_TXFF/U70  ( .A(\UART_TXFF/iFIFOMem[0][0] ), .B(
        \UART_TXFF/iFIFOMem[2][0] ), .C(\UART_TXFF/iFIFOMem[1][0] ), .D(
        \UART_TXFF/iFIFOMem[3][0] ), .S0(\UART_TXFF/n36 ), .S1(\UART_TXFF/N12 ), .Z(\UART_TXFF/n68 ) );
  notech_mux4 \UART_TXFF/U69  ( .A(\UART_TXFF/iFIFOMem[4][0] ), .B(
        \UART_TXFF/iFIFOMem[6][0] ), .C(\UART_TXFF/iFIFOMem[5][0] ), .D(
        \UART_TXFF/iFIFOMem[7][0] ), .S0(\UART_TXFF/n36 ), .S1(\UART_TXFF/N12 ), .Z(\UART_TXFF/n67 ) );
  notech_mux4 \UART_TXFF/U68  ( .A(\UART_TXFF/iFIFOMem[8][0] ), .B(
        \UART_TXFF/iFIFOMem[10][0] ), .C(\UART_TXFF/iFIFOMem[9][0] ), .D(
        \UART_TXFF/iFIFOMem[11][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n66 ) );
  notech_mux4 \UART_TXFF/U67  ( .A(\UART_TXFF/iFIFOMem[12][0] ), .B(
        \UART_TXFF/iFIFOMem[14][0] ), .C(\UART_TXFF/iFIFOMem[13][0] ), .D(
        \UART_TXFF/iFIFOMem[15][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n65 ) );
  notech_mux4 \UART_TXFF/U66  ( .A(\UART_TXFF/n63 ), .B(\UART_TXFF/n61 ), .C(
        \UART_TXFF/n62 ), .D(\UART_TXFF/n60 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n64 ) );
  notech_mux4 \UART_TXFF/U65  ( .A(\UART_TXFF/iFIFOMem[16][0] ), .B(
        \UART_TXFF/iFIFOMem[18][0] ), .C(\UART_TXFF/iFIFOMem[17][0] ), .D(
        \UART_TXFF/iFIFOMem[19][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n63 ) );
  notech_mux4 \UART_TXFF/U64  ( .A(\UART_TXFF/iFIFOMem[20][0] ), .B(
        \UART_TXFF/iFIFOMem[22][0] ), .C(\UART_TXFF/iFIFOMem[21][0] ), .D(
        \UART_TXFF/iFIFOMem[23][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n62 ) );
  notech_mux4 \UART_TXFF/U63  ( .A(\UART_TXFF/iFIFOMem[24][0] ), .B(
        \UART_TXFF/iFIFOMem[26][0] ), .C(\UART_TXFF/iFIFOMem[25][0] ), .D(
        \UART_TXFF/iFIFOMem[27][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n61 ) );
  notech_mux4 \UART_TXFF/U62  ( .A(\UART_TXFF/iFIFOMem[28][0] ), .B(
        \UART_TXFF/iFIFOMem[30][0] ), .C(\UART_TXFF/iFIFOMem[29][0] ), .D(
        \UART_TXFF/iFIFOMem[31][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n60 ) );
  notech_mux4 \UART_TXFF/U61  ( .A(\UART_TXFF/n58 ), .B(\UART_TXFF/n56 ), .C(
        \UART_TXFF/n57 ), .D(\UART_TXFF/n55 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n59 ) );
  notech_mux4 \UART_TXFF/U60  ( .A(\UART_TXFF/iFIFOMem[32][0] ), .B(
        \UART_TXFF/iFIFOMem[34][0] ), .C(\UART_TXFF/iFIFOMem[33][0] ), .D(
        \UART_TXFF/iFIFOMem[35][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n58 ) );
  notech_mux4 \UART_TXFF/U59  ( .A(\UART_TXFF/iFIFOMem[36][0] ), .B(
        \UART_TXFF/iFIFOMem[38][0] ), .C(\UART_TXFF/iFIFOMem[37][0] ), .D(
        \UART_TXFF/iFIFOMem[39][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n57 ) );
  notech_mux4 \UART_TXFF/U58  ( .A(\UART_TXFF/iFIFOMem[40][0] ), .B(
        \UART_TXFF/iFIFOMem[42][0] ), .C(\UART_TXFF/iFIFOMem[41][0] ), .D(
        \UART_TXFF/iFIFOMem[43][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/N12 ), .Z(\UART_TXFF/n56 ) );
  notech_mux4 \UART_TXFF/U57  ( .A(\UART_TXFF/iFIFOMem[44][0] ), .B(
        \UART_TXFF/iFIFOMem[46][0] ), .C(\UART_TXFF/iFIFOMem[45][0] ), .D(
        \UART_TXFF/iFIFOMem[47][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n43 ), .Z(\UART_TXFF/n55 ) );
  notech_mux4 \UART_TXFF/U56  ( .A(\UART_TXFF/n53 ), .B(\UART_TXFF/n51 ), .C(
        \UART_TXFF/n52 ), .D(\UART_TXFF/n50 ), .S0(\UART_TXFF/N15 ), .S1(
        \UART_TXFF/N14 ), .Z(\UART_TXFF/n54 ) );
  notech_mux4 \UART_TXFF/U55  ( .A(\UART_TXFF/iFIFOMem[48][0] ), .B(
        \UART_TXFF/iFIFOMem[50][0] ), .C(\UART_TXFF/iFIFOMem[49][0] ), .D(
        \UART_TXFF/iFIFOMem[51][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n47 ), .Z(\UART_TXFF/n53 ) );
  notech_mux4 \UART_TXFF/U54  ( .A(\UART_TXFF/iFIFOMem[52][0] ), .B(
        \UART_TXFF/iFIFOMem[54][0] ), .C(\UART_TXFF/iFIFOMem[53][0] ), .D(
        \UART_TXFF/iFIFOMem[55][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n48 ), .Z(\UART_TXFF/n52 ) );
  notech_mux4 \UART_TXFF/U53  ( .A(\UART_TXFF/iFIFOMem[56][0] ), .B(
        \UART_TXFF/iFIFOMem[58][0] ), .C(\UART_TXFF/iFIFOMem[57][0] ), .D(
        \UART_TXFF/iFIFOMem[59][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n44 ), .Z(\UART_TXFF/n51 ) );
  notech_mux4 \UART_TXFF/U52  ( .A(\UART_TXFF/iFIFOMem[60][0] ), .B(
        \UART_TXFF/iFIFOMem[62][0] ), .C(\UART_TXFF/iFIFOMem[61][0] ), .D(
        \UART_TXFF/iFIFOMem[63][0] ), .S0(\UART_TXFF/n36 ), .S1(
        \UART_TXFF/n45 ), .Z(\UART_TXFF/n50 ) );
  notech_inv \UART_TXFF/U51  ( .A(\UART_TXFF/N12 ), .Z(\UART_TXFF/n49 ) );
  notech_inv \UART_TXFF/U50  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n48 ) );
  notech_inv \UART_TXFF/U49  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n47 ) );
  notech_inv \UART_TXFF/U48  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n46 ) );
  notech_inv \UART_TXFF/U47  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n45 ) );
  notech_inv \UART_TXFF/U46  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n44 ) );
  notech_inv \UART_TXFF/U45  ( .A(\UART_TXFF/n49 ), .Z(\UART_TXFF/n43 ) );
  notech_inv \UART_TXFF/U44  ( .A(\UART_TXFF/N13 ), .Z(\UART_TXFF/n42 ) );
  notech_inv \UART_TXFF/U43  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n41 ) );
  notech_inv \UART_TXFF/U42  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n40 ) );
  notech_inv \UART_TXFF/U41  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n39 ) );
  notech_inv \UART_TXFF/U40  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n38 ) );
  notech_inv \UART_TXFF/U39  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n37 ) );
  notech_inv \UART_TXFF/U38  ( .A(\UART_TXFF/n42 ), .Z(\UART_TXFF/n36 ) );
  notech_inv \UART_TXFF/U37  ( .A(\UART_TXFF/n234 ), .Z(\UART_TXFF/n35 ) );
  notech_inv \UART_TXFF/U36  ( .A(\UART_TXFF/n232 ), .Z(\UART_TXFF/n34 ) );
  notech_inv \UART_TXFF/U34  ( .A(\UART_TXFF/n29 ), .Z(\UART_TXFF/n32 ) );
  notech_inv \UART_TXFF/U33  ( .A(\UART_TXFF/n29 ), .Z(\UART_TXFF/n31 ) );
  notech_inv \UART_TXFF/U32  ( .A(\UART_TXFF/n29 ), .Z(\UART_TXFF/n30 ) );
  notech_inv \UART_TXFF/U31  ( .A(iDIN[7]), .Z(\UART_TXFF/n29 ) );
  notech_inv \UART_TXFF/U30  ( .A(\UART_TXFF/n25 ), .Z(\UART_TXFF/n28 ) );
  notech_inv \UART_TXFF/U29  ( .A(\UART_TXFF/n25 ), .Z(\UART_TXFF/n27 ) );
  notech_inv \UART_TXFF/U28  ( .A(\UART_TXFF/n25 ), .Z(\UART_TXFF/n26 ) );
  notech_inv \UART_TXFF/U27  ( .A(iDIN[6]), .Z(\UART_TXFF/n25 ) );
  notech_inv \UART_TXFF/U26  ( .A(\UART_TXFF/n21 ), .Z(\UART_TXFF/n24 ) );
  notech_inv \UART_TXFF/U25  ( .A(\UART_TXFF/n21 ), .Z(\UART_TXFF/n23 ) );
  notech_inv \UART_TXFF/U24  ( .A(\UART_TXFF/n21 ), .Z(\UART_TXFF/n22 ) );
  notech_inv \UART_TXFF/U23  ( .A(iDIN[5]), .Z(\UART_TXFF/n21 ) );
  notech_inv \UART_TXFF/U22  ( .A(\UART_TXFF/n17 ), .Z(\UART_TXFF/n20 ) );
  notech_inv \UART_TXFF/U21  ( .A(\UART_TXFF/n17 ), .Z(\UART_TXFF/n19 ) );
  notech_inv \UART_TXFF/U20  ( .A(\UART_TXFF/n17 ), .Z(\UART_TXFF/n18 ) );
  notech_inv \UART_TXFF/U19  ( .A(iDIN[4]), .Z(\UART_TXFF/n17 ) );
  notech_inv \UART_TXFF/U18  ( .A(\UART_TXFF/n13 ), .Z(\UART_TXFF/n16 ) );
  notech_inv \UART_TXFF/U17  ( .A(\UART_TXFF/n13 ), .Z(\UART_TXFF/n15 ) );
  notech_inv \UART_TXFF/U16  ( .A(\UART_TXFF/n13 ), .Z(\UART_TXFF/n14 ) );
  notech_inv \UART_TXFF/U15  ( .A(iDIN[3]), .Z(\UART_TXFF/n13 ) );
  notech_inv \UART_TXFF/U14  ( .A(\UART_TXFF/n9 ), .Z(\UART_TXFF/n12 ) );
  notech_inv \UART_TXFF/U13  ( .A(\UART_TXFF/n9 ), .Z(\UART_TXFF/n11 ) );
  notech_inv \UART_TXFF/U12  ( .A(\UART_TXFF/n9 ), .Z(\UART_TXFF/n10 ) );
  notech_inv \UART_TXFF/U11  ( .A(iDIN[2]), .Z(\UART_TXFF/n9 ) );
  notech_inv \UART_TXFF/U10  ( .A(\UART_TXFF/n5 ), .Z(\UART_TXFF/n8 ) );
  notech_inv \UART_TXFF/U9  ( .A(\UART_TXFF/n5 ), .Z(\UART_TXFF/n7 ) );
  notech_inv \UART_TXFF/U8  ( .A(\UART_TXFF/n5 ), .Z(\UART_TXFF/n6 ) );
  notech_inv \UART_TXFF/U7  ( .A(iDIN[1]), .Z(\UART_TXFF/n5 ) );
  notech_inv \UART_TXFF/U6  ( .A(\UART_TXFF/n1 ), .Z(\UART_TXFF/n4 ) );
  notech_inv \UART_TXFF/U5  ( .A(\UART_TXFF/n1 ), .Z(\UART_TXFF/n3 ) );
  notech_inv \UART_TXFF/U4  ( .A(\UART_TXFF/n1 ), .Z(\UART_TXFF/n2 ) );
  notech_inv \UART_TXFF/U3  ( .A(iDIN[0]), .Z(\UART_TXFF/n1 ) );
  notech_reg \UART_TXFF/iUSAGE_reg[4]  ( .D(\UART_TXFF/n1287 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(\iTXFIFOUsage[4] ) );
  notech_reg \UART_TXFF/iUSAGE_reg[3]  ( .D(\UART_TXFF/n1288 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_TXFF/USAGE[3] ) );
  notech_reg \UART_TXFF/iUSAGE_reg[2]  ( .D(\UART_TXFF/n1289 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(\UART_TXFF/USAGE[2] ) );
  notech_reg \UART_TXFF/iUSAGE_reg[1]  ( .D(\UART_TXFF/n1290 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(\UART_TXFF/USAGE[1] ) );
  notech_reg \UART_TXFF/iUSAGE_reg[0]  ( .D(\UART_TXFF/n1291 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(\UART_TXFF/USAGE[0] ) );
  notech_reg \UART_TXFF/Q_reg[0]  ( .D(\UART_TXFF/n758 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[0]) );
  notech_reg \UART_TXFF/Q_reg[1]  ( .D(\UART_TXFF/n760 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[1]) );
  notech_reg \UART_TXFF/Q_reg[2]  ( .D(\UART_TXFF/n762 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[2]) );
  notech_reg \UART_TXFF/Q_reg[3]  ( .D(\UART_TXFF/n764 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[3]) );
  notech_reg \UART_TXFF/Q_reg[4]  ( .D(\UART_TXFF/n766 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[4]) );
  notech_reg \UART_TXFF/Q_reg[5]  ( .D(\UART_TXFF/n768 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[5]) );
  notech_reg \UART_TXFF/Q_reg[6]  ( .D(\UART_TXFF/n770 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[6]) );
  notech_reg \UART_TXFF/Q_reg[7]  ( .D(\UART_TXFF/n772 ), .CP(CLK), .CD(1'b1), 
        .Q(iTXFIFOQ[7]) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][0]  ( .D(\UART_TXFF/n1292 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][1]  ( .D(\UART_TXFF/n1293 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][2]  ( .D(\UART_TXFF/n1294 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][3]  ( .D(\UART_TXFF/n1295 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][4]  ( .D(\UART_TXFF/n1296 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][5]  ( .D(\UART_TXFF/n1297 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][6]  ( .D(\UART_TXFF/n1298 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[0][7]  ( .D(\UART_TXFF/n1299 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[0][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][0]  ( .D(\UART_TXFF/n1300 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][1]  ( .D(\UART_TXFF/n1301 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][2]  ( .D(\UART_TXFF/n1302 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][3]  ( .D(\UART_TXFF/n1303 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][4]  ( .D(\UART_TXFF/n1304 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][5]  ( .D(\UART_TXFF/n1305 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][6]  ( .D(\UART_TXFF/n1306 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[1][7]  ( .D(\UART_TXFF/n1307 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[1][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][0]  ( .D(\UART_TXFF/n1308 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][1]  ( .D(\UART_TXFF/n1309 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][2]  ( .D(\UART_TXFF/n1310 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][3]  ( .D(\UART_TXFF/n1311 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][4]  ( .D(\UART_TXFF/n1312 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][5]  ( .D(\UART_TXFF/n1313 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][6]  ( .D(\UART_TXFF/n1314 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[2][7]  ( .D(\UART_TXFF/n1315 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[2][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][0]  ( .D(\UART_TXFF/n1316 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][1]  ( .D(\UART_TXFF/n1317 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][2]  ( .D(\UART_TXFF/n1318 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][3]  ( .D(\UART_TXFF/n1319 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][4]  ( .D(\UART_TXFF/n1320 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][5]  ( .D(\UART_TXFF/n1321 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][6]  ( .D(\UART_TXFF/n1322 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[3][7]  ( .D(\UART_TXFF/n1323 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[3][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][0]  ( .D(\UART_TXFF/n1324 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][1]  ( .D(\UART_TXFF/n1325 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][2]  ( .D(\UART_TXFF/n1326 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][3]  ( .D(\UART_TXFF/n1327 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][4]  ( .D(\UART_TXFF/n1328 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][5]  ( .D(\UART_TXFF/n1329 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][6]  ( .D(\UART_TXFF/n1330 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[4][7]  ( .D(\UART_TXFF/n1331 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[4][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][0]  ( .D(\UART_TXFF/n1332 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][1]  ( .D(\UART_TXFF/n1333 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][2]  ( .D(\UART_TXFF/n1334 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][3]  ( .D(\UART_TXFF/n1335 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][4]  ( .D(\UART_TXFF/n1336 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][5]  ( .D(\UART_TXFF/n1337 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][6]  ( .D(\UART_TXFF/n1338 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[5][7]  ( .D(\UART_TXFF/n1339 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[5][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][0]  ( .D(\UART_TXFF/n1340 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][1]  ( .D(\UART_TXFF/n1341 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][2]  ( .D(\UART_TXFF/n1342 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][3]  ( .D(\UART_TXFF/n1343 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][4]  ( .D(\UART_TXFF/n1344 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][5]  ( .D(\UART_TXFF/n1345 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][6]  ( .D(\UART_TXFF/n1346 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[6][7]  ( .D(\UART_TXFF/n1347 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[6][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][0]  ( .D(\UART_TXFF/n1348 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][1]  ( .D(\UART_TXFF/n1349 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][2]  ( .D(\UART_TXFF/n1350 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][3]  ( .D(\UART_TXFF/n1351 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][4]  ( .D(\UART_TXFF/n1352 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][5]  ( .D(\UART_TXFF/n1353 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][6]  ( .D(\UART_TXFF/n1354 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[7][7]  ( .D(\UART_TXFF/n1355 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[7][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][0]  ( .D(\UART_TXFF/n1356 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][1]  ( .D(\UART_TXFF/n1357 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][2]  ( .D(\UART_TXFF/n1358 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][3]  ( .D(\UART_TXFF/n1359 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][4]  ( .D(\UART_TXFF/n1360 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][5]  ( .D(\UART_TXFF/n1361 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][6]  ( .D(\UART_TXFF/n1362 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[8][7]  ( .D(\UART_TXFF/n1363 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[8][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][0]  ( .D(\UART_TXFF/n1364 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][1]  ( .D(\UART_TXFF/n1365 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][2]  ( .D(\UART_TXFF/n1366 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][3]  ( .D(\UART_TXFF/n1367 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][4]  ( .D(\UART_TXFF/n1368 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][5]  ( .D(\UART_TXFF/n1369 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][6]  ( .D(\UART_TXFF/n1370 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[9][7]  ( .D(\UART_TXFF/n1371 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[9][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][0]  ( .D(\UART_TXFF/n1372 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][1]  ( .D(\UART_TXFF/n1373 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][2]  ( .D(\UART_TXFF/n1374 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][3]  ( .D(\UART_TXFF/n1375 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][4]  ( .D(\UART_TXFF/n1376 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][5]  ( .D(\UART_TXFF/n1377 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][6]  ( .D(\UART_TXFF/n1378 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[10][7]  ( .D(\UART_TXFF/n1379 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[10][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][0]  ( .D(\UART_TXFF/n1380 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][1]  ( .D(\UART_TXFF/n1381 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][2]  ( .D(\UART_TXFF/n1382 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][3]  ( .D(\UART_TXFF/n1383 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][4]  ( .D(\UART_TXFF/n1384 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][5]  ( .D(\UART_TXFF/n1385 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][6]  ( .D(\UART_TXFF/n1386 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[11][7]  ( .D(\UART_TXFF/n1387 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[11][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][0]  ( .D(\UART_TXFF/n1388 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][1]  ( .D(\UART_TXFF/n1389 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][2]  ( .D(\UART_TXFF/n1390 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][3]  ( .D(\UART_TXFF/n1391 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][4]  ( .D(\UART_TXFF/n1392 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][5]  ( .D(\UART_TXFF/n1393 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][6]  ( .D(\UART_TXFF/n1394 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[12][7]  ( .D(\UART_TXFF/n1395 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[12][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][0]  ( .D(\UART_TXFF/n1396 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][1]  ( .D(\UART_TXFF/n1397 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][2]  ( .D(\UART_TXFF/n1398 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][3]  ( .D(\UART_TXFF/n1399 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][4]  ( .D(\UART_TXFF/n1400 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][5]  ( .D(\UART_TXFF/n1401 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][6]  ( .D(\UART_TXFF/n1402 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[13][7]  ( .D(\UART_TXFF/n1403 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[13][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][0]  ( .D(\UART_TXFF/n1404 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][1]  ( .D(\UART_TXFF/n1405 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][2]  ( .D(\UART_TXFF/n1406 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][3]  ( .D(\UART_TXFF/n1407 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][4]  ( .D(\UART_TXFF/n1408 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][5]  ( .D(\UART_TXFF/n1409 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][6]  ( .D(\UART_TXFF/n1410 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[14][7]  ( .D(\UART_TXFF/n1411 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[14][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][0]  ( .D(\UART_TXFF/n1412 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][1]  ( .D(\UART_TXFF/n1413 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][2]  ( .D(\UART_TXFF/n1414 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][3]  ( .D(\UART_TXFF/n1415 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][4]  ( .D(\UART_TXFF/n1416 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][5]  ( .D(\UART_TXFF/n1417 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][6]  ( .D(\UART_TXFF/n1418 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[15][7]  ( .D(\UART_TXFF/n1419 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[15][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][0]  ( .D(\UART_TXFF/n1420 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][1]  ( .D(\UART_TXFF/n1421 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][2]  ( .D(\UART_TXFF/n1422 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][3]  ( .D(\UART_TXFF/n1423 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][4]  ( .D(\UART_TXFF/n1424 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][5]  ( .D(\UART_TXFF/n1425 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][6]  ( .D(\UART_TXFF/n1426 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[16][7]  ( .D(\UART_TXFF/n1427 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[16][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][0]  ( .D(\UART_TXFF/n1428 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][1]  ( .D(\UART_TXFF/n1429 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][2]  ( .D(\UART_TXFF/n1430 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][3]  ( .D(\UART_TXFF/n1431 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][4]  ( .D(\UART_TXFF/n1432 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][5]  ( .D(\UART_TXFF/n1433 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][6]  ( .D(\UART_TXFF/n1434 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[17][7]  ( .D(\UART_TXFF/n1435 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[17][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][0]  ( .D(\UART_TXFF/n1436 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][1]  ( .D(\UART_TXFF/n1437 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][2]  ( .D(\UART_TXFF/n1438 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][3]  ( .D(\UART_TXFF/n1439 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][4]  ( .D(\UART_TXFF/n1440 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][5]  ( .D(\UART_TXFF/n1441 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][6]  ( .D(\UART_TXFF/n1442 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[18][7]  ( .D(\UART_TXFF/n1443 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[18][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][0]  ( .D(\UART_TXFF/n1444 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][1]  ( .D(\UART_TXFF/n1445 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][2]  ( .D(\UART_TXFF/n1446 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][3]  ( .D(\UART_TXFF/n1447 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][4]  ( .D(\UART_TXFF/n1448 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][5]  ( .D(\UART_TXFF/n1449 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][6]  ( .D(\UART_TXFF/n1450 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[19][7]  ( .D(\UART_TXFF/n1451 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[19][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][0]  ( .D(\UART_TXFF/n1452 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][1]  ( .D(\UART_TXFF/n1453 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][2]  ( .D(\UART_TXFF/n1454 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][3]  ( .D(\UART_TXFF/n1455 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][4]  ( .D(\UART_TXFF/n1456 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][5]  ( .D(\UART_TXFF/n1457 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][6]  ( .D(\UART_TXFF/n1458 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[20][7]  ( .D(\UART_TXFF/n1459 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[20][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][0]  ( .D(\UART_TXFF/n1460 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][1]  ( .D(\UART_TXFF/n1461 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][2]  ( .D(\UART_TXFF/n1462 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][3]  ( .D(\UART_TXFF/n1463 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][4]  ( .D(\UART_TXFF/n1464 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][5]  ( .D(\UART_TXFF/n1465 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][6]  ( .D(\UART_TXFF/n1466 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[21][7]  ( .D(\UART_TXFF/n1467 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[21][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][0]  ( .D(\UART_TXFF/n1468 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][1]  ( .D(\UART_TXFF/n1469 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][2]  ( .D(\UART_TXFF/n1470 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][3]  ( .D(\UART_TXFF/n1471 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][4]  ( .D(\UART_TXFF/n1472 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][5]  ( .D(\UART_TXFF/n1473 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][6]  ( .D(\UART_TXFF/n1474 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[22][7]  ( .D(\UART_TXFF/n1475 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[22][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][0]  ( .D(\UART_TXFF/n1476 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][1]  ( .D(\UART_TXFF/n1477 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][2]  ( .D(\UART_TXFF/n1478 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][3]  ( .D(\UART_TXFF/n1479 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][4]  ( .D(\UART_TXFF/n1480 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][5]  ( .D(\UART_TXFF/n1481 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][6]  ( .D(\UART_TXFF/n1482 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[23][7]  ( .D(\UART_TXFF/n1483 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[23][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][0]  ( .D(\UART_TXFF/n1484 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][1]  ( .D(\UART_TXFF/n1485 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][2]  ( .D(\UART_TXFF/n1486 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][3]  ( .D(\UART_TXFF/n1487 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][4]  ( .D(\UART_TXFF/n1488 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][5]  ( .D(\UART_TXFF/n1489 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][6]  ( .D(\UART_TXFF/n1490 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[24][7]  ( .D(\UART_TXFF/n1491 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[24][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][0]  ( .D(\UART_TXFF/n1492 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][1]  ( .D(\UART_TXFF/n1493 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][2]  ( .D(\UART_TXFF/n1494 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][3]  ( .D(\UART_TXFF/n1495 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][4]  ( .D(\UART_TXFF/n1496 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][5]  ( .D(\UART_TXFF/n1497 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][6]  ( .D(\UART_TXFF/n1498 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[25][7]  ( .D(\UART_TXFF/n1499 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[25][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][0]  ( .D(\UART_TXFF/n1500 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][1]  ( .D(\UART_TXFF/n1501 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][2]  ( .D(\UART_TXFF/n1502 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][3]  ( .D(\UART_TXFF/n1503 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][4]  ( .D(\UART_TXFF/n1504 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][5]  ( .D(\UART_TXFF/n1505 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][6]  ( .D(\UART_TXFF/n1506 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[26][7]  ( .D(\UART_TXFF/n1507 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[26][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][0]  ( .D(\UART_TXFF/n1508 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][1]  ( .D(\UART_TXFF/n1509 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][2]  ( .D(\UART_TXFF/n1510 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][3]  ( .D(\UART_TXFF/n1511 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][4]  ( .D(\UART_TXFF/n1512 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][5]  ( .D(\UART_TXFF/n1513 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][6]  ( .D(\UART_TXFF/n1514 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[27][7]  ( .D(\UART_TXFF/n1515 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[27][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][0]  ( .D(\UART_TXFF/n1516 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][1]  ( .D(\UART_TXFF/n1517 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][2]  ( .D(\UART_TXFF/n1518 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][3]  ( .D(\UART_TXFF/n1519 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][4]  ( .D(\UART_TXFF/n1520 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][5]  ( .D(\UART_TXFF/n1521 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][6]  ( .D(\UART_TXFF/n1522 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[28][7]  ( .D(\UART_TXFF/n1523 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[28][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][0]  ( .D(\UART_TXFF/n1524 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][1]  ( .D(\UART_TXFF/n1525 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][2]  ( .D(\UART_TXFF/n1526 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][3]  ( .D(\UART_TXFF/n1527 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][4]  ( .D(\UART_TXFF/n1528 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][5]  ( .D(\UART_TXFF/n1529 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][6]  ( .D(\UART_TXFF/n1530 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[29][7]  ( .D(\UART_TXFF/n1531 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[29][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][0]  ( .D(\UART_TXFF/n1532 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][1]  ( .D(\UART_TXFF/n1533 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][2]  ( .D(\UART_TXFF/n1534 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][3]  ( .D(\UART_TXFF/n1535 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][4]  ( .D(\UART_TXFF/n1536 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][5]  ( .D(\UART_TXFF/n1537 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][6]  ( .D(\UART_TXFF/n1538 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[30][7]  ( .D(\UART_TXFF/n1539 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[30][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][0]  ( .D(\UART_TXFF/n1540 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][1]  ( .D(\UART_TXFF/n1541 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][2]  ( .D(\UART_TXFF/n1542 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][3]  ( .D(\UART_TXFF/n1543 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][4]  ( .D(\UART_TXFF/n1544 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][5]  ( .D(\UART_TXFF/n1545 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][6]  ( .D(\UART_TXFF/n1546 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[31][7]  ( .D(\UART_TXFF/n1547 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[31][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][0]  ( .D(\UART_TXFF/n1548 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][1]  ( .D(\UART_TXFF/n1549 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][2]  ( .D(\UART_TXFF/n1550 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][3]  ( .D(\UART_TXFF/n1551 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][4]  ( .D(\UART_TXFF/n1552 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][5]  ( .D(\UART_TXFF/n1553 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][6]  ( .D(\UART_TXFF/n1554 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[32][7]  ( .D(\UART_TXFF/n1555 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[32][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][0]  ( .D(\UART_TXFF/n1556 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][1]  ( .D(\UART_TXFF/n1557 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][2]  ( .D(\UART_TXFF/n1558 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][3]  ( .D(\UART_TXFF/n1559 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][4]  ( .D(\UART_TXFF/n1560 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][5]  ( .D(\UART_TXFF/n1561 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][6]  ( .D(\UART_TXFF/n1562 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[33][7]  ( .D(\UART_TXFF/n1563 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[33][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][0]  ( .D(\UART_TXFF/n1564 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][1]  ( .D(\UART_TXFF/n1565 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][2]  ( .D(\UART_TXFF/n1566 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][3]  ( .D(\UART_TXFF/n1567 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][4]  ( .D(\UART_TXFF/n1568 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][5]  ( .D(\UART_TXFF/n1569 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][6]  ( .D(\UART_TXFF/n1570 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[34][7]  ( .D(\UART_TXFF/n1571 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[34][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][0]  ( .D(\UART_TXFF/n1572 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][1]  ( .D(\UART_TXFF/n1573 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][2]  ( .D(\UART_TXFF/n1574 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][3]  ( .D(\UART_TXFF/n1575 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][4]  ( .D(\UART_TXFF/n1576 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][5]  ( .D(\UART_TXFF/n1577 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][6]  ( .D(\UART_TXFF/n1578 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[35][7]  ( .D(\UART_TXFF/n1579 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[35][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][0]  ( .D(\UART_TXFF/n1580 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][1]  ( .D(\UART_TXFF/n1581 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][2]  ( .D(\UART_TXFF/n1582 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][3]  ( .D(\UART_TXFF/n1583 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][4]  ( .D(\UART_TXFF/n1584 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][5]  ( .D(\UART_TXFF/n1585 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][6]  ( .D(\UART_TXFF/n1586 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[36][7]  ( .D(\UART_TXFF/n1587 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[36][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][0]  ( .D(\UART_TXFF/n1588 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][1]  ( .D(\UART_TXFF/n1589 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][2]  ( .D(\UART_TXFF/n1590 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][3]  ( .D(\UART_TXFF/n1591 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][4]  ( .D(\UART_TXFF/n1592 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][5]  ( .D(\UART_TXFF/n1593 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][6]  ( .D(\UART_TXFF/n1594 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[37][7]  ( .D(\UART_TXFF/n1595 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[37][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][0]  ( .D(\UART_TXFF/n1596 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][1]  ( .D(\UART_TXFF/n1597 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][2]  ( .D(\UART_TXFF/n1598 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][3]  ( .D(\UART_TXFF/n1599 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][4]  ( .D(\UART_TXFF/n1600 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][5]  ( .D(\UART_TXFF/n1601 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][6]  ( .D(\UART_TXFF/n1602 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[38][7]  ( .D(\UART_TXFF/n1603 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[38][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][0]  ( .D(\UART_TXFF/n1604 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][1]  ( .D(\UART_TXFF/n1605 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][2]  ( .D(\UART_TXFF/n1606 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][3]  ( .D(\UART_TXFF/n1607 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][4]  ( .D(\UART_TXFF/n1608 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][5]  ( .D(\UART_TXFF/n1609 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][6]  ( .D(\UART_TXFF/n1610 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[39][7]  ( .D(\UART_TXFF/n1611 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[39][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][0]  ( .D(\UART_TXFF/n1612 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][1]  ( .D(\UART_TXFF/n1613 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][2]  ( .D(\UART_TXFF/n1614 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][3]  ( .D(\UART_TXFF/n1615 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][4]  ( .D(\UART_TXFF/n1616 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][5]  ( .D(\UART_TXFF/n1617 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][6]  ( .D(\UART_TXFF/n1618 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[40][7]  ( .D(\UART_TXFF/n1619 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[40][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][0]  ( .D(\UART_TXFF/n1620 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][1]  ( .D(\UART_TXFF/n1621 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][2]  ( .D(\UART_TXFF/n1622 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][3]  ( .D(\UART_TXFF/n1623 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][4]  ( .D(\UART_TXFF/n1624 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][5]  ( .D(\UART_TXFF/n1625 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][6]  ( .D(\UART_TXFF/n1626 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[41][7]  ( .D(\UART_TXFF/n1627 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[41][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][0]  ( .D(\UART_TXFF/n1628 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][1]  ( .D(\UART_TXFF/n1629 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][2]  ( .D(\UART_TXFF/n1630 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][3]  ( .D(\UART_TXFF/n1631 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][4]  ( .D(\UART_TXFF/n1632 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][5]  ( .D(\UART_TXFF/n1633 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][6]  ( .D(\UART_TXFF/n1634 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[42][7]  ( .D(\UART_TXFF/n1635 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[42][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][0]  ( .D(\UART_TXFF/n1636 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][1]  ( .D(\UART_TXFF/n1637 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][2]  ( .D(\UART_TXFF/n1638 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][3]  ( .D(\UART_TXFF/n1639 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][4]  ( .D(\UART_TXFF/n1640 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][5]  ( .D(\UART_TXFF/n1641 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][6]  ( .D(\UART_TXFF/n1642 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[43][7]  ( .D(\UART_TXFF/n1643 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[43][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][0]  ( .D(\UART_TXFF/n1644 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][1]  ( .D(\UART_TXFF/n1645 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][2]  ( .D(\UART_TXFF/n1646 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][3]  ( .D(\UART_TXFF/n1647 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][4]  ( .D(\UART_TXFF/n1648 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][5]  ( .D(\UART_TXFF/n1649 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][6]  ( .D(\UART_TXFF/n1650 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[44][7]  ( .D(\UART_TXFF/n1651 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[44][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][0]  ( .D(\UART_TXFF/n1652 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][1]  ( .D(\UART_TXFF/n1653 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][2]  ( .D(\UART_TXFF/n1654 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][3]  ( .D(\UART_TXFF/n1655 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][4]  ( .D(\UART_TXFF/n1656 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][5]  ( .D(\UART_TXFF/n1657 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][6]  ( .D(\UART_TXFF/n1658 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[45][7]  ( .D(\UART_TXFF/n1659 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[45][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][0]  ( .D(\UART_TXFF/n1660 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][1]  ( .D(\UART_TXFF/n1661 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][2]  ( .D(\UART_TXFF/n1662 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][3]  ( .D(\UART_TXFF/n1663 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][4]  ( .D(\UART_TXFF/n1664 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][5]  ( .D(\UART_TXFF/n1665 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][6]  ( .D(\UART_TXFF/n1666 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[46][7]  ( .D(\UART_TXFF/n1667 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[46][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][0]  ( .D(\UART_TXFF/n1668 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][1]  ( .D(\UART_TXFF/n1669 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][2]  ( .D(\UART_TXFF/n1670 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][3]  ( .D(\UART_TXFF/n1671 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][4]  ( .D(\UART_TXFF/n1672 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][5]  ( .D(\UART_TXFF/n1673 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][6]  ( .D(\UART_TXFF/n1674 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[47][7]  ( .D(\UART_TXFF/n1675 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[47][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][0]  ( .D(\UART_TXFF/n1676 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][1]  ( .D(\UART_TXFF/n1677 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][2]  ( .D(\UART_TXFF/n1678 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][3]  ( .D(\UART_TXFF/n1679 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][4]  ( .D(\UART_TXFF/n1680 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][5]  ( .D(\UART_TXFF/n1681 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][6]  ( .D(\UART_TXFF/n1682 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[48][7]  ( .D(\UART_TXFF/n1683 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[48][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][0]  ( .D(\UART_TXFF/n1684 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][1]  ( .D(\UART_TXFF/n1685 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][2]  ( .D(\UART_TXFF/n1686 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][3]  ( .D(\UART_TXFF/n1687 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][4]  ( .D(\UART_TXFF/n1688 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][5]  ( .D(\UART_TXFF/n1689 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][6]  ( .D(\UART_TXFF/n1690 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[49][7]  ( .D(\UART_TXFF/n1691 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[49][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][0]  ( .D(\UART_TXFF/n1692 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][1]  ( .D(\UART_TXFF/n1693 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][2]  ( .D(\UART_TXFF/n1694 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][3]  ( .D(\UART_TXFF/n1695 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][4]  ( .D(\UART_TXFF/n1696 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][5]  ( .D(\UART_TXFF/n1697 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][6]  ( .D(\UART_TXFF/n1698 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[50][7]  ( .D(\UART_TXFF/n1699 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[50][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][0]  ( .D(\UART_TXFF/n1700 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][1]  ( .D(\UART_TXFF/n1701 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][2]  ( .D(\UART_TXFF/n1702 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][3]  ( .D(\UART_TXFF/n1703 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][4]  ( .D(\UART_TXFF/n1704 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][5]  ( .D(\UART_TXFF/n1705 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][6]  ( .D(\UART_TXFF/n1706 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[51][7]  ( .D(\UART_TXFF/n1707 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[51][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][0]  ( .D(\UART_TXFF/n1708 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][1]  ( .D(\UART_TXFF/n1709 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][2]  ( .D(\UART_TXFF/n1710 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][3]  ( .D(\UART_TXFF/n1711 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][4]  ( .D(\UART_TXFF/n1712 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][5]  ( .D(\UART_TXFF/n1713 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][6]  ( .D(\UART_TXFF/n1714 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[52][7]  ( .D(\UART_TXFF/n1715 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[52][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][0]  ( .D(\UART_TXFF/n1716 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][1]  ( .D(\UART_TXFF/n1717 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][2]  ( .D(\UART_TXFF/n1718 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][3]  ( .D(\UART_TXFF/n1719 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][4]  ( .D(\UART_TXFF/n1720 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][5]  ( .D(\UART_TXFF/n1721 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][6]  ( .D(\UART_TXFF/n1722 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[53][7]  ( .D(\UART_TXFF/n1723 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[53][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][0]  ( .D(\UART_TXFF/n1724 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][1]  ( .D(\UART_TXFF/n1725 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][2]  ( .D(\UART_TXFF/n1726 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][3]  ( .D(\UART_TXFF/n1727 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][4]  ( .D(\UART_TXFF/n1728 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][5]  ( .D(\UART_TXFF/n1729 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][6]  ( .D(\UART_TXFF/n1730 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[54][7]  ( .D(\UART_TXFF/n1731 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[54][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][0]  ( .D(\UART_TXFF/n1732 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][1]  ( .D(\UART_TXFF/n1733 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][2]  ( .D(\UART_TXFF/n1734 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][3]  ( .D(\UART_TXFF/n1735 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][4]  ( .D(\UART_TXFF/n1736 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][5]  ( .D(\UART_TXFF/n1737 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][6]  ( .D(\UART_TXFF/n1738 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[55][7]  ( .D(\UART_TXFF/n1739 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[55][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][0]  ( .D(\UART_TXFF/n1740 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][1]  ( .D(\UART_TXFF/n1741 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][2]  ( .D(\UART_TXFF/n1742 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][3]  ( .D(\UART_TXFF/n1743 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][4]  ( .D(\UART_TXFF/n1744 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][5]  ( .D(\UART_TXFF/n1745 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][6]  ( .D(\UART_TXFF/n1746 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[56][7]  ( .D(\UART_TXFF/n1747 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[56][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][0]  ( .D(\UART_TXFF/n1748 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][1]  ( .D(\UART_TXFF/n1749 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][2]  ( .D(\UART_TXFF/n1750 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][3]  ( .D(\UART_TXFF/n1751 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][4]  ( .D(\UART_TXFF/n1752 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][5]  ( .D(\UART_TXFF/n1753 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][6]  ( .D(\UART_TXFF/n1754 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[57][7]  ( .D(\UART_TXFF/n1755 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[57][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][0]  ( .D(\UART_TXFF/n1756 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][1]  ( .D(\UART_TXFF/n1757 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][2]  ( .D(\UART_TXFF/n1758 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][3]  ( .D(\UART_TXFF/n1759 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][4]  ( .D(\UART_TXFF/n1760 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][5]  ( .D(\UART_TXFF/n1761 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][6]  ( .D(\UART_TXFF/n1762 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[58][7]  ( .D(\UART_TXFF/n1763 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[58][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][0]  ( .D(\UART_TXFF/n1764 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][1]  ( .D(\UART_TXFF/n1765 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][2]  ( .D(\UART_TXFF/n1766 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][3]  ( .D(\UART_TXFF/n1767 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][4]  ( .D(\UART_TXFF/n1768 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][5]  ( .D(\UART_TXFF/n1769 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][6]  ( .D(\UART_TXFF/n1770 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[59][7]  ( .D(\UART_TXFF/n1771 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[59][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][0]  ( .D(\UART_TXFF/n1772 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][1]  ( .D(\UART_TXFF/n1773 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][2]  ( .D(\UART_TXFF/n1774 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][3]  ( .D(\UART_TXFF/n1775 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][4]  ( .D(\UART_TXFF/n1776 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][5]  ( .D(\UART_TXFF/n1777 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][6]  ( .D(\UART_TXFF/n1778 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[60][7]  ( .D(\UART_TXFF/n1779 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[60][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][0]  ( .D(\UART_TXFF/n1780 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][1]  ( .D(\UART_TXFF/n1781 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][2]  ( .D(\UART_TXFF/n1782 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][3]  ( .D(\UART_TXFF/n1783 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][4]  ( .D(\UART_TXFF/n1784 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][5]  ( .D(\UART_TXFF/n1785 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][6]  ( .D(\UART_TXFF/n1786 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[61][7]  ( .D(\UART_TXFF/n1787 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[61][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][0]  ( .D(\UART_TXFF/n1788 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][1]  ( .D(\UART_TXFF/n1789 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][2]  ( .D(\UART_TXFF/n1790 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][3]  ( .D(\UART_TXFF/n1791 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][4]  ( .D(\UART_TXFF/n1792 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][5]  ( .D(\UART_TXFF/n1793 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][6]  ( .D(\UART_TXFF/n1794 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[62][7]  ( .D(\UART_TXFF/n1795 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[62][7] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][0]  ( .D(\UART_TXFF/n1796 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][0] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][1]  ( .D(\UART_TXFF/n1797 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][1] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][2]  ( .D(\UART_TXFF/n1798 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][2] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][3]  ( .D(\UART_TXFF/n1799 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][3] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][4]  ( .D(\UART_TXFF/n1800 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][4] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][5]  ( .D(\UART_TXFF/n1801 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][5] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][6]  ( .D(\UART_TXFF/n1802 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][6] ) );
  notech_reg \UART_TXFF/iFIFOMem_reg[63][7]  ( .D(\UART_TXFF/n1803 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_TXFF/iFIFOMem[63][7] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[5]  ( .D(\UART_TXFF/n1810 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_TXFF/iWRAddr[5] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[4]  ( .D(\UART_TXFF/n1811 ), .CP(CLK), 
        .CD(\UART_IS_DSR/n1 ), .Q(\UART_TXFF/iWRAddr[4] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[3]  ( .D(\UART_TXFF/n1812 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_TXFF/iWRAddr[3] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[2]  ( .D(\UART_TXFF/n1813 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_TXFF/iWRAddr[2] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[1]  ( .D(\UART_TXFF/n1814 ), .CP(CLK), 
        .CD(\UART_IS_SIN/n1 ), .Q(\UART_TXFF/iWRAddr[1] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[0]  ( .D(\UART_TXFF/n1815 ), .CP(CLK), 
        .CD(\UART_IS_SIN/n1 ), .Q(\UART_TXFF/iWRAddr[0] ) );
  notech_reg \UART_TXFF/iWRAddr_reg[6]  ( .D(\UART_TXFF/n1816 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_TXFF/iWRAddr[6] ) );
  notech_reg \UART_TXFF/iRDAddr_reg[5]  ( .D(\UART_TXFF/n1804 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_TXFF/N17 ) );
  notech_reg \UART_TXFF/iRDAddr_reg[4]  ( .D(\UART_TXFF/n1805 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_TXFF/N16 ) );
  notech_reg \UART_TXFF/iRDAddr_reg[3]  ( .D(\UART_TXFF/n1806 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_TXFF/N15 ) );
  notech_reg \UART_TXFF/iRDAddr_reg[2]  ( .D(\UART_TXFF/n1807 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_TXFF/N14 ) );
  notech_reg \UART_TXFF/iRDAddr_reg[1]  ( .D(\UART_TXFF/n1808 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_TXFF/N13 ) );
  notech_reg \UART_TXFF/iRDAddr_reg[6]  ( .D(\UART_TXFF/n1809 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_TXFF/iRDAddr[6] ) );
  notech_reg_set \UART_TXFF/iEMPTY_reg  ( .D(\UART_TXFF/N56 ), .CP(CLK), .SD(
        \UART_IS_SIN/n1 ), .Q(iTXFIFOEmpty) );
  notech_reg \UART_TXFF/iRDAddr_reg[0]  ( .D(\UART_TXFF/n1817 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_TXFF/N12 ) );
  notech_xor2 \UART_TXFF/add_73/U1  ( .A(\UART_TXFF/add_73/carry [6]), .B(
        \UART_TXFF/iWRAddr[6] ), .Z(\UART_TXFF/N30 ) );
  notech_ha2 \UART_TXFF/add_73/U1_1_1  ( .A(\UART_TXFF/iWRAddr[1] ), .B(
        \UART_TXFF/iWRAddr[0] ), .CO(\UART_TXFF/add_73/carry [2]), .Z(
        \UART_TXFF/N25 ) );
  notech_ha2 \UART_TXFF/add_73/U1_1_2  ( .A(\UART_TXFF/iWRAddr[2] ), .B(
        \UART_TXFF/add_73/carry [2]), .CO(\UART_TXFF/add_73/carry [3]), .Z(
        \UART_TXFF/N26 ) );
  notech_ha2 \UART_TXFF/add_73/U1_1_3  ( .A(\UART_TXFF/iWRAddr[3] ), .B(
        \UART_TXFF/add_73/carry [3]), .CO(\UART_TXFF/add_73/carry [4]), .Z(
        \UART_TXFF/N27 ) );
  notech_ha2 \UART_TXFF/add_73/U1_1_4  ( .A(\UART_TXFF/iWRAddr[4] ), .B(
        \UART_TXFF/add_73/carry [4]), .CO(\UART_TXFF/add_73/carry [5]), .Z(
        \UART_TXFF/N28 ) );
  notech_ha2 \UART_TXFF/add_73/U1_1_5  ( .A(\UART_TXFF/iWRAddr[5] ), .B(
        \UART_TXFF/add_73/carry [5]), .CO(\UART_TXFF/add_73/carry [6]), .Z(
        \UART_TXFF/N29 ) );
  notech_xor2 \UART_TXFF/add_77/U1  ( .A(\UART_TXFF/add_77/carry [6]), .B(
        \UART_TXFF/iRDAddr[6] ), .Z(\UART_TXFF/N38 ) );
  notech_ha2 \UART_TXFF/add_77/U1_1_1  ( .A(\UART_TXFF/n36 ), .B(
        \UART_TXFF/n46 ), .CO(\UART_TXFF/add_77/carry [2]), .Z(\UART_TXFF/N33 ) );
  notech_ha2 \UART_TXFF/add_77/U1_1_2  ( .A(\UART_TXFF/N14 ), .B(
        \UART_TXFF/add_77/carry [2]), .CO(\UART_TXFF/add_77/carry [3]), .Z(
        \UART_TXFF/N34 ) );
  notech_ha2 \UART_TXFF/add_77/U1_1_3  ( .A(\UART_TXFF/N15 ), .B(
        \UART_TXFF/add_77/carry [3]), .CO(\UART_TXFF/add_77/carry [4]), .Z(
        \UART_TXFF/N35 ) );
  notech_ha2 \UART_TXFF/add_77/U1_1_4  ( .A(\UART_TXFF/N16 ), .B(
        \UART_TXFF/add_77/carry [4]), .CO(\UART_TXFF/add_77/carry [5]), .Z(
        \UART_TXFF/N36 ) );
  notech_ha2 \UART_TXFF/add_77/U1_1_5  ( .A(\UART_TXFF/N17 ), .B(
        \UART_TXFF/add_77/carry [5]), .CO(\UART_TXFF/add_77/carry [6]), .Z(
        \UART_TXFF/N37 ) );
  notech_xor2 \UART_RXFF/U1202  ( .A(\UART_RXFF/iWRAddr[1] ), .B(
        \UART_RXFF/N13 ), .Z(\UART_RXFF/n445 ) );
  notech_xor2 \UART_RXFF/U1201  ( .A(\UART_RXFF/iWRAddr[5] ), .B(
        \UART_RXFF/N17 ), .Z(\UART_RXFF/n446 ) );
  notech_xor2 \UART_RXFF/U1200  ( .A(\UART_RXFF/iWRAddr[0] ), .B(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n447 ) );
  notech_xor2 \UART_RXFF/U1199  ( .A(\UART_RXFF/n46 ), .B(
        \UART_RXFF/iWRAddr[2] ), .Z(\UART_RXFF/n449 ) );
  notech_xor2 \UART_RXFF/U1198  ( .A(\UART_RXFF/n49 ), .B(
        \UART_RXFF/iWRAddr[3] ), .Z(\UART_RXFF/n450 ) );
  notech_inv \UART_RXFF/U1197  ( .A(\UART_RXFF/N16 ), .Z(\UART_RXFF/n314 ) );
  notech_xor2 \UART_RXFF/U1196  ( .A(\UART_RXFF/n314 ), .B(
        \UART_RXFF/iWRAddr[4] ), .Z(\UART_RXFF/n451 ) );
  notech_nand3 \UART_RXFF/U1195  ( .A(\UART_RXFF/n449 ), .B(\UART_RXFF/n450 ), 
        .C(\UART_RXFF/n451 ), .Z(\UART_RXFF/n448 ) );
  notech_nor4 \UART_RXFF/U1194  ( .A(\UART_RXFF/n445 ), .B(\UART_RXFF/n446 ), 
        .C(\UART_RXFF/n447 ), .D(\UART_RXFF/n448 ), .Z(\UART_RXFF/n442 ) );
  notech_inv \UART_RXFF/U1193  ( .A(\UART_RXFF/n442 ), .Z(\UART_RXFF/n444 ) );
  notech_inv \UART_RXFF/U1192  ( .A(\UART_RXFF/iWRAddr[6] ), .Z(
        \UART_RXFF/n293 ) );
  notech_xor2 \UART_RXFF/U1191  ( .A(\UART_RXFF/iRDAddr[6] ), .B(
        \UART_RXFF/n293 ), .Z(\UART_RXFF/n443 ) );
  notech_nor2 \UART_RXFF/U1190  ( .A(\UART_RXFF/n444 ), .B(\UART_RXFF/n443 ), 
        .Z(iRXFIFO64Full) );
  notech_and2 \UART_RXFF/U1189  ( .A(\UART_RXFF/n442 ), .B(\UART_RXFF/n443 ), 
        .Z(\UART_RXFF/N56 ) );
  notech_and3 \UART_RXFF/U1188  ( .A(iRXFIFOUsage[2]), .B(\UART_RXFF/USAGE[0] ), .C(iRXFIFOUsage[1]), .Z(\UART_RXFF/n424 ) );
  notech_inv \UART_RXFF/U1187  ( .A(iRXFIFOWrite), .Z(\UART_RXFF/n441 ) );
  notech_nand3 \UART_RXFF/U1185  ( .A(\UART_RXFF/n441 ), .B(n371), .C(n438), 
        .Z(\UART_RXFF/n436 ) );
  notech_nor2 \UART_RXFF/U1184  ( .A(iRXFIFO64Full), .B(\UART_RXFF/n441 ), .Z(
        \UART_RXFF/n365 ) );
  notech_or2 \UART_RXFF/U1183  ( .A(\UART_RXFF/n365 ), .B(iRXFIFOClear), .Z(
        \UART_RXFF/n294 ) );
  notech_inv \UART_RXFF/U1182  ( .A(iRXFIFOClear), .Z(\UART_RXFF/n308 ) );
  notech_nand2 \UART_RXFF/U1181  ( .A(\UART_RXFF/n308 ), .B(n371), .Z(
        \UART_RXFF/n440 ) );
  notech_nand2 \UART_RXFF/U1180  ( .A(\UART_RXFF/n294 ), .B(\UART_RXFF/n440 ), 
        .Z(\UART_RXFF/n439 ) );
  notech_nand2 \UART_RXFF/U1179  ( .A(\UART_RXFF/n439 ), .B(\UART_RXFF/n436 ), 
        .Z(\UART_RXFF/n406 ) );
  notech_ao3 \UART_RXFF/U1178  ( .A(\UART_RXFF/n436 ), .B(\UART_RXFF/n406 ), 
        .C(iRXFIFOClear), .Z(\UART_RXFF/n412 ) );
  notech_and3 \UART_RXFF/U1177  ( .A(\UART_RXFF/n424 ), .B(iRXFIFOUsage[3]), 
        .C(\UART_RXFF/n412 ), .Z(\UART_RXFF/n427 ) );
  notech_and2 \UART_RXFF/U1176  ( .A(\UART_RXFF/n427 ), .B(iRXFIFOUsage[4]), 
        .Z(\UART_RXFF/n435 ) );
  notech_inv \UART_RXFF/U1175  ( .A(iRXFIFOUsage[1]), .Z(\UART_RXFF/n437 ) );
  notech_inv \UART_RXFF/U1174  ( .A(\UART_RXFF/USAGE[0] ), .Z(\UART_RXFF/n438 ) );
  notech_ao3 \UART_RXFF/U1173  ( .A(\UART_RXFF/n437 ), .B(\UART_RXFF/n438 ), 
        .C(iRXFIFOUsage[2]), .Z(\UART_RXFF/n415 ) );
  notech_or2 \UART_RXFF/U1172  ( .A(\UART_RXFF/n436 ), .B(iRXFIFOClear), .Z(
        \UART_RXFF/n408 ) );
  notech_inv \UART_RXFF/U1171  ( .A(\UART_RXFF/n408 ), .Z(\UART_RXFF/n411 ) );
  notech_nao3 \UART_RXFF/U1170  ( .C(iRXFIFOUsage[3]), .A(\UART_RXFF/n415 ), 
        .B(\UART_RXFF/n411 ), .Z(\UART_RXFF/n421 ) );
  notech_nor2 \UART_RXFF/U1169  ( .A(\UART_RXFF/n421 ), .B(iRXFIFOUsage[4]), 
        .Z(\UART_RXFF/n426 ) );
  notech_or2 \UART_RXFF/U1168  ( .A(\UART_RXFF/n435 ), .B(\UART_RXFF/n426 ), 
        .Z(\UART_RXFF/n429 ) );
  notech_or2 \UART_RXFF/U1167  ( .A(\UART_RXFF/n408 ), .B(\UART_RXFF/n415 ), 
        .Z(\UART_RXFF/n433 ) );
  notech_inv \UART_RXFF/U1166  ( .A(\UART_RXFF/n412 ), .Z(\UART_RXFF/n407 ) );
  notech_or2 \UART_RXFF/U1165  ( .A(\UART_RXFF/n407 ), .B(\UART_RXFF/n424 ), 
        .Z(\UART_RXFF/n434 ) );
  notech_and3 \UART_RXFF/U1164  ( .A(\UART_RXFF/n433 ), .B(\UART_RXFF/n434 ), 
        .C(\UART_RXFF/n406 ), .Z(\UART_RXFF/n423 ) );
  notech_mux2 \UART_RXFF/U1163  ( .A(\UART_RXFF/n407 ), .B(\UART_RXFF/n408 ), 
        .S(iRXFIFOUsage[3]), .Z(\UART_RXFF/n432 ) );
  notech_nand2 \UART_RXFF/U1162  ( .A(\UART_RXFF/n423 ), .B(\UART_RXFF/n432 ), 
        .Z(\UART_RXFF/n428 ) );
  notech_mux2 \UART_RXFF/U1161  ( .A(\UART_RXFF/n412 ), .B(\UART_RXFF/n411 ), 
        .S(iRXFIFOUsage[4]), .Z(\UART_RXFF/n431 ) );
  notech_or2 \UART_RXFF/U1160  ( .A(\UART_RXFF/n428 ), .B(\UART_RXFF/n431 ), 
        .Z(\UART_RXFF/n430 ) );
  notech_mux2 \UART_RXFF/U1159  ( .A(\UART_RXFF/n429 ), .B(\UART_RXFF/n430 ), 
        .S(iRXFIFOUsage[5]), .Z(\UART_RXFF/n1685 ) );
  notech_mux2 \UART_RXFF/U1158  ( .A(\UART_RXFF/n427 ), .B(\UART_RXFF/n428 ), 
        .S(iRXFIFOUsage[4]), .Z(\UART_RXFF/n425 ) );
  notech_or2 \UART_RXFF/U1157  ( .A(\UART_RXFF/n425 ), .B(\UART_RXFF/n426 ), 
        .Z(\UART_RXFF/n1686 ) );
  notech_nand2 \UART_RXFF/U1156  ( .A(\UART_RXFF/n412 ), .B(\UART_RXFF/n424 ), 
        .Z(\UART_RXFF/n422 ) );
  notech_mux2 \UART_RXFF/U1155  ( .A(\UART_RXFF/n422 ), .B(\UART_RXFF/n423 ), 
        .S(iRXFIFOUsage[3]), .Z(\UART_RXFF/n420 ) );
  notech_nand2 \UART_RXFF/U1154  ( .A(\UART_RXFF/n420 ), .B(\UART_RXFF/n421 ), 
        .Z(\UART_RXFF/n1687 ) );
  notech_nand3 \UART_RXFF/U1153  ( .A(\UART_RXFF/n412 ), .B(
        \UART_RXFF/USAGE[0] ), .C(iRXFIFOUsage[1]), .Z(\UART_RXFF/n416 ) );
  notech_mux2 \UART_RXFF/U1152  ( .A(\UART_RXFF/n407 ), .B(\UART_RXFF/n408 ), 
        .S(\UART_RXFF/USAGE[0] ), .Z(\UART_RXFF/n419 ) );
  notech_nand2 \UART_RXFF/U1151  ( .A(\UART_RXFF/n419 ), .B(\UART_RXFF/n406 ), 
        .Z(\UART_RXFF/n410 ) );
  notech_mux2 \UART_RXFF/U1150  ( .A(\UART_RXFF/n412 ), .B(\UART_RXFF/n411 ), 
        .S(iRXFIFOUsage[1]), .Z(\UART_RXFF/n418 ) );
  notech_nor2 \UART_RXFF/U1149  ( .A(\UART_RXFF/n410 ), .B(\UART_RXFF/n418 ), 
        .Z(\UART_RXFF/n417 ) );
  notech_mux2 \UART_RXFF/U1148  ( .A(\UART_RXFF/n416 ), .B(\UART_RXFF/n417 ), 
        .S(iRXFIFOUsage[2]), .Z(\UART_RXFF/n413 ) );
  notech_nand2 \UART_RXFF/U1147  ( .A(\UART_RXFF/n411 ), .B(\UART_RXFF/n415 ), 
        .Z(\UART_RXFF/n414 ) );
  notech_nand2 \UART_RXFF/U1146  ( .A(\UART_RXFF/n413 ), .B(\UART_RXFF/n414 ), 
        .Z(\UART_RXFF/n1688 ) );
  notech_mux2 \UART_RXFF/U1145  ( .A(\UART_RXFF/n411 ), .B(\UART_RXFF/n412 ), 
        .S(\UART_RXFF/USAGE[0] ), .Z(\UART_RXFF/n409 ) );
  notech_mux2 \UART_RXFF/U1144  ( .A(\UART_RXFF/n409 ), .B(\UART_RXFF/n410 ), 
        .S(iRXFIFOUsage[1]), .Z(\UART_RXFF/n1689 ) );
  notech_nand2 \UART_RXFF/U1143  ( .A(\UART_RXFF/n407 ), .B(\UART_RXFF/n408 ), 
        .Z(\UART_RXFF/n404 ) );
  notech_inv \UART_RXFF/U1142  ( .A(\UART_RXFF/n406 ), .Z(\UART_RXFF/n405 ) );
  notech_mux2 \UART_RXFF/U1141  ( .A(\UART_RXFF/n404 ), .B(\UART_RXFF/n405 ), 
        .S(\UART_RXFF/USAGE[0] ), .Z(\UART_RXFF/n1690 ) );
  notech_inv \UART_RXFF/U1140  ( .A(\UART_RXFF/iWRAddr[3] ), .Z(
        \UART_RXFF/n302 ) );
  notech_ao3 \UART_RXFF/U1138  ( .A(\UART_IS_RI/n1 ), .B(\UART_RXFF/n365 ), 
        .C(\UART_RXFF/iWRAddr[5] ), .Z(\UART_RXFF/n375 ) );
  notech_ao3 \UART_RXFF/U1137  ( .A(\UART_RXFF/n302 ), .B(\UART_RXFF/n375 ), 
        .C(\UART_RXFF/iWRAddr[4] ), .Z(\UART_RXFF/n395 ) );
  notech_inv \UART_RXFF/U1136  ( .A(\UART_RXFF/iWRAddr[0] ), .Z(
        \UART_RXFF/n397 ) );
  notech_inv \UART_RXFF/U1135  ( .A(\UART_RXFF/iWRAddr[2] ), .Z(
        \UART_RXFF/n300 ) );
  notech_inv \UART_RXFF/U1134  ( .A(\UART_RXFF/iWRAddr[1] ), .Z(
        \UART_RXFF/n298 ) );
  notech_and3 \UART_RXFF/U1133  ( .A(\UART_RXFF/n397 ), .B(\UART_RXFF/n300 ), 
        .C(\UART_RXFF/n298 ), .Z(\UART_RXFF/n336 ) );
  notech_and2 \UART_RXFF/U1132  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n403 ) );
  notech_mux2 \UART_RXFF/U1131  ( .A(\UART_RXFF/iFIFOMem[0][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1691 ) );
  notech_mux2 \UART_RXFF/U1130  ( .A(\UART_RXFF/iFIFOMem[0][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1692 ) );
  notech_mux2 \UART_RXFF/U1129  ( .A(\UART_RXFF/iFIFOMem[0][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1693 ) );
  notech_mux2 \UART_RXFF/U1128  ( .A(\UART_RXFF/iFIFOMem[0][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1694 ) );
  notech_mux2 \UART_RXFF/U1127  ( .A(\UART_RXFF/iFIFOMem[0][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1695 ) );
  notech_mux2 \UART_RXFF/U1126  ( .A(\UART_RXFF/iFIFOMem[0][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1696 ) );
  notech_mux2 \UART_RXFF/U1125  ( .A(\UART_RXFF/iFIFOMem[0][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1697 ) );
  notech_mux2 \UART_RXFF/U1124  ( .A(\UART_RXFF/iFIFOMem[0][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1698 ) );
  notech_mux2 \UART_RXFF/U1123  ( .A(\UART_RXFF/iFIFOMem[0][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1699 ) );
  notech_mux2 \UART_RXFF/U1122  ( .A(\UART_RXFF/iFIFOMem[0][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1700 ) );
  notech_mux2 \UART_RXFF/U1121  ( .A(\UART_RXFF/iFIFOMem[0][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n403 ), .Z(\UART_RXFF/n1701 ) );
  notech_and3 \UART_RXFF/U1120  ( .A(\UART_RXFF/iWRAddr[0] ), .B(
        \UART_RXFF/n300 ), .C(\UART_RXFF/n298 ), .Z(\UART_RXFF/n334 ) );
  notech_and2 \UART_RXFF/U1119  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n402 ) );
  notech_mux2 \UART_RXFF/U1118  ( .A(\UART_RXFF/iFIFOMem[1][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1702 ) );
  notech_mux2 \UART_RXFF/U1117  ( .A(\UART_RXFF/iFIFOMem[1][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1703 ) );
  notech_mux2 \UART_RXFF/U1116  ( .A(\UART_RXFF/iFIFOMem[1][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1704 ) );
  notech_mux2 \UART_RXFF/U1115  ( .A(\UART_RXFF/iFIFOMem[1][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1705 ) );
  notech_mux2 \UART_RXFF/U1114  ( .A(\UART_RXFF/iFIFOMem[1][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1706 ) );
  notech_mux2 \UART_RXFF/U1113  ( .A(\UART_RXFF/iFIFOMem[1][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1707 ) );
  notech_mux2 \UART_RXFF/U1112  ( .A(\UART_RXFF/iFIFOMem[1][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1708 ) );
  notech_mux2 \UART_RXFF/U1111  ( .A(\UART_RXFF/iFIFOMem[1][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1709 ) );
  notech_mux2 \UART_RXFF/U1110  ( .A(\UART_RXFF/iFIFOMem[1][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1710 ) );
  notech_mux2 \UART_RXFF/U1109  ( .A(\UART_RXFF/iFIFOMem[1][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1711 ) );
  notech_mux2 \UART_RXFF/U1108  ( .A(\UART_RXFF/iFIFOMem[1][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n402 ), .Z(\UART_RXFF/n1712 ) );
  notech_and3 \UART_RXFF/U1107  ( .A(\UART_RXFF/iWRAddr[1] ), .B(
        \UART_RXFF/n300 ), .C(\UART_RXFF/n397 ), .Z(\UART_RXFF/n332 ) );
  notech_and2 \UART_RXFF/U1106  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n401 ) );
  notech_mux2 \UART_RXFF/U1105  ( .A(\UART_RXFF/iFIFOMem[2][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1713 ) );
  notech_mux2 \UART_RXFF/U1104  ( .A(\UART_RXFF/iFIFOMem[2][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1714 ) );
  notech_mux2 \UART_RXFF/U1103  ( .A(\UART_RXFF/iFIFOMem[2][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1715 ) );
  notech_mux2 \UART_RXFF/U1102  ( .A(\UART_RXFF/iFIFOMem[2][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1716 ) );
  notech_mux2 \UART_RXFF/U1101  ( .A(\UART_RXFF/iFIFOMem[2][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1717 ) );
  notech_mux2 \UART_RXFF/U1100  ( .A(\UART_RXFF/iFIFOMem[2][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1718 ) );
  notech_mux2 \UART_RXFF/U1099  ( .A(\UART_RXFF/iFIFOMem[2][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1719 ) );
  notech_mux2 \UART_RXFF/U1098  ( .A(\UART_RXFF/iFIFOMem[2][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1720 ) );
  notech_mux2 \UART_RXFF/U1097  ( .A(\UART_RXFF/iFIFOMem[2][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1721 ) );
  notech_mux2 \UART_RXFF/U1096  ( .A(\UART_RXFF/iFIFOMem[2][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1722 ) );
  notech_mux2 \UART_RXFF/U1095  ( .A(\UART_RXFF/iFIFOMem[2][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n401 ), .Z(\UART_RXFF/n1723 ) );
  notech_and3 \UART_RXFF/U1094  ( .A(\UART_RXFF/iWRAddr[0] ), .B(
        \UART_RXFF/iWRAddr[1] ), .C(\UART_RXFF/n300 ), .Z(\UART_RXFF/n330 ) );
  notech_and2 \UART_RXFF/U1093  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n400 ) );
  notech_mux2 \UART_RXFF/U1092  ( .A(\UART_RXFF/iFIFOMem[3][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1724 ) );
  notech_mux2 \UART_RXFF/U1091  ( .A(\UART_RXFF/iFIFOMem[3][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1725 ) );
  notech_mux2 \UART_RXFF/U1090  ( .A(\UART_RXFF/iFIFOMem[3][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1726 ) );
  notech_mux2 \UART_RXFF/U1089  ( .A(\UART_RXFF/iFIFOMem[3][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1727 ) );
  notech_mux2 \UART_RXFF/U1088  ( .A(\UART_RXFF/iFIFOMem[3][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1728 ) );
  notech_mux2 \UART_RXFF/U1087  ( .A(\UART_RXFF/iFIFOMem[3][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1729 ) );
  notech_mux2 \UART_RXFF/U1086  ( .A(\UART_RXFF/iFIFOMem[3][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1730 ) );
  notech_mux2 \UART_RXFF/U1085  ( .A(\UART_RXFF/iFIFOMem[3][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1731 ) );
  notech_mux2 \UART_RXFF/U1084  ( .A(\UART_RXFF/iFIFOMem[3][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1732 ) );
  notech_mux2 \UART_RXFF/U1083  ( .A(\UART_RXFF/iFIFOMem[3][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1733 ) );
  notech_mux2 \UART_RXFF/U1082  ( .A(\UART_RXFF/iFIFOMem[3][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n400 ), .Z(\UART_RXFF/n1734 ) );
  notech_and3 \UART_RXFF/U1081  ( .A(\UART_RXFF/iWRAddr[2] ), .B(
        \UART_RXFF/n298 ), .C(\UART_RXFF/n397 ), .Z(\UART_RXFF/n328 ) );
  notech_and2 \UART_RXFF/U1080  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n399 ) );
  notech_mux2 \UART_RXFF/U1079  ( .A(\UART_RXFF/iFIFOMem[4][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1735 ) );
  notech_mux2 \UART_RXFF/U1078  ( .A(\UART_RXFF/iFIFOMem[4][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1736 ) );
  notech_mux2 \UART_RXFF/U1077  ( .A(\UART_RXFF/iFIFOMem[4][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1737 ) );
  notech_mux2 \UART_RXFF/U1076  ( .A(\UART_RXFF/iFIFOMem[4][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1738 ) );
  notech_mux2 \UART_RXFF/U1075  ( .A(\UART_RXFF/iFIFOMem[4][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1739 ) );
  notech_mux2 \UART_RXFF/U1074  ( .A(\UART_RXFF/iFIFOMem[4][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1740 ) );
  notech_mux2 \UART_RXFF/U1073  ( .A(\UART_RXFF/iFIFOMem[4][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1741 ) );
  notech_mux2 \UART_RXFF/U1072  ( .A(\UART_RXFF/iFIFOMem[4][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1742 ) );
  notech_mux2 \UART_RXFF/U1071  ( .A(\UART_RXFF/iFIFOMem[4][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1743 ) );
  notech_mux2 \UART_RXFF/U1070  ( .A(\UART_RXFF/iFIFOMem[4][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1744 ) );
  notech_mux2 \UART_RXFF/U1069  ( .A(\UART_RXFF/iFIFOMem[4][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n399 ), .Z(\UART_RXFF/n1745 ) );
  notech_and3 \UART_RXFF/U1068  ( .A(\UART_RXFF/iWRAddr[0] ), .B(
        \UART_RXFF/iWRAddr[2] ), .C(\UART_RXFF/n298 ), .Z(\UART_RXFF/n326 ) );
  notech_and2 \UART_RXFF/U1067  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n398 ) );
  notech_mux2 \UART_RXFF/U1066  ( .A(\UART_RXFF/iFIFOMem[5][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1746 ) );
  notech_mux2 \UART_RXFF/U1065  ( .A(\UART_RXFF/iFIFOMem[5][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1747 ) );
  notech_mux2 \UART_RXFF/U1064  ( .A(\UART_RXFF/iFIFOMem[5][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1748 ) );
  notech_mux2 \UART_RXFF/U1063  ( .A(\UART_RXFF/iFIFOMem[5][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1749 ) );
  notech_mux2 \UART_RXFF/U1062  ( .A(\UART_RXFF/iFIFOMem[5][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1750 ) );
  notech_mux2 \UART_RXFF/U1061  ( .A(\UART_RXFF/iFIFOMem[5][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1751 ) );
  notech_mux2 \UART_RXFF/U1060  ( .A(\UART_RXFF/iFIFOMem[5][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1752 ) );
  notech_mux2 \UART_RXFF/U1059  ( .A(\UART_RXFF/iFIFOMem[5][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1753 ) );
  notech_mux2 \UART_RXFF/U1058  ( .A(\UART_RXFF/iFIFOMem[5][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1754 ) );
  notech_mux2 \UART_RXFF/U1057  ( .A(\UART_RXFF/iFIFOMem[5][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1755 ) );
  notech_mux2 \UART_RXFF/U1056  ( .A(\UART_RXFF/iFIFOMem[5][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n398 ), .Z(\UART_RXFF/n1756 ) );
  notech_and3 \UART_RXFF/U1055  ( .A(\UART_RXFF/iWRAddr[1] ), .B(
        \UART_RXFF/iWRAddr[2] ), .C(\UART_RXFF/n397 ), .Z(\UART_RXFF/n324 ) );
  notech_and2 \UART_RXFF/U1054  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n396 ) );
  notech_mux2 \UART_RXFF/U1053  ( .A(\UART_RXFF/iFIFOMem[6][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1757 ) );
  notech_mux2 \UART_RXFF/U1052  ( .A(\UART_RXFF/iFIFOMem[6][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1758 ) );
  notech_mux2 \UART_RXFF/U1051  ( .A(\UART_RXFF/iFIFOMem[6][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1759 ) );
  notech_mux2 \UART_RXFF/U1050  ( .A(\UART_RXFF/iFIFOMem[6][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1760 ) );
  notech_mux2 \UART_RXFF/U1049  ( .A(\UART_RXFF/iFIFOMem[6][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1761 ) );
  notech_mux2 \UART_RXFF/U1048  ( .A(\UART_RXFF/iFIFOMem[6][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1762 ) );
  notech_mux2 \UART_RXFF/U1047  ( .A(\UART_RXFF/iFIFOMem[6][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1763 ) );
  notech_mux2 \UART_RXFF/U1046  ( .A(\UART_RXFF/iFIFOMem[6][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1764 ) );
  notech_mux2 \UART_RXFF/U1045  ( .A(\UART_RXFF/iFIFOMem[6][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1765 ) );
  notech_mux2 \UART_RXFF/U1044  ( .A(\UART_RXFF/iFIFOMem[6][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1766 ) );
  notech_mux2 \UART_RXFF/U1043  ( .A(\UART_RXFF/iFIFOMem[6][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n396 ), .Z(\UART_RXFF/n1767 ) );
  notech_and3 \UART_RXFF/U1042  ( .A(\UART_RXFF/iWRAddr[0] ), .B(
        \UART_RXFF/iWRAddr[2] ), .C(\UART_RXFF/iWRAddr[1] ), .Z(
        \UART_RXFF/n322 ) );
  notech_and2 \UART_RXFF/U1041  ( .A(\UART_RXFF/n395 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n394 ) );
  notech_mux2 \UART_RXFF/U1040  ( .A(\UART_RXFF/iFIFOMem[7][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1768 ) );
  notech_mux2 \UART_RXFF/U1039  ( .A(\UART_RXFF/iFIFOMem[7][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1769 ) );
  notech_mux2 \UART_RXFF/U1038  ( .A(\UART_RXFF/iFIFOMem[7][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1770 ) );
  notech_mux2 \UART_RXFF/U1037  ( .A(\UART_RXFF/iFIFOMem[7][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1771 ) );
  notech_mux2 \UART_RXFF/U1036  ( .A(\UART_RXFF/iFIFOMem[7][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1772 ) );
  notech_mux2 \UART_RXFF/U1035  ( .A(\UART_RXFF/iFIFOMem[7][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1773 ) );
  notech_mux2 \UART_RXFF/U1034  ( .A(\UART_RXFF/iFIFOMem[7][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1774 ) );
  notech_mux2 \UART_RXFF/U1033  ( .A(\UART_RXFF/iFIFOMem[7][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1775 ) );
  notech_mux2 \UART_RXFF/U1032  ( .A(\UART_RXFF/iFIFOMem[7][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1776 ) );
  notech_mux2 \UART_RXFF/U1031  ( .A(\UART_RXFF/iFIFOMem[7][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1777 ) );
  notech_mux2 \UART_RXFF/U1030  ( .A(\UART_RXFF/iFIFOMem[7][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n394 ), .Z(\UART_RXFF/n1778 ) );
  notech_ao3 \UART_RXFF/U1029  ( .A(\UART_RXFF/iWRAddr[3] ), .B(
        \UART_RXFF/n375 ), .C(\UART_RXFF/iWRAddr[4] ), .Z(\UART_RXFF/n386 ) );
  notech_and2 \UART_RXFF/U1028  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n393 ) );
  notech_mux2 \UART_RXFF/U1027  ( .A(\UART_RXFF/iFIFOMem[8][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1779 ) );
  notech_mux2 \UART_RXFF/U1026  ( .A(\UART_RXFF/iFIFOMem[8][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1780 ) );
  notech_mux2 \UART_RXFF/U1025  ( .A(\UART_RXFF/iFIFOMem[8][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1781 ) );
  notech_mux2 \UART_RXFF/U1024  ( .A(\UART_RXFF/iFIFOMem[8][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1782 ) );
  notech_mux2 \UART_RXFF/U1023  ( .A(\UART_RXFF/iFIFOMem[8][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1783 ) );
  notech_mux2 \UART_RXFF/U1022  ( .A(\UART_RXFF/iFIFOMem[8][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1784 ) );
  notech_mux2 \UART_RXFF/U1021  ( .A(\UART_RXFF/iFIFOMem[8][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1785 ) );
  notech_mux2 \UART_RXFF/U1020  ( .A(\UART_RXFF/iFIFOMem[8][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1786 ) );
  notech_mux2 \UART_RXFF/U1019  ( .A(\UART_RXFF/iFIFOMem[8][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1787 ) );
  notech_mux2 \UART_RXFF/U1018  ( .A(\UART_RXFF/iFIFOMem[8][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1788 ) );
  notech_mux2 \UART_RXFF/U1017  ( .A(\UART_RXFF/iFIFOMem[8][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n393 ), .Z(\UART_RXFF/n1789 ) );
  notech_and2 \UART_RXFF/U1016  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n392 ) );
  notech_mux2 \UART_RXFF/U1015  ( .A(\UART_RXFF/iFIFOMem[9][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1790 ) );
  notech_mux2 \UART_RXFF/U1014  ( .A(\UART_RXFF/iFIFOMem[9][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1791 ) );
  notech_mux2 \UART_RXFF/U1013  ( .A(\UART_RXFF/iFIFOMem[9][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1792 ) );
  notech_mux2 \UART_RXFF/U1012  ( .A(\UART_RXFF/iFIFOMem[9][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1793 ) );
  notech_mux2 \UART_RXFF/U1011  ( .A(\UART_RXFF/iFIFOMem[9][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1794 ) );
  notech_mux2 \UART_RXFF/U1010  ( .A(\UART_RXFF/iFIFOMem[9][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1795 ) );
  notech_mux2 \UART_RXFF/U1009  ( .A(\UART_RXFF/iFIFOMem[9][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1796 ) );
  notech_mux2 \UART_RXFF/U1008  ( .A(\UART_RXFF/iFIFOMem[9][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1797 ) );
  notech_mux2 \UART_RXFF/U1007  ( .A(\UART_RXFF/iFIFOMem[9][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1798 ) );
  notech_mux2 \UART_RXFF/U1006  ( .A(\UART_RXFF/iFIFOMem[9][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1799 ) );
  notech_mux2 \UART_RXFF/U1005  ( .A(\UART_RXFF/iFIFOMem[9][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n392 ), .Z(\UART_RXFF/n1800 ) );
  notech_and2 \UART_RXFF/U1004  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n391 ) );
  notech_mux2 \UART_RXFF/U1003  ( .A(\UART_RXFF/iFIFOMem[10][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1801 ) );
  notech_mux2 \UART_RXFF/U1002  ( .A(\UART_RXFF/iFIFOMem[10][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1802 ) );
  notech_mux2 \UART_RXFF/U1001  ( .A(\UART_RXFF/iFIFOMem[10][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1803 ) );
  notech_mux2 \UART_RXFF/U1000  ( .A(\UART_RXFF/iFIFOMem[10][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1804 ) );
  notech_mux2 \UART_RXFF/U999  ( .A(\UART_RXFF/iFIFOMem[10][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1805 ) );
  notech_mux2 \UART_RXFF/U998  ( .A(\UART_RXFF/iFIFOMem[10][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1806 ) );
  notech_mux2 \UART_RXFF/U997  ( .A(\UART_RXFF/iFIFOMem[10][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1807 ) );
  notech_mux2 \UART_RXFF/U996  ( .A(\UART_RXFF/iFIFOMem[10][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1808 ) );
  notech_mux2 \UART_RXFF/U995  ( .A(\UART_RXFF/iFIFOMem[10][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1809 ) );
  notech_mux2 \UART_RXFF/U994  ( .A(\UART_RXFF/iFIFOMem[10][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1810 ) );
  notech_mux2 \UART_RXFF/U993  ( .A(\UART_RXFF/iFIFOMem[10][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n391 ), .Z(\UART_RXFF/n1811 ) );
  notech_and2 \UART_RXFF/U992  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n390 ) );
  notech_mux2 \UART_RXFF/U991  ( .A(\UART_RXFF/iFIFOMem[11][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1812 ) );
  notech_mux2 \UART_RXFF/U990  ( .A(\UART_RXFF/iFIFOMem[11][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1813 ) );
  notech_mux2 \UART_RXFF/U989  ( .A(\UART_RXFF/iFIFOMem[11][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1814 ) );
  notech_mux2 \UART_RXFF/U988  ( .A(\UART_RXFF/iFIFOMem[11][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1815 ) );
  notech_mux2 \UART_RXFF/U987  ( .A(\UART_RXFF/iFIFOMem[11][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1816 ) );
  notech_mux2 \UART_RXFF/U986  ( .A(\UART_RXFF/iFIFOMem[11][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1817 ) );
  notech_mux2 \UART_RXFF/U985  ( .A(\UART_RXFF/iFIFOMem[11][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1818 ) );
  notech_mux2 \UART_RXFF/U984  ( .A(\UART_RXFF/iFIFOMem[11][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1819 ) );
  notech_mux2 \UART_RXFF/U983  ( .A(\UART_RXFF/iFIFOMem[11][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1820 ) );
  notech_mux2 \UART_RXFF/U982  ( .A(\UART_RXFF/iFIFOMem[11][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1821 ) );
  notech_mux2 \UART_RXFF/U981  ( .A(\UART_RXFF/iFIFOMem[11][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n390 ), .Z(\UART_RXFF/n1822 ) );
  notech_and2 \UART_RXFF/U980  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n389 ) );
  notech_mux2 \UART_RXFF/U979  ( .A(\UART_RXFF/iFIFOMem[12][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1823 ) );
  notech_mux2 \UART_RXFF/U978  ( .A(\UART_RXFF/iFIFOMem[12][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1824 ) );
  notech_mux2 \UART_RXFF/U977  ( .A(\UART_RXFF/iFIFOMem[12][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1825 ) );
  notech_mux2 \UART_RXFF/U976  ( .A(\UART_RXFF/iFIFOMem[12][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1826 ) );
  notech_mux2 \UART_RXFF/U975  ( .A(\UART_RXFF/iFIFOMem[12][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1827 ) );
  notech_mux2 \UART_RXFF/U974  ( .A(\UART_RXFF/iFIFOMem[12][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1828 ) );
  notech_mux2 \UART_RXFF/U973  ( .A(\UART_RXFF/iFIFOMem[12][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1829 ) );
  notech_mux2 \UART_RXFF/U972  ( .A(\UART_RXFF/iFIFOMem[12][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1830 ) );
  notech_mux2 \UART_RXFF/U971  ( .A(\UART_RXFF/iFIFOMem[12][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1831 ) );
  notech_mux2 \UART_RXFF/U970  ( .A(\UART_RXFF/iFIFOMem[12][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1832 ) );
  notech_mux2 \UART_RXFF/U969  ( .A(\UART_RXFF/iFIFOMem[12][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n389 ), .Z(\UART_RXFF/n1833 ) );
  notech_and2 \UART_RXFF/U968  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n388 ) );
  notech_mux2 \UART_RXFF/U967  ( .A(\UART_RXFF/iFIFOMem[13][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1834 ) );
  notech_mux2 \UART_RXFF/U966  ( .A(\UART_RXFF/iFIFOMem[13][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1835 ) );
  notech_mux2 \UART_RXFF/U965  ( .A(\UART_RXFF/iFIFOMem[13][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1836 ) );
  notech_mux2 \UART_RXFF/U964  ( .A(\UART_RXFF/iFIFOMem[13][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1837 ) );
  notech_mux2 \UART_RXFF/U963  ( .A(\UART_RXFF/iFIFOMem[13][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1838 ) );
  notech_mux2 \UART_RXFF/U962  ( .A(\UART_RXFF/iFIFOMem[13][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1839 ) );
  notech_mux2 \UART_RXFF/U961  ( .A(\UART_RXFF/iFIFOMem[13][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1840 ) );
  notech_mux2 \UART_RXFF/U960  ( .A(\UART_RXFF/iFIFOMem[13][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1841 ) );
  notech_mux2 \UART_RXFF/U959  ( .A(\UART_RXFF/iFIFOMem[13][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1842 ) );
  notech_mux2 \UART_RXFF/U958  ( .A(\UART_RXFF/iFIFOMem[13][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1843 ) );
  notech_mux2 \UART_RXFF/U957  ( .A(\UART_RXFF/iFIFOMem[13][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n388 ), .Z(\UART_RXFF/n1844 ) );
  notech_and2 \UART_RXFF/U956  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n387 ) );
  notech_mux2 \UART_RXFF/U955  ( .A(\UART_RXFF/iFIFOMem[14][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1845 ) );
  notech_mux2 \UART_RXFF/U954  ( .A(\UART_RXFF/iFIFOMem[14][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1846 ) );
  notech_mux2 \UART_RXFF/U953  ( .A(\UART_RXFF/iFIFOMem[14][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1847 ) );
  notech_mux2 \UART_RXFF/U952  ( .A(\UART_RXFF/iFIFOMem[14][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1848 ) );
  notech_mux2 \UART_RXFF/U951  ( .A(\UART_RXFF/iFIFOMem[14][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1849 ) );
  notech_mux2 \UART_RXFF/U950  ( .A(\UART_RXFF/iFIFOMem[14][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1850 ) );
  notech_mux2 \UART_RXFF/U949  ( .A(\UART_RXFF/iFIFOMem[14][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1851 ) );
  notech_mux2 \UART_RXFF/U948  ( .A(\UART_RXFF/iFIFOMem[14][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1852 ) );
  notech_mux2 \UART_RXFF/U947  ( .A(\UART_RXFF/iFIFOMem[14][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1853 ) );
  notech_mux2 \UART_RXFF/U946  ( .A(\UART_RXFF/iFIFOMem[14][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1854 ) );
  notech_mux2 \UART_RXFF/U945  ( .A(\UART_RXFF/iFIFOMem[14][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n387 ), .Z(\UART_RXFF/n1855 ) );
  notech_and2 \UART_RXFF/U944  ( .A(\UART_RXFF/n386 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n385 ) );
  notech_mux2 \UART_RXFF/U943  ( .A(\UART_RXFF/iFIFOMem[15][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1856 ) );
  notech_mux2 \UART_RXFF/U942  ( .A(\UART_RXFF/iFIFOMem[15][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1857 ) );
  notech_mux2 \UART_RXFF/U941  ( .A(\UART_RXFF/iFIFOMem[15][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1858 ) );
  notech_mux2 \UART_RXFF/U940  ( .A(\UART_RXFF/iFIFOMem[15][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1859 ) );
  notech_mux2 \UART_RXFF/U939  ( .A(\UART_RXFF/iFIFOMem[15][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1860 ) );
  notech_mux2 \UART_RXFF/U938  ( .A(\UART_RXFF/iFIFOMem[15][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1861 ) );
  notech_mux2 \UART_RXFF/U937  ( .A(\UART_RXFF/iFIFOMem[15][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1862 ) );
  notech_mux2 \UART_RXFF/U936  ( .A(\UART_RXFF/iFIFOMem[15][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1863 ) );
  notech_mux2 \UART_RXFF/U935  ( .A(\UART_RXFF/iFIFOMem[15][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1864 ) );
  notech_mux2 \UART_RXFF/U934  ( .A(\UART_RXFF/iFIFOMem[15][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1865 ) );
  notech_mux2 \UART_RXFF/U933  ( .A(\UART_RXFF/iFIFOMem[15][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n385 ), .Z(\UART_RXFF/n1866 ) );
  notech_ao3 \UART_RXFF/U932  ( .A(\UART_RXFF/iWRAddr[4] ), .B(
        \UART_RXFF/n375 ), .C(\UART_RXFF/iWRAddr[3] ), .Z(\UART_RXFF/n377 ) );
  notech_and2 \UART_RXFF/U931  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n384 ) );
  notech_mux2 \UART_RXFF/U930  ( .A(\UART_RXFF/iFIFOMem[16][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1867 ) );
  notech_mux2 \UART_RXFF/U929  ( .A(\UART_RXFF/iFIFOMem[16][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1868 ) );
  notech_mux2 \UART_RXFF/U928  ( .A(\UART_RXFF/iFIFOMem[16][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1869 ) );
  notech_mux2 \UART_RXFF/U927  ( .A(\UART_RXFF/iFIFOMem[16][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1870 ) );
  notech_mux2 \UART_RXFF/U926  ( .A(\UART_RXFF/iFIFOMem[16][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1871 ) );
  notech_mux2 \UART_RXFF/U925  ( .A(\UART_RXFF/iFIFOMem[16][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1872 ) );
  notech_mux2 \UART_RXFF/U924  ( .A(\UART_RXFF/iFIFOMem[16][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1873 ) );
  notech_mux2 \UART_RXFF/U923  ( .A(\UART_RXFF/iFIFOMem[16][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1874 ) );
  notech_mux2 \UART_RXFF/U922  ( .A(\UART_RXFF/iFIFOMem[16][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1875 ) );
  notech_mux2 \UART_RXFF/U921  ( .A(\UART_RXFF/iFIFOMem[16][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1876 ) );
  notech_mux2 \UART_RXFF/U920  ( .A(\UART_RXFF/iFIFOMem[16][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n384 ), .Z(\UART_RXFF/n1877 ) );
  notech_and2 \UART_RXFF/U919  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n383 ) );
  notech_mux2 \UART_RXFF/U918  ( .A(\UART_RXFF/iFIFOMem[17][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1878 ) );
  notech_mux2 \UART_RXFF/U917  ( .A(\UART_RXFF/iFIFOMem[17][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1879 ) );
  notech_mux2 \UART_RXFF/U916  ( .A(\UART_RXFF/iFIFOMem[17][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1880 ) );
  notech_mux2 \UART_RXFF/U915  ( .A(\UART_RXFF/iFIFOMem[17][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1881 ) );
  notech_mux2 \UART_RXFF/U914  ( .A(\UART_RXFF/iFIFOMem[17][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1882 ) );
  notech_mux2 \UART_RXFF/U913  ( .A(\UART_RXFF/iFIFOMem[17][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1883 ) );
  notech_mux2 \UART_RXFF/U912  ( .A(\UART_RXFF/iFIFOMem[17][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1884 ) );
  notech_mux2 \UART_RXFF/U911  ( .A(\UART_RXFF/iFIFOMem[17][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1885 ) );
  notech_mux2 \UART_RXFF/U910  ( .A(\UART_RXFF/iFIFOMem[17][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1886 ) );
  notech_mux2 \UART_RXFF/U909  ( .A(\UART_RXFF/iFIFOMem[17][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1887 ) );
  notech_mux2 \UART_RXFF/U908  ( .A(\UART_RXFF/iFIFOMem[17][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n383 ), .Z(\UART_RXFF/n1888 ) );
  notech_and2 \UART_RXFF/U907  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n382 ) );
  notech_mux2 \UART_RXFF/U906  ( .A(\UART_RXFF/iFIFOMem[18][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1889 ) );
  notech_mux2 \UART_RXFF/U905  ( .A(\UART_RXFF/iFIFOMem[18][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1890 ) );
  notech_mux2 \UART_RXFF/U904  ( .A(\UART_RXFF/iFIFOMem[18][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1891 ) );
  notech_mux2 \UART_RXFF/U903  ( .A(\UART_RXFF/iFIFOMem[18][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1892 ) );
  notech_mux2 \UART_RXFF/U902  ( .A(\UART_RXFF/iFIFOMem[18][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1893 ) );
  notech_mux2 \UART_RXFF/U901  ( .A(\UART_RXFF/iFIFOMem[18][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1894 ) );
  notech_mux2 \UART_RXFF/U900  ( .A(\UART_RXFF/iFIFOMem[18][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1895 ) );
  notech_mux2 \UART_RXFF/U899  ( .A(\UART_RXFF/iFIFOMem[18][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1896 ) );
  notech_mux2 \UART_RXFF/U898  ( .A(\UART_RXFF/iFIFOMem[18][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1897 ) );
  notech_mux2 \UART_RXFF/U897  ( .A(\UART_RXFF/iFIFOMem[18][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1898 ) );
  notech_mux2 \UART_RXFF/U896  ( .A(\UART_RXFF/iFIFOMem[18][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n382 ), .Z(\UART_RXFF/n1899 ) );
  notech_and2 \UART_RXFF/U895  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n381 ) );
  notech_mux2 \UART_RXFF/U894  ( .A(\UART_RXFF/iFIFOMem[19][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1900 ) );
  notech_mux2 \UART_RXFF/U893  ( .A(\UART_RXFF/iFIFOMem[19][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1901 ) );
  notech_mux2 \UART_RXFF/U892  ( .A(\UART_RXFF/iFIFOMem[19][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1902 ) );
  notech_mux2 \UART_RXFF/U891  ( .A(\UART_RXFF/iFIFOMem[19][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1903 ) );
  notech_mux2 \UART_RXFF/U890  ( .A(\UART_RXFF/iFIFOMem[19][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1904 ) );
  notech_mux2 \UART_RXFF/U889  ( .A(\UART_RXFF/iFIFOMem[19][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1905 ) );
  notech_mux2 \UART_RXFF/U888  ( .A(\UART_RXFF/iFIFOMem[19][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1906 ) );
  notech_mux2 \UART_RXFF/U887  ( .A(\UART_RXFF/iFIFOMem[19][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1907 ) );
  notech_mux2 \UART_RXFF/U886  ( .A(\UART_RXFF/iFIFOMem[19][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1908 ) );
  notech_mux2 \UART_RXFF/U885  ( .A(\UART_RXFF/iFIFOMem[19][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1909 ) );
  notech_mux2 \UART_RXFF/U884  ( .A(\UART_RXFF/iFIFOMem[19][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n381 ), .Z(\UART_RXFF/n1910 ) );
  notech_and2 \UART_RXFF/U883  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n380 ) );
  notech_mux2 \UART_RXFF/U882  ( .A(\UART_RXFF/iFIFOMem[20][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1911 ) );
  notech_mux2 \UART_RXFF/U881  ( .A(\UART_RXFF/iFIFOMem[20][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1912 ) );
  notech_mux2 \UART_RXFF/U880  ( .A(\UART_RXFF/iFIFOMem[20][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1913 ) );
  notech_mux2 \UART_RXFF/U879  ( .A(\UART_RXFF/iFIFOMem[20][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1914 ) );
  notech_mux2 \UART_RXFF/U878  ( .A(\UART_RXFF/iFIFOMem[20][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1915 ) );
  notech_mux2 \UART_RXFF/U877  ( .A(\UART_RXFF/iFIFOMem[20][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1916 ) );
  notech_mux2 \UART_RXFF/U876  ( .A(\UART_RXFF/iFIFOMem[20][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1917 ) );
  notech_mux2 \UART_RXFF/U875  ( .A(\UART_RXFF/iFIFOMem[20][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1918 ) );
  notech_mux2 \UART_RXFF/U874  ( .A(\UART_RXFF/iFIFOMem[20][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1919 ) );
  notech_mux2 \UART_RXFF/U873  ( .A(\UART_RXFF/iFIFOMem[20][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1920 ) );
  notech_mux2 \UART_RXFF/U872  ( .A(\UART_RXFF/iFIFOMem[20][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n380 ), .Z(\UART_RXFF/n1921 ) );
  notech_and2 \UART_RXFF/U871  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n379 ) );
  notech_mux2 \UART_RXFF/U870  ( .A(\UART_RXFF/iFIFOMem[21][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1922 ) );
  notech_mux2 \UART_RXFF/U869  ( .A(\UART_RXFF/iFIFOMem[21][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1923 ) );
  notech_mux2 \UART_RXFF/U868  ( .A(\UART_RXFF/iFIFOMem[21][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1924 ) );
  notech_mux2 \UART_RXFF/U867  ( .A(\UART_RXFF/iFIFOMem[21][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1925 ) );
  notech_mux2 \UART_RXFF/U866  ( .A(\UART_RXFF/iFIFOMem[21][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1926 ) );
  notech_mux2 \UART_RXFF/U865  ( .A(\UART_RXFF/iFIFOMem[21][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1927 ) );
  notech_mux2 \UART_RXFF/U864  ( .A(\UART_RXFF/iFIFOMem[21][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1928 ) );
  notech_mux2 \UART_RXFF/U863  ( .A(\UART_RXFF/iFIFOMem[21][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1929 ) );
  notech_mux2 \UART_RXFF/U862  ( .A(\UART_RXFF/iFIFOMem[21][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1930 ) );
  notech_mux2 \UART_RXFF/U861  ( .A(\UART_RXFF/iFIFOMem[21][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1931 ) );
  notech_mux2 \UART_RXFF/U860  ( .A(\UART_RXFF/iFIFOMem[21][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n379 ), .Z(\UART_RXFF/n1932 ) );
  notech_and2 \UART_RXFF/U859  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n378 ) );
  notech_mux2 \UART_RXFF/U858  ( .A(\UART_RXFF/iFIFOMem[22][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1933 ) );
  notech_mux2 \UART_RXFF/U857  ( .A(\UART_RXFF/iFIFOMem[22][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1934 ) );
  notech_mux2 \UART_RXFF/U856  ( .A(\UART_RXFF/iFIFOMem[22][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1935 ) );
  notech_mux2 \UART_RXFF/U855  ( .A(\UART_RXFF/iFIFOMem[22][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1936 ) );
  notech_mux2 \UART_RXFF/U854  ( .A(\UART_RXFF/iFIFOMem[22][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1937 ) );
  notech_mux2 \UART_RXFF/U853  ( .A(\UART_RXFF/iFIFOMem[22][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1938 ) );
  notech_mux2 \UART_RXFF/U852  ( .A(\UART_RXFF/iFIFOMem[22][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1939 ) );
  notech_mux2 \UART_RXFF/U851  ( .A(\UART_RXFF/iFIFOMem[22][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1940 ) );
  notech_mux2 \UART_RXFF/U850  ( .A(\UART_RXFF/iFIFOMem[22][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1941 ) );
  notech_mux2 \UART_RXFF/U849  ( .A(\UART_RXFF/iFIFOMem[22][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1942 ) );
  notech_mux2 \UART_RXFF/U848  ( .A(\UART_RXFF/iFIFOMem[22][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n378 ), .Z(\UART_RXFF/n1943 ) );
  notech_and2 \UART_RXFF/U847  ( .A(\UART_RXFF/n377 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n376 ) );
  notech_mux2 \UART_RXFF/U846  ( .A(\UART_RXFF/iFIFOMem[23][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1944 ) );
  notech_mux2 \UART_RXFF/U845  ( .A(\UART_RXFF/iFIFOMem[23][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1945 ) );
  notech_mux2 \UART_RXFF/U844  ( .A(\UART_RXFF/iFIFOMem[23][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1946 ) );
  notech_mux2 \UART_RXFF/U843  ( .A(\UART_RXFF/iFIFOMem[23][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1947 ) );
  notech_mux2 \UART_RXFF/U842  ( .A(\UART_RXFF/iFIFOMem[23][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1948 ) );
  notech_mux2 \UART_RXFF/U841  ( .A(\UART_RXFF/iFIFOMem[23][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1949 ) );
  notech_mux2 \UART_RXFF/U840  ( .A(\UART_RXFF/iFIFOMem[23][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1950 ) );
  notech_mux2 \UART_RXFF/U839  ( .A(\UART_RXFF/iFIFOMem[23][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1951 ) );
  notech_mux2 \UART_RXFF/U838  ( .A(\UART_RXFF/iFIFOMem[23][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1952 ) );
  notech_mux2 \UART_RXFF/U837  ( .A(\UART_RXFF/iFIFOMem[23][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1953 ) );
  notech_mux2 \UART_RXFF/U836  ( .A(\UART_RXFF/iFIFOMem[23][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n376 ), .Z(\UART_RXFF/n1954 ) );
  notech_ao3 \UART_RXFF/U835  ( .A(\UART_RXFF/iWRAddr[4] ), .B(
        \UART_RXFF/n375 ), .C(\UART_RXFF/n302 ), .Z(\UART_RXFF/n367 ) );
  notech_and2 \UART_RXFF/U834  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n374 ) );
  notech_mux2 \UART_RXFF/U833  ( .A(\UART_RXFF/iFIFOMem[24][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1955 ) );
  notech_mux2 \UART_RXFF/U832  ( .A(\UART_RXFF/iFIFOMem[24][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1956 ) );
  notech_mux2 \UART_RXFF/U831  ( .A(\UART_RXFF/iFIFOMem[24][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1957 ) );
  notech_mux2 \UART_RXFF/U830  ( .A(\UART_RXFF/iFIFOMem[24][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1958 ) );
  notech_mux2 \UART_RXFF/U829  ( .A(\UART_RXFF/iFIFOMem[24][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1959 ) );
  notech_mux2 \UART_RXFF/U828  ( .A(\UART_RXFF/iFIFOMem[24][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1960 ) );
  notech_mux2 \UART_RXFF/U827  ( .A(\UART_RXFF/iFIFOMem[24][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1961 ) );
  notech_mux2 \UART_RXFF/U826  ( .A(\UART_RXFF/iFIFOMem[24][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1962 ) );
  notech_mux2 \UART_RXFF/U825  ( .A(\UART_RXFF/iFIFOMem[24][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1963 ) );
  notech_mux2 \UART_RXFF/U824  ( .A(\UART_RXFF/iFIFOMem[24][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1964 ) );
  notech_mux2 \UART_RXFF/U823  ( .A(\UART_RXFF/iFIFOMem[24][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n374 ), .Z(\UART_RXFF/n1965 ) );
  notech_and2 \UART_RXFF/U822  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n373 ) );
  notech_mux2 \UART_RXFF/U821  ( .A(\UART_RXFF/iFIFOMem[25][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1966 ) );
  notech_mux2 \UART_RXFF/U820  ( .A(\UART_RXFF/iFIFOMem[25][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1967 ) );
  notech_mux2 \UART_RXFF/U819  ( .A(\UART_RXFF/iFIFOMem[25][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1968 ) );
  notech_mux2 \UART_RXFF/U818  ( .A(\UART_RXFF/iFIFOMem[25][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1969 ) );
  notech_mux2 \UART_RXFF/U817  ( .A(\UART_RXFF/iFIFOMem[25][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1970 ) );
  notech_mux2 \UART_RXFF/U816  ( .A(\UART_RXFF/iFIFOMem[25][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1971 ) );
  notech_mux2 \UART_RXFF/U815  ( .A(\UART_RXFF/iFIFOMem[25][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1972 ) );
  notech_mux2 \UART_RXFF/U814  ( .A(\UART_RXFF/iFIFOMem[25][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1973 ) );
  notech_mux2 \UART_RXFF/U813  ( .A(\UART_RXFF/iFIFOMem[25][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1974 ) );
  notech_mux2 \UART_RXFF/U812  ( .A(\UART_RXFF/iFIFOMem[25][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1975 ) );
  notech_mux2 \UART_RXFF/U811  ( .A(\UART_RXFF/iFIFOMem[25][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n373 ), .Z(\UART_RXFF/n1976 ) );
  notech_and2 \UART_RXFF/U810  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n372 ) );
  notech_mux2 \UART_RXFF/U809  ( .A(\UART_RXFF/iFIFOMem[26][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1977 ) );
  notech_mux2 \UART_RXFF/U808  ( .A(\UART_RXFF/iFIFOMem[26][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1978 ) );
  notech_mux2 \UART_RXFF/U807  ( .A(\UART_RXFF/iFIFOMem[26][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1979 ) );
  notech_mux2 \UART_RXFF/U806  ( .A(\UART_RXFF/iFIFOMem[26][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1980 ) );
  notech_mux2 \UART_RXFF/U805  ( .A(\UART_RXFF/iFIFOMem[26][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1981 ) );
  notech_mux2 \UART_RXFF/U804  ( .A(\UART_RXFF/iFIFOMem[26][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1982 ) );
  notech_mux2 \UART_RXFF/U803  ( .A(\UART_RXFF/iFIFOMem[26][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1983 ) );
  notech_mux2 \UART_RXFF/U802  ( .A(\UART_RXFF/iFIFOMem[26][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1984 ) );
  notech_mux2 \UART_RXFF/U801  ( .A(\UART_RXFF/iFIFOMem[26][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1985 ) );
  notech_mux2 \UART_RXFF/U800  ( .A(\UART_RXFF/iFIFOMem[26][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1986 ) );
  notech_mux2 \UART_RXFF/U799  ( .A(\UART_RXFF/iFIFOMem[26][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n372 ), .Z(\UART_RXFF/n1987 ) );
  notech_and2 \UART_RXFF/U798  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n371 ) );
  notech_mux2 \UART_RXFF/U797  ( .A(\UART_RXFF/iFIFOMem[27][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1988 ) );
  notech_mux2 \UART_RXFF/U796  ( .A(\UART_RXFF/iFIFOMem[27][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1989 ) );
  notech_mux2 \UART_RXFF/U795  ( .A(\UART_RXFF/iFIFOMem[27][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1990 ) );
  notech_mux2 \UART_RXFF/U794  ( .A(\UART_RXFF/iFIFOMem[27][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1991 ) );
  notech_mux2 \UART_RXFF/U793  ( .A(\UART_RXFF/iFIFOMem[27][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1992 ) );
  notech_mux2 \UART_RXFF/U792  ( .A(\UART_RXFF/iFIFOMem[27][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1993 ) );
  notech_mux2 \UART_RXFF/U791  ( .A(\UART_RXFF/iFIFOMem[27][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1994 ) );
  notech_mux2 \UART_RXFF/U790  ( .A(\UART_RXFF/iFIFOMem[27][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1995 ) );
  notech_mux2 \UART_RXFF/U789  ( .A(\UART_RXFF/iFIFOMem[27][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1996 ) );
  notech_mux2 \UART_RXFF/U788  ( .A(\UART_RXFF/iFIFOMem[27][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1997 ) );
  notech_mux2 \UART_RXFF/U787  ( .A(\UART_RXFF/iFIFOMem[27][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n371 ), .Z(\UART_RXFF/n1998 ) );
  notech_and2 \UART_RXFF/U786  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n370 ) );
  notech_mux2 \UART_RXFF/U785  ( .A(\UART_RXFF/iFIFOMem[28][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n1999 ) );
  notech_mux2 \UART_RXFF/U784  ( .A(\UART_RXFF/iFIFOMem[28][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2000 ) );
  notech_mux2 \UART_RXFF/U783  ( .A(\UART_RXFF/iFIFOMem[28][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2001 ) );
  notech_mux2 \UART_RXFF/U782  ( .A(\UART_RXFF/iFIFOMem[28][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2002 ) );
  notech_mux2 \UART_RXFF/U781  ( .A(\UART_RXFF/iFIFOMem[28][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2003 ) );
  notech_mux2 \UART_RXFF/U780  ( .A(\UART_RXFF/iFIFOMem[28][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2004 ) );
  notech_mux2 \UART_RXFF/U779  ( .A(\UART_RXFF/iFIFOMem[28][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2005 ) );
  notech_mux2 \UART_RXFF/U778  ( .A(\UART_RXFF/iFIFOMem[28][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2006 ) );
  notech_mux2 \UART_RXFF/U777  ( .A(\UART_RXFF/iFIFOMem[28][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2007 ) );
  notech_mux2 \UART_RXFF/U776  ( .A(\UART_RXFF/iFIFOMem[28][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2008 ) );
  notech_mux2 \UART_RXFF/U775  ( .A(\UART_RXFF/iFIFOMem[28][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n370 ), .Z(\UART_RXFF/n2009 ) );
  notech_and2 \UART_RXFF/U774  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n369 ) );
  notech_mux2 \UART_RXFF/U773  ( .A(\UART_RXFF/iFIFOMem[29][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2010 ) );
  notech_mux2 \UART_RXFF/U772  ( .A(\UART_RXFF/iFIFOMem[29][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2011 ) );
  notech_mux2 \UART_RXFF/U771  ( .A(\UART_RXFF/iFIFOMem[29][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2012 ) );
  notech_mux2 \UART_RXFF/U770  ( .A(\UART_RXFF/iFIFOMem[29][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2013 ) );
  notech_mux2 \UART_RXFF/U769  ( .A(\UART_RXFF/iFIFOMem[29][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2014 ) );
  notech_mux2 \UART_RXFF/U768  ( .A(\UART_RXFF/iFIFOMem[29][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2015 ) );
  notech_mux2 \UART_RXFF/U767  ( .A(\UART_RXFF/iFIFOMem[29][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2016 ) );
  notech_mux2 \UART_RXFF/U766  ( .A(\UART_RXFF/iFIFOMem[29][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2017 ) );
  notech_mux2 \UART_RXFF/U765  ( .A(\UART_RXFF/iFIFOMem[29][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2018 ) );
  notech_mux2 \UART_RXFF/U764  ( .A(\UART_RXFF/iFIFOMem[29][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2019 ) );
  notech_mux2 \UART_RXFF/U763  ( .A(\UART_RXFF/iFIFOMem[29][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n369 ), .Z(\UART_RXFF/n2020 ) );
  notech_and2 \UART_RXFF/U762  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n368 ) );
  notech_mux2 \UART_RXFF/U761  ( .A(\UART_RXFF/iFIFOMem[30][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2021 ) );
  notech_mux2 \UART_RXFF/U760  ( .A(\UART_RXFF/iFIFOMem[30][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2022 ) );
  notech_mux2 \UART_RXFF/U759  ( .A(\UART_RXFF/iFIFOMem[30][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2023 ) );
  notech_mux2 \UART_RXFF/U758  ( .A(\UART_RXFF/iFIFOMem[30][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2024 ) );
  notech_mux2 \UART_RXFF/U757  ( .A(\UART_RXFF/iFIFOMem[30][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2025 ) );
  notech_mux2 \UART_RXFF/U756  ( .A(\UART_RXFF/iFIFOMem[30][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2026 ) );
  notech_mux2 \UART_RXFF/U755  ( .A(\UART_RXFF/iFIFOMem[30][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2027 ) );
  notech_mux2 \UART_RXFF/U754  ( .A(\UART_RXFF/iFIFOMem[30][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2028 ) );
  notech_mux2 \UART_RXFF/U753  ( .A(\UART_RXFF/iFIFOMem[30][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2029 ) );
  notech_mux2 \UART_RXFF/U752  ( .A(\UART_RXFF/iFIFOMem[30][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2030 ) );
  notech_mux2 \UART_RXFF/U751  ( .A(\UART_RXFF/iFIFOMem[30][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n368 ), .Z(\UART_RXFF/n2031 ) );
  notech_and2 \UART_RXFF/U750  ( .A(\UART_RXFF/n367 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n366 ) );
  notech_mux2 \UART_RXFF/U749  ( .A(\UART_RXFF/iFIFOMem[31][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2032 ) );
  notech_mux2 \UART_RXFF/U748  ( .A(\UART_RXFF/iFIFOMem[31][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2033 ) );
  notech_mux2 \UART_RXFF/U747  ( .A(\UART_RXFF/iFIFOMem[31][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2034 ) );
  notech_mux2 \UART_RXFF/U746  ( .A(\UART_RXFF/iFIFOMem[31][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2035 ) );
  notech_mux2 \UART_RXFF/U745  ( .A(\UART_RXFF/iFIFOMem[31][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2036 ) );
  notech_mux2 \UART_RXFF/U744  ( .A(\UART_RXFF/iFIFOMem[31][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2037 ) );
  notech_mux2 \UART_RXFF/U743  ( .A(\UART_RXFF/iFIFOMem[31][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2038 ) );
  notech_mux2 \UART_RXFF/U742  ( .A(\UART_RXFF/iFIFOMem[31][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2039 ) );
  notech_mux2 \UART_RXFF/U741  ( .A(\UART_RXFF/iFIFOMem[31][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2040 ) );
  notech_mux2 \UART_RXFF/U740  ( .A(\UART_RXFF/iFIFOMem[31][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2041 ) );
  notech_mux2 \UART_RXFF/U739  ( .A(\UART_RXFF/iFIFOMem[31][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n366 ), .Z(\UART_RXFF/n2042 ) );
  notech_ao3 \UART_RXFF/U738  ( .A(\UART_RXFF/iWRAddr[5] ), .B(
        \UART_RXFF/n365 ), .C(RST), .Z(\UART_RXFF/n337 ) );
  notech_ao3 \UART_RXFF/U737  ( .A(\UART_RXFF/n302 ), .B(\UART_RXFF/n337 ), 
        .C(\UART_RXFF/iWRAddr[4] ), .Z(\UART_RXFF/n357 ) );
  notech_and2 \UART_RXFF/U736  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n364 ) );
  notech_mux2 \UART_RXFF/U735  ( .A(\UART_RXFF/iFIFOMem[32][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2043 ) );
  notech_mux2 \UART_RXFF/U734  ( .A(\UART_RXFF/iFIFOMem[32][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2044 ) );
  notech_mux2 \UART_RXFF/U733  ( .A(\UART_RXFF/iFIFOMem[32][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2045 ) );
  notech_mux2 \UART_RXFF/U732  ( .A(\UART_RXFF/iFIFOMem[32][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2046 ) );
  notech_mux2 \UART_RXFF/U731  ( .A(\UART_RXFF/iFIFOMem[32][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2047 ) );
  notech_mux2 \UART_RXFF/U730  ( .A(\UART_RXFF/iFIFOMem[32][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2048 ) );
  notech_mux2 \UART_RXFF/U729  ( .A(\UART_RXFF/iFIFOMem[32][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2049 ) );
  notech_mux2 \UART_RXFF/U728  ( .A(\UART_RXFF/iFIFOMem[32][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2050 ) );
  notech_mux2 \UART_RXFF/U727  ( .A(\UART_RXFF/iFIFOMem[32][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2051 ) );
  notech_mux2 \UART_RXFF/U726  ( .A(\UART_RXFF/iFIFOMem[32][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2052 ) );
  notech_mux2 \UART_RXFF/U725  ( .A(\UART_RXFF/iFIFOMem[32][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n364 ), .Z(\UART_RXFF/n2053 ) );
  notech_and2 \UART_RXFF/U724  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n363 ) );
  notech_mux2 \UART_RXFF/U723  ( .A(\UART_RXFF/iFIFOMem[33][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2054 ) );
  notech_mux2 \UART_RXFF/U722  ( .A(\UART_RXFF/iFIFOMem[33][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2055 ) );
  notech_mux2 \UART_RXFF/U721  ( .A(\UART_RXFF/iFIFOMem[33][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2056 ) );
  notech_mux2 \UART_RXFF/U720  ( .A(\UART_RXFF/iFIFOMem[33][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2057 ) );
  notech_mux2 \UART_RXFF/U719  ( .A(\UART_RXFF/iFIFOMem[33][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2058 ) );
  notech_mux2 \UART_RXFF/U718  ( .A(\UART_RXFF/iFIFOMem[33][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2059 ) );
  notech_mux2 \UART_RXFF/U717  ( .A(\UART_RXFF/iFIFOMem[33][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2060 ) );
  notech_mux2 \UART_RXFF/U716  ( .A(\UART_RXFF/iFIFOMem[33][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2061 ) );
  notech_mux2 \UART_RXFF/U715  ( .A(\UART_RXFF/iFIFOMem[33][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2062 ) );
  notech_mux2 \UART_RXFF/U714  ( .A(\UART_RXFF/iFIFOMem[33][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2063 ) );
  notech_mux2 \UART_RXFF/U713  ( .A(\UART_RXFF/iFIFOMem[33][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n363 ), .Z(\UART_RXFF/n2064 ) );
  notech_and2 \UART_RXFF/U712  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n362 ) );
  notech_mux2 \UART_RXFF/U711  ( .A(\UART_RXFF/iFIFOMem[34][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2065 ) );
  notech_mux2 \UART_RXFF/U710  ( .A(\UART_RXFF/iFIFOMem[34][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2066 ) );
  notech_mux2 \UART_RXFF/U709  ( .A(\UART_RXFF/iFIFOMem[34][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2067 ) );
  notech_mux2 \UART_RXFF/U708  ( .A(\UART_RXFF/iFIFOMem[34][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2068 ) );
  notech_mux2 \UART_RXFF/U707  ( .A(\UART_RXFF/iFIFOMem[34][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2069 ) );
  notech_mux2 \UART_RXFF/U706  ( .A(\UART_RXFF/iFIFOMem[34][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2070 ) );
  notech_mux2 \UART_RXFF/U705  ( .A(\UART_RXFF/iFIFOMem[34][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2071 ) );
  notech_mux2 \UART_RXFF/U704  ( .A(\UART_RXFF/iFIFOMem[34][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2072 ) );
  notech_mux2 \UART_RXFF/U703  ( .A(\UART_RXFF/iFIFOMem[34][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2073 ) );
  notech_mux2 \UART_RXFF/U702  ( .A(\UART_RXFF/iFIFOMem[34][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2074 ) );
  notech_mux2 \UART_RXFF/U701  ( .A(\UART_RXFF/iFIFOMem[34][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n362 ), .Z(\UART_RXFF/n2075 ) );
  notech_and2 \UART_RXFF/U700  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n361 ) );
  notech_mux2 \UART_RXFF/U699  ( .A(\UART_RXFF/iFIFOMem[35][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2076 ) );
  notech_mux2 \UART_RXFF/U698  ( .A(\UART_RXFF/iFIFOMem[35][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2077 ) );
  notech_mux2 \UART_RXFF/U697  ( .A(\UART_RXFF/iFIFOMem[35][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2078 ) );
  notech_mux2 \UART_RXFF/U696  ( .A(\UART_RXFF/iFIFOMem[35][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2079 ) );
  notech_mux2 \UART_RXFF/U695  ( .A(\UART_RXFF/iFIFOMem[35][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2080 ) );
  notech_mux2 \UART_RXFF/U694  ( .A(\UART_RXFF/iFIFOMem[35][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2081 ) );
  notech_mux2 \UART_RXFF/U693  ( .A(\UART_RXFF/iFIFOMem[35][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2082 ) );
  notech_mux2 \UART_RXFF/U692  ( .A(\UART_RXFF/iFIFOMem[35][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2083 ) );
  notech_mux2 \UART_RXFF/U691  ( .A(\UART_RXFF/iFIFOMem[35][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2084 ) );
  notech_mux2 \UART_RXFF/U690  ( .A(\UART_RXFF/iFIFOMem[35][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2085 ) );
  notech_mux2 \UART_RXFF/U689  ( .A(\UART_RXFF/iFIFOMem[35][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n361 ), .Z(\UART_RXFF/n2086 ) );
  notech_and2 \UART_RXFF/U688  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n360 ) );
  notech_mux2 \UART_RXFF/U687  ( .A(\UART_RXFF/iFIFOMem[36][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2087 ) );
  notech_mux2 \UART_RXFF/U686  ( .A(\UART_RXFF/iFIFOMem[36][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2088 ) );
  notech_mux2 \UART_RXFF/U685  ( .A(\UART_RXFF/iFIFOMem[36][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2089 ) );
  notech_mux2 \UART_RXFF/U684  ( .A(\UART_RXFF/iFIFOMem[36][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2090 ) );
  notech_mux2 \UART_RXFF/U683  ( .A(\UART_RXFF/iFIFOMem[36][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2091 ) );
  notech_mux2 \UART_RXFF/U682  ( .A(\UART_RXFF/iFIFOMem[36][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2092 ) );
  notech_mux2 \UART_RXFF/U681  ( .A(\UART_RXFF/iFIFOMem[36][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2093 ) );
  notech_mux2 \UART_RXFF/U680  ( .A(\UART_RXFF/iFIFOMem[36][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2094 ) );
  notech_mux2 \UART_RXFF/U679  ( .A(\UART_RXFF/iFIFOMem[36][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2095 ) );
  notech_mux2 \UART_RXFF/U678  ( .A(\UART_RXFF/iFIFOMem[36][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2096 ) );
  notech_mux2 \UART_RXFF/U677  ( .A(\UART_RXFF/iFIFOMem[36][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n360 ), .Z(\UART_RXFF/n2097 ) );
  notech_and2 \UART_RXFF/U676  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n359 ) );
  notech_mux2 \UART_RXFF/U675  ( .A(\UART_RXFF/iFIFOMem[37][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2098 ) );
  notech_mux2 \UART_RXFF/U674  ( .A(\UART_RXFF/iFIFOMem[37][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2099 ) );
  notech_mux2 \UART_RXFF/U673  ( .A(\UART_RXFF/iFIFOMem[37][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2100 ) );
  notech_mux2 \UART_RXFF/U672  ( .A(\UART_RXFF/iFIFOMem[37][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2101 ) );
  notech_mux2 \UART_RXFF/U671  ( .A(\UART_RXFF/iFIFOMem[37][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2102 ) );
  notech_mux2 \UART_RXFF/U670  ( .A(\UART_RXFF/iFIFOMem[37][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2103 ) );
  notech_mux2 \UART_RXFF/U669  ( .A(\UART_RXFF/iFIFOMem[37][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2104 ) );
  notech_mux2 \UART_RXFF/U668  ( .A(\UART_RXFF/iFIFOMem[37][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2105 ) );
  notech_mux2 \UART_RXFF/U667  ( .A(\UART_RXFF/iFIFOMem[37][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2106 ) );
  notech_mux2 \UART_RXFF/U666  ( .A(\UART_RXFF/iFIFOMem[37][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2107 ) );
  notech_mux2 \UART_RXFF/U665  ( .A(\UART_RXFF/iFIFOMem[37][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n359 ), .Z(\UART_RXFF/n2108 ) );
  notech_and2 \UART_RXFF/U664  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n358 ) );
  notech_mux2 \UART_RXFF/U663  ( .A(\UART_RXFF/iFIFOMem[38][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2109 ) );
  notech_mux2 \UART_RXFF/U662  ( .A(\UART_RXFF/iFIFOMem[38][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2110 ) );
  notech_mux2 \UART_RXFF/U661  ( .A(\UART_RXFF/iFIFOMem[38][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2111 ) );
  notech_mux2 \UART_RXFF/U660  ( .A(\UART_RXFF/iFIFOMem[38][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2112 ) );
  notech_mux2 \UART_RXFF/U659  ( .A(\UART_RXFF/iFIFOMem[38][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2113 ) );
  notech_mux2 \UART_RXFF/U658  ( .A(\UART_RXFF/iFIFOMem[38][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2114 ) );
  notech_mux2 \UART_RXFF/U657  ( .A(\UART_RXFF/iFIFOMem[38][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2115 ) );
  notech_mux2 \UART_RXFF/U656  ( .A(\UART_RXFF/iFIFOMem[38][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2116 ) );
  notech_mux2 \UART_RXFF/U655  ( .A(\UART_RXFF/iFIFOMem[38][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2117 ) );
  notech_mux2 \UART_RXFF/U654  ( .A(\UART_RXFF/iFIFOMem[38][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2118 ) );
  notech_mux2 \UART_RXFF/U653  ( .A(\UART_RXFF/iFIFOMem[38][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n358 ), .Z(\UART_RXFF/n2119 ) );
  notech_and2 \UART_RXFF/U652  ( .A(\UART_RXFF/n357 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n356 ) );
  notech_mux2 \UART_RXFF/U651  ( .A(\UART_RXFF/iFIFOMem[39][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2120 ) );
  notech_mux2 \UART_RXFF/U650  ( .A(\UART_RXFF/iFIFOMem[39][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2121 ) );
  notech_mux2 \UART_RXFF/U649  ( .A(\UART_RXFF/iFIFOMem[39][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2122 ) );
  notech_mux2 \UART_RXFF/U648  ( .A(\UART_RXFF/iFIFOMem[39][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2123 ) );
  notech_mux2 \UART_RXFF/U647  ( .A(\UART_RXFF/iFIFOMem[39][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2124 ) );
  notech_mux2 \UART_RXFF/U646  ( .A(\UART_RXFF/iFIFOMem[39][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2125 ) );
  notech_mux2 \UART_RXFF/U645  ( .A(\UART_RXFF/iFIFOMem[39][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2126 ) );
  notech_mux2 \UART_RXFF/U644  ( .A(\UART_RXFF/iFIFOMem[39][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2127 ) );
  notech_mux2 \UART_RXFF/U643  ( .A(\UART_RXFF/iFIFOMem[39][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2128 ) );
  notech_mux2 \UART_RXFF/U642  ( .A(\UART_RXFF/iFIFOMem[39][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2129 ) );
  notech_mux2 \UART_RXFF/U641  ( .A(\UART_RXFF/iFIFOMem[39][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n356 ), .Z(\UART_RXFF/n2130 ) );
  notech_ao3 \UART_RXFF/U640  ( .A(\UART_RXFF/iWRAddr[3] ), .B(
        \UART_RXFF/n337 ), .C(\UART_RXFF/iWRAddr[4] ), .Z(\UART_RXFF/n348 ) );
  notech_and2 \UART_RXFF/U639  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n355 ) );
  notech_mux2 \UART_RXFF/U638  ( .A(\UART_RXFF/iFIFOMem[40][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2131 ) );
  notech_mux2 \UART_RXFF/U637  ( .A(\UART_RXFF/iFIFOMem[40][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2132 ) );
  notech_mux2 \UART_RXFF/U636  ( .A(\UART_RXFF/iFIFOMem[40][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2133 ) );
  notech_mux2 \UART_RXFF/U635  ( .A(\UART_RXFF/iFIFOMem[40][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2134 ) );
  notech_mux2 \UART_RXFF/U634  ( .A(\UART_RXFF/iFIFOMem[40][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2135 ) );
  notech_mux2 \UART_RXFF/U633  ( .A(\UART_RXFF/iFIFOMem[40][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2136 ) );
  notech_mux2 \UART_RXFF/U632  ( .A(\UART_RXFF/iFIFOMem[40][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2137 ) );
  notech_mux2 \UART_RXFF/U631  ( .A(\UART_RXFF/iFIFOMem[40][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2138 ) );
  notech_mux2 \UART_RXFF/U630  ( .A(\UART_RXFF/iFIFOMem[40][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2139 ) );
  notech_mux2 \UART_RXFF/U629  ( .A(\UART_RXFF/iFIFOMem[40][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2140 ) );
  notech_mux2 \UART_RXFF/U628  ( .A(\UART_RXFF/iFIFOMem[40][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n355 ), .Z(\UART_RXFF/n2141 ) );
  notech_and2 \UART_RXFF/U627  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n354 ) );
  notech_mux2 \UART_RXFF/U626  ( .A(\UART_RXFF/iFIFOMem[41][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2142 ) );
  notech_mux2 \UART_RXFF/U625  ( .A(\UART_RXFF/iFIFOMem[41][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2143 ) );
  notech_mux2 \UART_RXFF/U624  ( .A(\UART_RXFF/iFIFOMem[41][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2144 ) );
  notech_mux2 \UART_RXFF/U623  ( .A(\UART_RXFF/iFIFOMem[41][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2145 ) );
  notech_mux2 \UART_RXFF/U622  ( .A(\UART_RXFF/iFIFOMem[41][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2146 ) );
  notech_mux2 \UART_RXFF/U621  ( .A(\UART_RXFF/iFIFOMem[41][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2147 ) );
  notech_mux2 \UART_RXFF/U620  ( .A(\UART_RXFF/iFIFOMem[41][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2148 ) );
  notech_mux2 \UART_RXFF/U619  ( .A(\UART_RXFF/iFIFOMem[41][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2149 ) );
  notech_mux2 \UART_RXFF/U618  ( .A(\UART_RXFF/iFIFOMem[41][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2150 ) );
  notech_mux2 \UART_RXFF/U617  ( .A(\UART_RXFF/iFIFOMem[41][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2151 ) );
  notech_mux2 \UART_RXFF/U616  ( .A(\UART_RXFF/iFIFOMem[41][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n354 ), .Z(\UART_RXFF/n2152 ) );
  notech_and2 \UART_RXFF/U615  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n353 ) );
  notech_mux2 \UART_RXFF/U614  ( .A(\UART_RXFF/iFIFOMem[42][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2153 ) );
  notech_mux2 \UART_RXFF/U613  ( .A(\UART_RXFF/iFIFOMem[42][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2154 ) );
  notech_mux2 \UART_RXFF/U612  ( .A(\UART_RXFF/iFIFOMem[42][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2155 ) );
  notech_mux2 \UART_RXFF/U611  ( .A(\UART_RXFF/iFIFOMem[42][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2156 ) );
  notech_mux2 \UART_RXFF/U610  ( .A(\UART_RXFF/iFIFOMem[42][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2157 ) );
  notech_mux2 \UART_RXFF/U609  ( .A(\UART_RXFF/iFIFOMem[42][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2158 ) );
  notech_mux2 \UART_RXFF/U608  ( .A(\UART_RXFF/iFIFOMem[42][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2159 ) );
  notech_mux2 \UART_RXFF/U607  ( .A(\UART_RXFF/iFIFOMem[42][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2160 ) );
  notech_mux2 \UART_RXFF/U606  ( .A(\UART_RXFF/iFIFOMem[42][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2161 ) );
  notech_mux2 \UART_RXFF/U605  ( .A(\UART_RXFF/iFIFOMem[42][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2162 ) );
  notech_mux2 \UART_RXFF/U604  ( .A(\UART_RXFF/iFIFOMem[42][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n353 ), .Z(\UART_RXFF/n2163 ) );
  notech_and2 \UART_RXFF/U603  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n352 ) );
  notech_mux2 \UART_RXFF/U602  ( .A(\UART_RXFF/iFIFOMem[43][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2164 ) );
  notech_mux2 \UART_RXFF/U601  ( .A(\UART_RXFF/iFIFOMem[43][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2165 ) );
  notech_mux2 \UART_RXFF/U600  ( .A(\UART_RXFF/iFIFOMem[43][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2166 ) );
  notech_mux2 \UART_RXFF/U599  ( .A(\UART_RXFF/iFIFOMem[43][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2167 ) );
  notech_mux2 \UART_RXFF/U598  ( .A(\UART_RXFF/iFIFOMem[43][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2168 ) );
  notech_mux2 \UART_RXFF/U597  ( .A(\UART_RXFF/iFIFOMem[43][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2169 ) );
  notech_mux2 \UART_RXFF/U596  ( .A(\UART_RXFF/iFIFOMem[43][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2170 ) );
  notech_mux2 \UART_RXFF/U595  ( .A(\UART_RXFF/iFIFOMem[43][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2171 ) );
  notech_mux2 \UART_RXFF/U594  ( .A(\UART_RXFF/iFIFOMem[43][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2172 ) );
  notech_mux2 \UART_RXFF/U593  ( .A(\UART_RXFF/iFIFOMem[43][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2173 ) );
  notech_mux2 \UART_RXFF/U592  ( .A(\UART_RXFF/iFIFOMem[43][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n352 ), .Z(\UART_RXFF/n2174 ) );
  notech_and2 \UART_RXFF/U591  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n351 ) );
  notech_mux2 \UART_RXFF/U590  ( .A(\UART_RXFF/iFIFOMem[44][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2175 ) );
  notech_mux2 \UART_RXFF/U589  ( .A(\UART_RXFF/iFIFOMem[44][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2176 ) );
  notech_mux2 \UART_RXFF/U588  ( .A(\UART_RXFF/iFIFOMem[44][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2177 ) );
  notech_mux2 \UART_RXFF/U587  ( .A(\UART_RXFF/iFIFOMem[44][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2178 ) );
  notech_mux2 \UART_RXFF/U586  ( .A(\UART_RXFF/iFIFOMem[44][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2179 ) );
  notech_mux2 \UART_RXFF/U585  ( .A(\UART_RXFF/iFIFOMem[44][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2180 ) );
  notech_mux2 \UART_RXFF/U584  ( .A(\UART_RXFF/iFIFOMem[44][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2181 ) );
  notech_mux2 \UART_RXFF/U583  ( .A(\UART_RXFF/iFIFOMem[44][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2182 ) );
  notech_mux2 \UART_RXFF/U582  ( .A(\UART_RXFF/iFIFOMem[44][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2183 ) );
  notech_mux2 \UART_RXFF/U581  ( .A(\UART_RXFF/iFIFOMem[44][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2184 ) );
  notech_mux2 \UART_RXFF/U580  ( .A(\UART_RXFF/iFIFOMem[44][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n351 ), .Z(\UART_RXFF/n2185 ) );
  notech_and2 \UART_RXFF/U579  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n350 ) );
  notech_mux2 \UART_RXFF/U578  ( .A(\UART_RXFF/iFIFOMem[45][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2186 ) );
  notech_mux2 \UART_RXFF/U577  ( .A(\UART_RXFF/iFIFOMem[45][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2187 ) );
  notech_mux2 \UART_RXFF/U576  ( .A(\UART_RXFF/iFIFOMem[45][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2188 ) );
  notech_mux2 \UART_RXFF/U575  ( .A(\UART_RXFF/iFIFOMem[45][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2189 ) );
  notech_mux2 \UART_RXFF/U574  ( .A(\UART_RXFF/iFIFOMem[45][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2190 ) );
  notech_mux2 \UART_RXFF/U573  ( .A(\UART_RXFF/iFIFOMem[45][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2191 ) );
  notech_mux2 \UART_RXFF/U572  ( .A(\UART_RXFF/iFIFOMem[45][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2192 ) );
  notech_mux2 \UART_RXFF/U571  ( .A(\UART_RXFF/iFIFOMem[45][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2193 ) );
  notech_mux2 \UART_RXFF/U570  ( .A(\UART_RXFF/iFIFOMem[45][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2194 ) );
  notech_mux2 \UART_RXFF/U569  ( .A(\UART_RXFF/iFIFOMem[45][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2195 ) );
  notech_mux2 \UART_RXFF/U568  ( .A(\UART_RXFF/iFIFOMem[45][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n350 ), .Z(\UART_RXFF/n2196 ) );
  notech_and2 \UART_RXFF/U567  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n349 ) );
  notech_mux2 \UART_RXFF/U566  ( .A(\UART_RXFF/iFIFOMem[46][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2197 ) );
  notech_mux2 \UART_RXFF/U565  ( .A(\UART_RXFF/iFIFOMem[46][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2198 ) );
  notech_mux2 \UART_RXFF/U564  ( .A(\UART_RXFF/iFIFOMem[46][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2199 ) );
  notech_mux2 \UART_RXFF/U563  ( .A(\UART_RXFF/iFIFOMem[46][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2200 ) );
  notech_mux2 \UART_RXFF/U562  ( .A(\UART_RXFF/iFIFOMem[46][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2201 ) );
  notech_mux2 \UART_RXFF/U561  ( .A(\UART_RXFF/iFIFOMem[46][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2202 ) );
  notech_mux2 \UART_RXFF/U560  ( .A(\UART_RXFF/iFIFOMem[46][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2203 ) );
  notech_mux2 \UART_RXFF/U559  ( .A(\UART_RXFF/iFIFOMem[46][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2204 ) );
  notech_mux2 \UART_RXFF/U558  ( .A(\UART_RXFF/iFIFOMem[46][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2205 ) );
  notech_mux2 \UART_RXFF/U557  ( .A(\UART_RXFF/iFIFOMem[46][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2206 ) );
  notech_mux2 \UART_RXFF/U556  ( .A(\UART_RXFF/iFIFOMem[46][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n349 ), .Z(\UART_RXFF/n2207 ) );
  notech_and2 \UART_RXFF/U555  ( .A(\UART_RXFF/n348 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n347 ) );
  notech_mux2 \UART_RXFF/U554  ( .A(\UART_RXFF/iFIFOMem[47][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2208 ) );
  notech_mux2 \UART_RXFF/U553  ( .A(\UART_RXFF/iFIFOMem[47][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2209 ) );
  notech_mux2 \UART_RXFF/U552  ( .A(\UART_RXFF/iFIFOMem[47][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2210 ) );
  notech_mux2 \UART_RXFF/U551  ( .A(\UART_RXFF/iFIFOMem[47][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2211 ) );
  notech_mux2 \UART_RXFF/U550  ( .A(\UART_RXFF/iFIFOMem[47][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2212 ) );
  notech_mux2 \UART_RXFF/U549  ( .A(\UART_RXFF/iFIFOMem[47][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2213 ) );
  notech_mux2 \UART_RXFF/U548  ( .A(\UART_RXFF/iFIFOMem[47][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2214 ) );
  notech_mux2 \UART_RXFF/U547  ( .A(\UART_RXFF/iFIFOMem[47][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2215 ) );
  notech_mux2 \UART_RXFF/U546  ( .A(\UART_RXFF/iFIFOMem[47][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2216 ) );
  notech_mux2 \UART_RXFF/U545  ( .A(\UART_RXFF/iFIFOMem[47][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2217 ) );
  notech_mux2 \UART_RXFF/U544  ( .A(\UART_RXFF/iFIFOMem[47][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n347 ), .Z(\UART_RXFF/n2218 ) );
  notech_ao3 \UART_RXFF/U543  ( .A(\UART_RXFF/iWRAddr[4] ), .B(
        \UART_RXFF/n337 ), .C(\UART_RXFF/iWRAddr[3] ), .Z(\UART_RXFF/n339 ) );
  notech_and2 \UART_RXFF/U542  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n346 ) );
  notech_mux2 \UART_RXFF/U541  ( .A(\UART_RXFF/iFIFOMem[48][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2219 ) );
  notech_mux2 \UART_RXFF/U540  ( .A(\UART_RXFF/iFIFOMem[48][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2220 ) );
  notech_mux2 \UART_RXFF/U539  ( .A(\UART_RXFF/iFIFOMem[48][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2221 ) );
  notech_mux2 \UART_RXFF/U538  ( .A(\UART_RXFF/iFIFOMem[48][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2222 ) );
  notech_mux2 \UART_RXFF/U537  ( .A(\UART_RXFF/iFIFOMem[48][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2223 ) );
  notech_mux2 \UART_RXFF/U536  ( .A(\UART_RXFF/iFIFOMem[48][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2224 ) );
  notech_mux2 \UART_RXFF/U535  ( .A(\UART_RXFF/iFIFOMem[48][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2225 ) );
  notech_mux2 \UART_RXFF/U534  ( .A(\UART_RXFF/iFIFOMem[48][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2226 ) );
  notech_mux2 \UART_RXFF/U533  ( .A(\UART_RXFF/iFIFOMem[48][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2227 ) );
  notech_mux2 \UART_RXFF/U532  ( .A(\UART_RXFF/iFIFOMem[48][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2228 ) );
  notech_mux2 \UART_RXFF/U531  ( .A(\UART_RXFF/iFIFOMem[48][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n346 ), .Z(\UART_RXFF/n2229 ) );
  notech_and2 \UART_RXFF/U530  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n345 ) );
  notech_mux2 \UART_RXFF/U529  ( .A(\UART_RXFF/iFIFOMem[49][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2230 ) );
  notech_mux2 \UART_RXFF/U528  ( .A(\UART_RXFF/iFIFOMem[49][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2231 ) );
  notech_mux2 \UART_RXFF/U527  ( .A(\UART_RXFF/iFIFOMem[49][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2232 ) );
  notech_mux2 \UART_RXFF/U526  ( .A(\UART_RXFF/iFIFOMem[49][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2233 ) );
  notech_mux2 \UART_RXFF/U525  ( .A(\UART_RXFF/iFIFOMem[49][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2234 ) );
  notech_mux2 \UART_RXFF/U524  ( .A(\UART_RXFF/iFIFOMem[49][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2235 ) );
  notech_mux2 \UART_RXFF/U523  ( .A(\UART_RXFF/iFIFOMem[49][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2236 ) );
  notech_mux2 \UART_RXFF/U522  ( .A(\UART_RXFF/iFIFOMem[49][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2237 ) );
  notech_mux2 \UART_RXFF/U521  ( .A(\UART_RXFF/iFIFOMem[49][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2238 ) );
  notech_mux2 \UART_RXFF/U520  ( .A(\UART_RXFF/iFIFOMem[49][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2239 ) );
  notech_mux2 \UART_RXFF/U519  ( .A(\UART_RXFF/iFIFOMem[49][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n345 ), .Z(\UART_RXFF/n2240 ) );
  notech_and2 \UART_RXFF/U518  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n344 ) );
  notech_mux2 \UART_RXFF/U517  ( .A(\UART_RXFF/iFIFOMem[50][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2241 ) );
  notech_mux2 \UART_RXFF/U516  ( .A(\UART_RXFF/iFIFOMem[50][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2242 ) );
  notech_mux2 \UART_RXFF/U515  ( .A(\UART_RXFF/iFIFOMem[50][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2243 ) );
  notech_mux2 \UART_RXFF/U514  ( .A(\UART_RXFF/iFIFOMem[50][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2244 ) );
  notech_mux2 \UART_RXFF/U513  ( .A(\UART_RXFF/iFIFOMem[50][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2245 ) );
  notech_mux2 \UART_RXFF/U512  ( .A(\UART_RXFF/iFIFOMem[50][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2246 ) );
  notech_mux2 \UART_RXFF/U511  ( .A(\UART_RXFF/iFIFOMem[50][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2247 ) );
  notech_mux2 \UART_RXFF/U510  ( .A(\UART_RXFF/iFIFOMem[50][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2248 ) );
  notech_mux2 \UART_RXFF/U509  ( .A(\UART_RXFF/iFIFOMem[50][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2249 ) );
  notech_mux2 \UART_RXFF/U508  ( .A(\UART_RXFF/iFIFOMem[50][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2250 ) );
  notech_mux2 \UART_RXFF/U507  ( .A(\UART_RXFF/iFIFOMem[50][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n344 ), .Z(\UART_RXFF/n2251 ) );
  notech_and2 \UART_RXFF/U506  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n343 ) );
  notech_mux2 \UART_RXFF/U505  ( .A(\UART_RXFF/iFIFOMem[51][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2252 ) );
  notech_mux2 \UART_RXFF/U504  ( .A(\UART_RXFF/iFIFOMem[51][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2253 ) );
  notech_mux2 \UART_RXFF/U503  ( .A(\UART_RXFF/iFIFOMem[51][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2254 ) );
  notech_mux2 \UART_RXFF/U502  ( .A(\UART_RXFF/iFIFOMem[51][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2255 ) );
  notech_mux2 \UART_RXFF/U501  ( .A(\UART_RXFF/iFIFOMem[51][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2256 ) );
  notech_mux2 \UART_RXFF/U500  ( .A(\UART_RXFF/iFIFOMem[51][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2257 ) );
  notech_mux2 \UART_RXFF/U499  ( .A(\UART_RXFF/iFIFOMem[51][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2258 ) );
  notech_mux2 \UART_RXFF/U498  ( .A(\UART_RXFF/iFIFOMem[51][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2259 ) );
  notech_mux2 \UART_RXFF/U497  ( .A(\UART_RXFF/iFIFOMem[51][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2260 ) );
  notech_mux2 \UART_RXFF/U496  ( .A(\UART_RXFF/iFIFOMem[51][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2261 ) );
  notech_mux2 \UART_RXFF/U495  ( .A(\UART_RXFF/iFIFOMem[51][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n343 ), .Z(\UART_RXFF/n2262 ) );
  notech_and2 \UART_RXFF/U494  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n342 ) );
  notech_mux2 \UART_RXFF/U493  ( .A(\UART_RXFF/iFIFOMem[52][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2263 ) );
  notech_mux2 \UART_RXFF/U492  ( .A(\UART_RXFF/iFIFOMem[52][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2264 ) );
  notech_mux2 \UART_RXFF/U491  ( .A(\UART_RXFF/iFIFOMem[52][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2265 ) );
  notech_mux2 \UART_RXFF/U490  ( .A(\UART_RXFF/iFIFOMem[52][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2266 ) );
  notech_mux2 \UART_RXFF/U489  ( .A(\UART_RXFF/iFIFOMem[52][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2267 ) );
  notech_mux2 \UART_RXFF/U488  ( .A(\UART_RXFF/iFIFOMem[52][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2268 ) );
  notech_mux2 \UART_RXFF/U487  ( .A(\UART_RXFF/iFIFOMem[52][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2269 ) );
  notech_mux2 \UART_RXFF/U486  ( .A(\UART_RXFF/iFIFOMem[52][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2270 ) );
  notech_mux2 \UART_RXFF/U485  ( .A(\UART_RXFF/iFIFOMem[52][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2271 ) );
  notech_mux2 \UART_RXFF/U484  ( .A(\UART_RXFF/iFIFOMem[52][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2272 ) );
  notech_mux2 \UART_RXFF/U483  ( .A(\UART_RXFF/iFIFOMem[52][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n342 ), .Z(\UART_RXFF/n2273 ) );
  notech_and2 \UART_RXFF/U482  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n341 ) );
  notech_mux2 \UART_RXFF/U481  ( .A(\UART_RXFF/iFIFOMem[53][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2274 ) );
  notech_mux2 \UART_RXFF/U480  ( .A(\UART_RXFF/iFIFOMem[53][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2275 ) );
  notech_mux2 \UART_RXFF/U479  ( .A(\UART_RXFF/iFIFOMem[53][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2276 ) );
  notech_mux2 \UART_RXFF/U478  ( .A(\UART_RXFF/iFIFOMem[53][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2277 ) );
  notech_mux2 \UART_RXFF/U477  ( .A(\UART_RXFF/iFIFOMem[53][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2278 ) );
  notech_mux2 \UART_RXFF/U476  ( .A(\UART_RXFF/iFIFOMem[53][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2279 ) );
  notech_mux2 \UART_RXFF/U475  ( .A(\UART_RXFF/iFIFOMem[53][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2280 ) );
  notech_mux2 \UART_RXFF/U474  ( .A(\UART_RXFF/iFIFOMem[53][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2281 ) );
  notech_mux2 \UART_RXFF/U473  ( .A(\UART_RXFF/iFIFOMem[53][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2282 ) );
  notech_mux2 \UART_RXFF/U472  ( .A(\UART_RXFF/iFIFOMem[53][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2283 ) );
  notech_mux2 \UART_RXFF/U471  ( .A(\UART_RXFF/iFIFOMem[53][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n341 ), .Z(\UART_RXFF/n2284 ) );
  notech_and2 \UART_RXFF/U470  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n340 ) );
  notech_mux2 \UART_RXFF/U469  ( .A(\UART_RXFF/iFIFOMem[54][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2285 ) );
  notech_mux2 \UART_RXFF/U468  ( .A(\UART_RXFF/iFIFOMem[54][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2286 ) );
  notech_mux2 \UART_RXFF/U467  ( .A(\UART_RXFF/iFIFOMem[54][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2287 ) );
  notech_mux2 \UART_RXFF/U466  ( .A(\UART_RXFF/iFIFOMem[54][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2288 ) );
  notech_mux2 \UART_RXFF/U465  ( .A(\UART_RXFF/iFIFOMem[54][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2289 ) );
  notech_mux2 \UART_RXFF/U464  ( .A(\UART_RXFF/iFIFOMem[54][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2290 ) );
  notech_mux2 \UART_RXFF/U463  ( .A(\UART_RXFF/iFIFOMem[54][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2291 ) );
  notech_mux2 \UART_RXFF/U462  ( .A(\UART_RXFF/iFIFOMem[54][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2292 ) );
  notech_mux2 \UART_RXFF/U461  ( .A(\UART_RXFF/iFIFOMem[54][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2293 ) );
  notech_mux2 \UART_RXFF/U460  ( .A(\UART_RXFF/iFIFOMem[54][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2294 ) );
  notech_mux2 \UART_RXFF/U459  ( .A(\UART_RXFF/iFIFOMem[54][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n340 ), .Z(\UART_RXFF/n2295 ) );
  notech_and2 \UART_RXFF/U458  ( .A(\UART_RXFF/n339 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n338 ) );
  notech_mux2 \UART_RXFF/U457  ( .A(\UART_RXFF/iFIFOMem[55][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2296 ) );
  notech_mux2 \UART_RXFF/U456  ( .A(\UART_RXFF/iFIFOMem[55][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2297 ) );
  notech_mux2 \UART_RXFF/U455  ( .A(\UART_RXFF/iFIFOMem[55][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2298 ) );
  notech_mux2 \UART_RXFF/U454  ( .A(\UART_RXFF/iFIFOMem[55][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2299 ) );
  notech_mux2 \UART_RXFF/U453  ( .A(\UART_RXFF/iFIFOMem[55][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2300 ) );
  notech_mux2 \UART_RXFF/U452  ( .A(\UART_RXFF/iFIFOMem[55][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2301 ) );
  notech_mux2 \UART_RXFF/U451  ( .A(\UART_RXFF/iFIFOMem[55][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2302 ) );
  notech_mux2 \UART_RXFF/U450  ( .A(\UART_RXFF/iFIFOMem[55][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2303 ) );
  notech_mux2 \UART_RXFF/U449  ( .A(\UART_RXFF/iFIFOMem[55][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2304 ) );
  notech_mux2 \UART_RXFF/U448  ( .A(\UART_RXFF/iFIFOMem[55][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2305 ) );
  notech_mux2 \UART_RXFF/U447  ( .A(\UART_RXFF/iFIFOMem[55][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n338 ), .Z(\UART_RXFF/n2306 ) );
  notech_and3 \UART_RXFF/U446  ( .A(\UART_RXFF/iWRAddr[4] ), .B(
        \UART_RXFF/n337 ), .C(\UART_RXFF/iWRAddr[3] ), .Z(\UART_RXFF/n321 ) );
  notech_and2 \UART_RXFF/U445  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n336 ), 
        .Z(\UART_RXFF/n335 ) );
  notech_mux2 \UART_RXFF/U444  ( .A(\UART_RXFF/iFIFOMem[56][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2307 ) );
  notech_mux2 \UART_RXFF/U443  ( .A(\UART_RXFF/iFIFOMem[56][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2308 ) );
  notech_mux2 \UART_RXFF/U442  ( .A(\UART_RXFF/iFIFOMem[56][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2309 ) );
  notech_mux2 \UART_RXFF/U441  ( .A(\UART_RXFF/iFIFOMem[56][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2310 ) );
  notech_mux2 \UART_RXFF/U440  ( .A(\UART_RXFF/iFIFOMem[56][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2311 ) );
  notech_mux2 \UART_RXFF/U439  ( .A(\UART_RXFF/iFIFOMem[56][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2312 ) );
  notech_mux2 \UART_RXFF/U438  ( .A(\UART_RXFF/iFIFOMem[56][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2313 ) );
  notech_mux2 \UART_RXFF/U437  ( .A(\UART_RXFF/iFIFOMem[56][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2314 ) );
  notech_mux2 \UART_RXFF/U436  ( .A(\UART_RXFF/iFIFOMem[56][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2315 ) );
  notech_mux2 \UART_RXFF/U435  ( .A(\UART_RXFF/iFIFOMem[56][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2316 ) );
  notech_mux2 \UART_RXFF/U434  ( .A(\UART_RXFF/iFIFOMem[56][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n335 ), .Z(\UART_RXFF/n2317 ) );
  notech_and2 \UART_RXFF/U433  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n334 ), 
        .Z(\UART_RXFF/n333 ) );
  notech_mux2 \UART_RXFF/U432  ( .A(\UART_RXFF/iFIFOMem[57][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2318 ) );
  notech_mux2 \UART_RXFF/U431  ( .A(\UART_RXFF/iFIFOMem[57][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2319 ) );
  notech_mux2 \UART_RXFF/U430  ( .A(\UART_RXFF/iFIFOMem[57][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2320 ) );
  notech_mux2 \UART_RXFF/U429  ( .A(\UART_RXFF/iFIFOMem[57][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2321 ) );
  notech_mux2 \UART_RXFF/U428  ( .A(\UART_RXFF/iFIFOMem[57][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2322 ) );
  notech_mux2 \UART_RXFF/U427  ( .A(\UART_RXFF/iFIFOMem[57][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2323 ) );
  notech_mux2 \UART_RXFF/U426  ( .A(\UART_RXFF/iFIFOMem[57][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2324 ) );
  notech_mux2 \UART_RXFF/U425  ( .A(\UART_RXFF/iFIFOMem[57][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2325 ) );
  notech_mux2 \UART_RXFF/U424  ( .A(\UART_RXFF/iFIFOMem[57][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2326 ) );
  notech_mux2 \UART_RXFF/U423  ( .A(\UART_RXFF/iFIFOMem[57][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2327 ) );
  notech_mux2 \UART_RXFF/U422  ( .A(\UART_RXFF/iFIFOMem[57][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n333 ), .Z(\UART_RXFF/n2328 ) );
  notech_and2 \UART_RXFF/U421  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n332 ), 
        .Z(\UART_RXFF/n331 ) );
  notech_mux2 \UART_RXFF/U420  ( .A(\UART_RXFF/iFIFOMem[58][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2329 ) );
  notech_mux2 \UART_RXFF/U419  ( .A(\UART_RXFF/iFIFOMem[58][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2330 ) );
  notech_mux2 \UART_RXFF/U418  ( .A(\UART_RXFF/iFIFOMem[58][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2331 ) );
  notech_mux2 \UART_RXFF/U417  ( .A(\UART_RXFF/iFIFOMem[58][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2332 ) );
  notech_mux2 \UART_RXFF/U416  ( .A(\UART_RXFF/iFIFOMem[58][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2333 ) );
  notech_mux2 \UART_RXFF/U415  ( .A(\UART_RXFF/iFIFOMem[58][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2334 ) );
  notech_mux2 \UART_RXFF/U414  ( .A(\UART_RXFF/iFIFOMem[58][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2335 ) );
  notech_mux2 \UART_RXFF/U413  ( .A(\UART_RXFF/iFIFOMem[58][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2336 ) );
  notech_mux2 \UART_RXFF/U412  ( .A(\UART_RXFF/iFIFOMem[58][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2337 ) );
  notech_mux2 \UART_RXFF/U411  ( .A(\UART_RXFF/iFIFOMem[58][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2338 ) );
  notech_mux2 \UART_RXFF/U410  ( .A(\UART_RXFF/iFIFOMem[58][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n331 ), .Z(\UART_RXFF/n2339 ) );
  notech_and2 \UART_RXFF/U409  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n330 ), 
        .Z(\UART_RXFF/n329 ) );
  notech_mux2 \UART_RXFF/U408  ( .A(\UART_RXFF/iFIFOMem[59][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2340 ) );
  notech_mux2 \UART_RXFF/U407  ( .A(\UART_RXFF/iFIFOMem[59][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2341 ) );
  notech_mux2 \UART_RXFF/U406  ( .A(\UART_RXFF/iFIFOMem[59][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2342 ) );
  notech_mux2 \UART_RXFF/U405  ( .A(\UART_RXFF/iFIFOMem[59][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2343 ) );
  notech_mux2 \UART_RXFF/U404  ( .A(\UART_RXFF/iFIFOMem[59][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2344 ) );
  notech_mux2 \UART_RXFF/U403  ( .A(\UART_RXFF/iFIFOMem[59][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2345 ) );
  notech_mux2 \UART_RXFF/U402  ( .A(\UART_RXFF/iFIFOMem[59][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2346 ) );
  notech_mux2 \UART_RXFF/U401  ( .A(\UART_RXFF/iFIFOMem[59][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2347 ) );
  notech_mux2 \UART_RXFF/U400  ( .A(\UART_RXFF/iFIFOMem[59][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2348 ) );
  notech_mux2 \UART_RXFF/U399  ( .A(\UART_RXFF/iFIFOMem[59][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2349 ) );
  notech_mux2 \UART_RXFF/U398  ( .A(\UART_RXFF/iFIFOMem[59][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n329 ), .Z(\UART_RXFF/n2350 ) );
  notech_and2 \UART_RXFF/U397  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n328 ), 
        .Z(\UART_RXFF/n327 ) );
  notech_mux2 \UART_RXFF/U396  ( .A(\UART_RXFF/iFIFOMem[60][0] ), .B(
        iRXFIFOD[0]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2351 ) );
  notech_mux2 \UART_RXFF/U395  ( .A(\UART_RXFF/iFIFOMem[60][1] ), .B(
        iRXFIFOD[1]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2352 ) );
  notech_mux2 \UART_RXFF/U394  ( .A(\UART_RXFF/iFIFOMem[60][2] ), .B(
        iRXFIFOD[2]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2353 ) );
  notech_mux2 \UART_RXFF/U393  ( .A(\UART_RXFF/iFIFOMem[60][3] ), .B(
        iRXFIFOD[3]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2354 ) );
  notech_mux2 \UART_RXFF/U392  ( .A(\UART_RXFF/iFIFOMem[60][4] ), .B(
        iRXFIFOD[4]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2355 ) );
  notech_mux2 \UART_RXFF/U391  ( .A(\UART_RXFF/iFIFOMem[60][5] ), .B(
        iRXFIFOD[5]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2356 ) );
  notech_mux2 \UART_RXFF/U390  ( .A(\UART_RXFF/iFIFOMem[60][6] ), .B(
        iRXFIFOD[6]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2357 ) );
  notech_mux2 \UART_RXFF/U389  ( .A(\UART_RXFF/iFIFOMem[60][7] ), .B(
        iRXFIFOD[7]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2358 ) );
  notech_mux2 \UART_RXFF/U388  ( .A(\UART_RXFF/iFIFOMem[60][8] ), .B(
        iRXFIFOD[8]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2359 ) );
  notech_mux2 \UART_RXFF/U387  ( .A(\UART_RXFF/iFIFOMem[60][9] ), .B(
        iRXFIFOD[9]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2360 ) );
  notech_mux2 \UART_RXFF/U386  ( .A(\UART_RXFF/iFIFOMem[60][10] ), .B(
        iRXFIFOD[10]), .S(\UART_RXFF/n327 ), .Z(\UART_RXFF/n2361 ) );
  notech_and2 \UART_RXFF/U385  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n326 ), 
        .Z(\UART_RXFF/n325 ) );
  notech_mux2 \UART_RXFF/U384  ( .A(\UART_RXFF/iFIFOMem[61][0] ), .B(
        \UART_RXFF/n4 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2362 ) );
  notech_mux2 \UART_RXFF/U383  ( .A(\UART_RXFF/iFIFOMem[61][1] ), .B(
        \UART_RXFF/n8 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2363 ) );
  notech_mux2 \UART_RXFF/U382  ( .A(\UART_RXFF/iFIFOMem[61][2] ), .B(
        \UART_RXFF/n12 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2364 ) );
  notech_mux2 \UART_RXFF/U381  ( .A(\UART_RXFF/iFIFOMem[61][3] ), .B(
        \UART_RXFF/n16 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2365 ) );
  notech_mux2 \UART_RXFF/U380  ( .A(\UART_RXFF/iFIFOMem[61][4] ), .B(
        \UART_RXFF/n20 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2366 ) );
  notech_mux2 \UART_RXFF/U379  ( .A(\UART_RXFF/iFIFOMem[61][5] ), .B(
        \UART_RXFF/n24 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2367 ) );
  notech_mux2 \UART_RXFF/U378  ( .A(\UART_RXFF/iFIFOMem[61][6] ), .B(
        \UART_RXFF/n28 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2368 ) );
  notech_mux2 \UART_RXFF/U377  ( .A(\UART_RXFF/iFIFOMem[61][7] ), .B(
        \UART_RXFF/n32 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2369 ) );
  notech_mux2 \UART_RXFF/U376  ( .A(\UART_RXFF/iFIFOMem[61][8] ), .B(
        \UART_RXFF/n36 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2370 ) );
  notech_mux2 \UART_RXFF/U375  ( .A(\UART_RXFF/iFIFOMem[61][9] ), .B(
        \UART_RXFF/n40 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2371 ) );
  notech_mux2 \UART_RXFF/U374  ( .A(\UART_RXFF/iFIFOMem[61][10] ), .B(
        \UART_RXFF/n44 ), .S(\UART_RXFF/n325 ), .Z(\UART_RXFF/n2372 ) );
  notech_and2 \UART_RXFF/U373  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n324 ), 
        .Z(\UART_RXFF/n323 ) );
  notech_mux2 \UART_RXFF/U372  ( .A(\UART_RXFF/iFIFOMem[62][0] ), .B(
        \UART_RXFF/n3 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2373 ) );
  notech_mux2 \UART_RXFF/U371  ( .A(\UART_RXFF/iFIFOMem[62][1] ), .B(
        \UART_RXFF/n7 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2374 ) );
  notech_mux2 \UART_RXFF/U370  ( .A(\UART_RXFF/iFIFOMem[62][2] ), .B(
        \UART_RXFF/n11 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2375 ) );
  notech_mux2 \UART_RXFF/U369  ( .A(\UART_RXFF/iFIFOMem[62][3] ), .B(
        \UART_RXFF/n15 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2376 ) );
  notech_mux2 \UART_RXFF/U368  ( .A(\UART_RXFF/iFIFOMem[62][4] ), .B(
        \UART_RXFF/n19 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2377 ) );
  notech_mux2 \UART_RXFF/U367  ( .A(\UART_RXFF/iFIFOMem[62][5] ), .B(
        \UART_RXFF/n23 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2378 ) );
  notech_mux2 \UART_RXFF/U366  ( .A(\UART_RXFF/iFIFOMem[62][6] ), .B(
        \UART_RXFF/n27 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2379 ) );
  notech_mux2 \UART_RXFF/U365  ( .A(\UART_RXFF/iFIFOMem[62][7] ), .B(
        \UART_RXFF/n31 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2380 ) );
  notech_mux2 \UART_RXFF/U364  ( .A(\UART_RXFF/iFIFOMem[62][8] ), .B(
        \UART_RXFF/n35 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2381 ) );
  notech_mux2 \UART_RXFF/U363  ( .A(\UART_RXFF/iFIFOMem[62][9] ), .B(
        \UART_RXFF/n39 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2382 ) );
  notech_mux2 \UART_RXFF/U362  ( .A(\UART_RXFF/iFIFOMem[62][10] ), .B(
        \UART_RXFF/n43 ), .S(\UART_RXFF/n323 ), .Z(\UART_RXFF/n2383 ) );
  notech_and2 \UART_RXFF/U361  ( .A(\UART_RXFF/n321 ), .B(\UART_RXFF/n322 ), 
        .Z(\UART_RXFF/n320 ) );
  notech_mux2 \UART_RXFF/U360  ( .A(\UART_RXFF/iFIFOMem[63][0] ), .B(
        \UART_RXFF/n2 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2384 ) );
  notech_mux2 \UART_RXFF/U359  ( .A(\UART_RXFF/iFIFOMem[63][1] ), .B(
        \UART_RXFF/n6 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2385 ) );
  notech_mux2 \UART_RXFF/U358  ( .A(\UART_RXFF/iFIFOMem[63][2] ), .B(
        \UART_RXFF/n10 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2386 ) );
  notech_mux2 \UART_RXFF/U357  ( .A(\UART_RXFF/iFIFOMem[63][3] ), .B(
        \UART_RXFF/n14 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2387 ) );
  notech_mux2 \UART_RXFF/U356  ( .A(\UART_RXFF/iFIFOMem[63][4] ), .B(
        \UART_RXFF/n18 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2388 ) );
  notech_mux2 \UART_RXFF/U355  ( .A(\UART_RXFF/iFIFOMem[63][5] ), .B(
        \UART_RXFF/n22 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2389 ) );
  notech_mux2 \UART_RXFF/U354  ( .A(\UART_RXFF/iFIFOMem[63][6] ), .B(
        \UART_RXFF/n26 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2390 ) );
  notech_mux2 \UART_RXFF/U353  ( .A(\UART_RXFF/iFIFOMem[63][7] ), .B(
        \UART_RXFF/n30 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2391 ) );
  notech_mux2 \UART_RXFF/U352  ( .A(\UART_RXFF/iFIFOMem[63][8] ), .B(
        \UART_RXFF/n34 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2392 ) );
  notech_mux2 \UART_RXFF/U351  ( .A(\UART_RXFF/iFIFOMem[63][9] ), .B(
        \UART_RXFF/n38 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2393 ) );
  notech_mux2 \UART_RXFF/U350  ( .A(\UART_RXFF/iFIFOMem[63][10] ), .B(
        \UART_RXFF/n42 ), .S(\UART_RXFF/n320 ), .Z(\UART_RXFF/n2394 ) );
  notech_and2 \UART_RXFF/U349  ( .A(n371), .B(n438), .Z(\UART_RXFF/n318 ) );
  notech_or2 \UART_RXFF/U348  ( .A(\UART_RXFF/n318 ), .B(iRXFIFOClear), .Z(
        \UART_RXFF/n292 ) );
  notech_inv \UART_RXFF/U347  ( .A(\UART_RXFF/N17 ), .Z(\UART_RXFF/n316 ) );
  notech_nand2 \UART_RXFF/U346  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n308 ), 
        .Z(\UART_RXFF/n291 ) );
  notech_inv \UART_RXFF/U345  ( .A(\UART_RXFF/N37 ), .Z(\UART_RXFF/n317 ) );
  notech_nao4 \UART_RXFF/U344  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n316 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n317 ), .Z(\UART_RXFF/n2395 ) );
  notech_inv \UART_RXFF/U343  ( .A(\UART_RXFF/N36 ), .Z(\UART_RXFF/n315 ) );
  notech_nao4 \UART_RXFF/U342  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n314 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n315 ), .Z(\UART_RXFF/n2396 ) );
  notech_inv \UART_RXFF/U341  ( .A(\UART_RXFF/N35 ), .Z(\UART_RXFF/n313 ) );
  notech_nao4 \UART_RXFF/U340  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n49 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n313 ), .Z(\UART_RXFF/n2397 ) );
  notech_inv \UART_RXFF/U339  ( .A(\UART_RXFF/N34 ), .Z(\UART_RXFF/n312 ) );
  notech_nao4 \UART_RXFF/U338  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n46 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n312 ), .Z(\UART_RXFF/n2398 ) );
  notech_inv \UART_RXFF/U337  ( .A(\UART_RXFF/N33 ), .Z(\UART_RXFF/n311 ) );
  notech_nao4 \UART_RXFF/U336  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n60 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n311 ), .Z(\UART_RXFF/n2399 ) );
  notech_inv \UART_RXFF/U335  ( .A(\UART_RXFF/iRDAddr[6] ), .Z(
        \UART_RXFF/n309 ) );
  notech_inv \UART_RXFF/U334  ( .A(\UART_RXFF/N38 ), .Z(\UART_RXFF/n310 ) );
  notech_nao4 \UART_RXFF/U333  ( .A(\UART_RXFF/n292 ), .B(\UART_RXFF/n309 ), 
        .C(\UART_RXFF/n291 ), .D(\UART_RXFF/n310 ), .Z(\UART_RXFF/n2400 ) );
  notech_inv \UART_RXFF/U332  ( .A(\UART_RXFF/iWRAddr[5] ), .Z(
        \UART_RXFF/n306 ) );
  notech_nand2 \UART_RXFF/U331  ( .A(\UART_RXFF/n294 ), .B(\UART_RXFF/n308 ), 
        .Z(\UART_RXFF/n295 ) );
  notech_inv \UART_RXFF/U330  ( .A(\UART_RXFF/N29 ), .Z(\UART_RXFF/n307 ) );
  notech_nao4 \UART_RXFF/U329  ( .A(\UART_RXFF/n306 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n307 ), .Z(\UART_RXFF/n2401 ) );
  notech_inv \UART_RXFF/U328  ( .A(\UART_RXFF/iWRAddr[4] ), .Z(
        \UART_RXFF/n304 ) );
  notech_inv \UART_RXFF/U327  ( .A(\UART_RXFF/N28 ), .Z(\UART_RXFF/n305 ) );
  notech_nao4 \UART_RXFF/U326  ( .A(\UART_RXFF/n304 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n305 ), .Z(\UART_RXFF/n2402 ) );
  notech_inv \UART_RXFF/U325  ( .A(\UART_RXFF/N27 ), .Z(\UART_RXFF/n303 ) );
  notech_nao4 \UART_RXFF/U324  ( .A(\UART_RXFF/n302 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n303 ), .Z(\UART_RXFF/n2403 ) );
  notech_inv \UART_RXFF/U323  ( .A(\UART_RXFF/N26 ), .Z(\UART_RXFF/n301 ) );
  notech_nao4 \UART_RXFF/U322  ( .A(\UART_RXFF/n300 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n301 ), .Z(\UART_RXFF/n2404 ) );
  notech_inv \UART_RXFF/U321  ( .A(\UART_RXFF/N25 ), .Z(\UART_RXFF/n299 ) );
  notech_nao4 \UART_RXFF/U320  ( .A(\UART_RXFF/n298 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n299 ), .Z(\UART_RXFF/n2405 ) );
  notech_mux2 \UART_RXFF/U319  ( .A(\UART_RXFF/n295 ), .B(\UART_RXFF/n294 ), 
        .S(\UART_RXFF/iWRAddr[0] ), .Z(\UART_RXFF/n297 ) );
  notech_inv \UART_RXFF/U318  ( .A(\UART_RXFF/n297 ), .Z(\UART_RXFF/n2406 ) );
  notech_inv \UART_RXFF/U317  ( .A(\UART_RXFF/N30 ), .Z(\UART_RXFF/n296 ) );
  notech_nao4 \UART_RXFF/U316  ( .A(\UART_RXFF/n293 ), .B(\UART_RXFF/n294 ), 
        .C(\UART_RXFF/n295 ), .D(\UART_RXFF/n296 ), .Z(\UART_RXFF/n2407 ) );
  notech_mux2 \UART_RXFF/U315  ( .A(\UART_RXFF/n291 ), .B(\UART_RXFF/n292 ), 
        .S(\UART_RXFF/n64 ), .Z(\UART_RXFF/n290 ) );
  notech_inv \UART_RXFF/U314  ( .A(\UART_RXFF/n290 ), .Z(\UART_RXFF/n2408 ) );
  notech_mux2 \UART_RXFF/U313  ( .A(\UART_RXFF/N133 ), .B(iRXFIFOQ[0]), .S(RST), .Z(\UART_RXFF/n959 ) );
  notech_mux2 \UART_RXFF/U312  ( .A(\UART_RXFF/N132 ), .B(iRXFIFOQ[1]), .S(RST), .Z(\UART_RXFF/n961 ) );
  notech_mux2 \UART_RXFF/U311  ( .A(\UART_RXFF/N131 ), .B(iRXFIFOQ[2]), .S(RST), .Z(\UART_RXFF/n963 ) );
  notech_mux2 \UART_RXFF/U310  ( .A(\UART_RXFF/N130 ), .B(iRXFIFOQ[3]), .S(RST), .Z(\UART_RXFF/n965 ) );
  notech_mux2 \UART_RXFF/U309  ( .A(\UART_RXFF/N129 ), .B(iRXFIFOQ[4]), .S(RST), .Z(\UART_RXFF/n967 ) );
  notech_mux2 \UART_RXFF/U308  ( .A(\UART_RXFF/N128 ), .B(iRXFIFOQ[5]), .S(RST), .Z(\UART_RXFF/n969 ) );
  notech_mux2 \UART_RXFF/U307  ( .A(\UART_RXFF/N127 ), .B(iRXFIFOQ[6]), .S(RST), .Z(\UART_RXFF/n971 ) );
  notech_mux2 \UART_RXFF/U306  ( .A(\UART_RXFF/N126 ), .B(iRXFIFOQ[7]), .S(RST), .Z(\UART_RXFF/n973 ) );
  notech_mux2 \UART_RXFF/U305  ( .A(\UART_RXFF/N125 ), .B(iRXFIFOQ[8]), .S(RST), .Z(\UART_RXFF/n975 ) );
  notech_mux2 \UART_RXFF/U304  ( .A(\UART_RXFF/N124 ), .B(iRXFIFOQ[9]), .S(RST), .Z(\UART_RXFF/n977 ) );
  notech_mux2 \UART_RXFF/U303  ( .A(\UART_RXFF/N123 ), .B(iRXFIFOQ[10]), .S(
        RST), .Z(\UART_RXFF/n979 ) );
  notech_mux4 \UART_RXFF/U302  ( .A(\UART_RXFF/n289 ), .B(\UART_RXFF/n279 ), 
        .C(\UART_RXFF/n284 ), .D(\UART_RXFF/n274 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N123 ) );
  notech_mux4 \UART_RXFF/U301  ( .A(\UART_RXFF/n288 ), .B(\UART_RXFF/n286 ), 
        .C(\UART_RXFF/n287 ), .D(\UART_RXFF/n285 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n289 ) );
  notech_mux4 \UART_RXFF/U300  ( .A(\UART_RXFF/iFIFOMem[0][10] ), .B(
        \UART_RXFF/iFIFOMem[2][10] ), .C(\UART_RXFF/iFIFOMem[1][10] ), .D(
        \UART_RXFF/iFIFOMem[3][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n288 ) );
  notech_mux4 \UART_RXFF/U299  ( .A(\UART_RXFF/iFIFOMem[4][10] ), .B(
        \UART_RXFF/iFIFOMem[6][10] ), .C(\UART_RXFF/iFIFOMem[5][10] ), .D(
        \UART_RXFF/iFIFOMem[7][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n287 ) );
  notech_mux4 \UART_RXFF/U298  ( .A(\UART_RXFF/iFIFOMem[8][10] ), .B(
        \UART_RXFF/iFIFOMem[10][10] ), .C(\UART_RXFF/iFIFOMem[9][10] ), .D(
        \UART_RXFF/iFIFOMem[11][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n286 ) );
  notech_mux4 \UART_RXFF/U297  ( .A(\UART_RXFF/iFIFOMem[12][10] ), .B(
        \UART_RXFF/iFIFOMem[14][10] ), .C(\UART_RXFF/iFIFOMem[13][10] ), .D(
        \UART_RXFF/iFIFOMem[15][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n285 ) );
  notech_mux4 \UART_RXFF/U296  ( .A(\UART_RXFF/n283 ), .B(\UART_RXFF/n281 ), 
        .C(\UART_RXFF/n282 ), .D(\UART_RXFF/n280 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n284 ) );
  notech_mux4 \UART_RXFF/U295  ( .A(\UART_RXFF/iFIFOMem[16][10] ), .B(
        \UART_RXFF/iFIFOMem[18][10] ), .C(\UART_RXFF/iFIFOMem[17][10] ), .D(
        \UART_RXFF/iFIFOMem[19][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n283 ) );
  notech_mux4 \UART_RXFF/U294  ( .A(\UART_RXFF/iFIFOMem[20][10] ), .B(
        \UART_RXFF/iFIFOMem[22][10] ), .C(\UART_RXFF/iFIFOMem[21][10] ), .D(
        \UART_RXFF/iFIFOMem[23][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n282 ) );
  notech_mux4 \UART_RXFF/U293  ( .A(\UART_RXFF/iFIFOMem[24][10] ), .B(
        \UART_RXFF/iFIFOMem[26][10] ), .C(\UART_RXFF/iFIFOMem[25][10] ), .D(
        \UART_RXFF/iFIFOMem[27][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n281 ) );
  notech_mux4 \UART_RXFF/U292  ( .A(\UART_RXFF/iFIFOMem[28][10] ), .B(
        \UART_RXFF/iFIFOMem[30][10] ), .C(\UART_RXFF/iFIFOMem[29][10] ), .D(
        \UART_RXFF/iFIFOMem[31][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n280 ) );
  notech_mux4 \UART_RXFF/U291  ( .A(\UART_RXFF/n278 ), .B(\UART_RXFF/n276 ), 
        .C(\UART_RXFF/n277 ), .D(\UART_RXFF/n275 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n279 ) );
  notech_mux4 \UART_RXFF/U290  ( .A(\UART_RXFF/iFIFOMem[32][10] ), .B(
        \UART_RXFF/iFIFOMem[34][10] ), .C(\UART_RXFF/iFIFOMem[33][10] ), .D(
        \UART_RXFF/iFIFOMem[35][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n278 ) );
  notech_mux4 \UART_RXFF/U289  ( .A(\UART_RXFF/iFIFOMem[36][10] ), .B(
        \UART_RXFF/iFIFOMem[38][10] ), .C(\UART_RXFF/iFIFOMem[37][10] ), .D(
        \UART_RXFF/iFIFOMem[39][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n277 ) );
  notech_mux4 \UART_RXFF/U288  ( .A(\UART_RXFF/iFIFOMem[40][10] ), .B(
        \UART_RXFF/iFIFOMem[42][10] ), .C(\UART_RXFF/iFIFOMem[41][10] ), .D(
        \UART_RXFF/iFIFOMem[43][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n276 ) );
  notech_mux4 \UART_RXFF/U287  ( .A(\UART_RXFF/iFIFOMem[44][10] ), .B(
        \UART_RXFF/iFIFOMem[46][10] ), .C(\UART_RXFF/iFIFOMem[45][10] ), .D(
        \UART_RXFF/iFIFOMem[47][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n275 ) );
  notech_mux4 \UART_RXFF/U286  ( .A(\UART_RXFF/n273 ), .B(\UART_RXFF/n271 ), 
        .C(\UART_RXFF/n272 ), .D(\UART_RXFF/n270 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n274 ) );
  notech_mux4 \UART_RXFF/U285  ( .A(\UART_RXFF/iFIFOMem[48][10] ), .B(
        \UART_RXFF/iFIFOMem[50][10] ), .C(\UART_RXFF/iFIFOMem[49][10] ), .D(
        \UART_RXFF/iFIFOMem[51][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n273 ) );
  notech_mux4 \UART_RXFF/U284  ( .A(\UART_RXFF/iFIFOMem[52][10] ), .B(
        \UART_RXFF/iFIFOMem[54][10] ), .C(\UART_RXFF/iFIFOMem[53][10] ), .D(
        \UART_RXFF/iFIFOMem[55][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n272 ) );
  notech_mux4 \UART_RXFF/U283  ( .A(\UART_RXFF/iFIFOMem[56][10] ), .B(
        \UART_RXFF/iFIFOMem[58][10] ), .C(\UART_RXFF/iFIFOMem[57][10] ), .D(
        \UART_RXFF/iFIFOMem[59][10] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n271 ) );
  notech_mux4 \UART_RXFF/U282  ( .A(\UART_RXFF/iFIFOMem[60][10] ), .B(
        \UART_RXFF/iFIFOMem[62][10] ), .C(\UART_RXFF/iFIFOMem[61][10] ), .D(
        \UART_RXFF/iFIFOMem[63][10] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n270 ) );
  notech_mux4 \UART_RXFF/U281  ( .A(\UART_RXFF/n269 ), .B(\UART_RXFF/n259 ), 
        .C(\UART_RXFF/n264 ), .D(\UART_RXFF/n254 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N124 ) );
  notech_mux4 \UART_RXFF/U280  ( .A(\UART_RXFF/n268 ), .B(\UART_RXFF/n266 ), 
        .C(\UART_RXFF/n267 ), .D(\UART_RXFF/n265 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n269 ) );
  notech_mux4 \UART_RXFF/U279  ( .A(\UART_RXFF/iFIFOMem[0][9] ), .B(
        \UART_RXFF/iFIFOMem[2][9] ), .C(\UART_RXFF/iFIFOMem[1][9] ), .D(
        \UART_RXFF/iFIFOMem[3][9] ), .S0(\UART_RXFF/n59 ), .S1(\UART_RXFF/n68 ), .Z(\UART_RXFF/n268 ) );
  notech_mux4 \UART_RXFF/U278  ( .A(\UART_RXFF/iFIFOMem[4][9] ), .B(
        \UART_RXFF/iFIFOMem[6][9] ), .C(\UART_RXFF/iFIFOMem[5][9] ), .D(
        \UART_RXFF/iFIFOMem[7][9] ), .S0(\UART_RXFF/n59 ), .S1(\UART_RXFF/n68 ), .Z(\UART_RXFF/n267 ) );
  notech_mux4 \UART_RXFF/U277  ( .A(\UART_RXFF/iFIFOMem[8][9] ), .B(
        \UART_RXFF/iFIFOMem[10][9] ), .C(\UART_RXFF/iFIFOMem[9][9] ), .D(
        \UART_RXFF/iFIFOMem[11][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n266 ) );
  notech_mux4 \UART_RXFF/U276  ( .A(\UART_RXFF/iFIFOMem[12][9] ), .B(
        \UART_RXFF/iFIFOMem[14][9] ), .C(\UART_RXFF/iFIFOMem[13][9] ), .D(
        \UART_RXFF/iFIFOMem[15][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n265 ) );
  notech_mux4 \UART_RXFF/U275  ( .A(\UART_RXFF/n263 ), .B(\UART_RXFF/n261 ), 
        .C(\UART_RXFF/n262 ), .D(\UART_RXFF/n260 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n264 ) );
  notech_mux4 \UART_RXFF/U274  ( .A(\UART_RXFF/iFIFOMem[16][9] ), .B(
        \UART_RXFF/iFIFOMem[18][9] ), .C(\UART_RXFF/iFIFOMem[17][9] ), .D(
        \UART_RXFF/iFIFOMem[19][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n263 ) );
  notech_mux4 \UART_RXFF/U273  ( .A(\UART_RXFF/iFIFOMem[20][9] ), .B(
        \UART_RXFF/iFIFOMem[22][9] ), .C(\UART_RXFF/iFIFOMem[21][9] ), .D(
        \UART_RXFF/iFIFOMem[23][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n262 ) );
  notech_mux4 \UART_RXFF/U272  ( .A(\UART_RXFF/iFIFOMem[24][9] ), .B(
        \UART_RXFF/iFIFOMem[26][9] ), .C(\UART_RXFF/iFIFOMem[25][9] ), .D(
        \UART_RXFF/iFIFOMem[27][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n261 ) );
  notech_mux4 \UART_RXFF/U271  ( .A(\UART_RXFF/iFIFOMem[28][9] ), .B(
        \UART_RXFF/iFIFOMem[30][9] ), .C(\UART_RXFF/iFIFOMem[29][9] ), .D(
        \UART_RXFF/iFIFOMem[31][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n260 ) );
  notech_mux4 \UART_RXFF/U270  ( .A(\UART_RXFF/n258 ), .B(\UART_RXFF/n256 ), 
        .C(\UART_RXFF/n257 ), .D(\UART_RXFF/n255 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n259 ) );
  notech_mux4 \UART_RXFF/U269  ( .A(\UART_RXFF/iFIFOMem[32][9] ), .B(
        \UART_RXFF/iFIFOMem[34][9] ), .C(\UART_RXFF/iFIFOMem[33][9] ), .D(
        \UART_RXFF/iFIFOMem[35][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n258 ) );
  notech_mux4 \UART_RXFF/U268  ( .A(\UART_RXFF/iFIFOMem[36][9] ), .B(
        \UART_RXFF/iFIFOMem[38][9] ), .C(\UART_RXFF/iFIFOMem[37][9] ), .D(
        \UART_RXFF/iFIFOMem[39][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n257 ) );
  notech_mux4 \UART_RXFF/U267  ( .A(\UART_RXFF/iFIFOMem[40][9] ), .B(
        \UART_RXFF/iFIFOMem[42][9] ), .C(\UART_RXFF/iFIFOMem[41][9] ), .D(
        \UART_RXFF/iFIFOMem[43][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n256 ) );
  notech_mux4 \UART_RXFF/U266  ( .A(\UART_RXFF/iFIFOMem[44][9] ), .B(
        \UART_RXFF/iFIFOMem[46][9] ), .C(\UART_RXFF/iFIFOMem[45][9] ), .D(
        \UART_RXFF/iFIFOMem[47][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n255 ) );
  notech_mux4 \UART_RXFF/U265  ( .A(\UART_RXFF/n253 ), .B(\UART_RXFF/n251 ), 
        .C(\UART_RXFF/n252 ), .D(\UART_RXFF/n250 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n254 ) );
  notech_mux4 \UART_RXFF/U264  ( .A(\UART_RXFF/iFIFOMem[48][9] ), .B(
        \UART_RXFF/iFIFOMem[50][9] ), .C(\UART_RXFF/iFIFOMem[49][9] ), .D(
        \UART_RXFF/iFIFOMem[51][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n253 ) );
  notech_mux4 \UART_RXFF/U263  ( .A(\UART_RXFF/iFIFOMem[52][9] ), .B(
        \UART_RXFF/iFIFOMem[54][9] ), .C(\UART_RXFF/iFIFOMem[53][9] ), .D(
        \UART_RXFF/iFIFOMem[55][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n252 ) );
  notech_mux4 \UART_RXFF/U262  ( .A(\UART_RXFF/iFIFOMem[56][9] ), .B(
        \UART_RXFF/iFIFOMem[58][9] ), .C(\UART_RXFF/iFIFOMem[57][9] ), .D(
        \UART_RXFF/iFIFOMem[59][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n251 ) );
  notech_mux4 \UART_RXFF/U261  ( .A(\UART_RXFF/iFIFOMem[60][9] ), .B(
        \UART_RXFF/iFIFOMem[62][9] ), .C(\UART_RXFF/iFIFOMem[61][9] ), .D(
        \UART_RXFF/iFIFOMem[63][9] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n68 ), .Z(\UART_RXFF/n250 ) );
  notech_mux4 \UART_RXFF/U260  ( .A(\UART_RXFF/n249 ), .B(\UART_RXFF/n239 ), 
        .C(\UART_RXFF/n244 ), .D(\UART_RXFF/n234 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N125 ) );
  notech_mux4 \UART_RXFF/U259  ( .A(\UART_RXFF/n248 ), .B(\UART_RXFF/n246 ), 
        .C(\UART_RXFF/n247 ), .D(\UART_RXFF/n245 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n249 ) );
  notech_mux4 \UART_RXFF/U258  ( .A(\UART_RXFF/iFIFOMem[0][8] ), .B(
        \UART_RXFF/iFIFOMem[2][8] ), .C(\UART_RXFF/iFIFOMem[1][8] ), .D(
        \UART_RXFF/iFIFOMem[3][8] ), .S0(\UART_RXFF/n59 ), .S1(\UART_RXFF/n68 ), .Z(\UART_RXFF/n248 ) );
  notech_mux4 \UART_RXFF/U257  ( .A(\UART_RXFF/iFIFOMem[4][8] ), .B(
        \UART_RXFF/iFIFOMem[6][8] ), .C(\UART_RXFF/iFIFOMem[5][8] ), .D(
        \UART_RXFF/iFIFOMem[7][8] ), .S0(\UART_RXFF/N13 ), .S1(\UART_RXFF/n68 ), .Z(\UART_RXFF/n247 ) );
  notech_mux4 \UART_RXFF/U256  ( .A(\UART_RXFF/iFIFOMem[8][8] ), .B(
        \UART_RXFF/iFIFOMem[10][8] ), .C(\UART_RXFF/iFIFOMem[9][8] ), .D(
        \UART_RXFF/iFIFOMem[11][8] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n246 ) );
  notech_mux4 \UART_RXFF/U255  ( .A(\UART_RXFF/iFIFOMem[12][8] ), .B(
        \UART_RXFF/iFIFOMem[14][8] ), .C(\UART_RXFF/iFIFOMem[13][8] ), .D(
        \UART_RXFF/iFIFOMem[15][8] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n245 ) );
  notech_mux4 \UART_RXFF/U254  ( .A(\UART_RXFF/n243 ), .B(\UART_RXFF/n241 ), 
        .C(\UART_RXFF/n242 ), .D(\UART_RXFF/n240 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n244 ) );
  notech_mux4 \UART_RXFF/U253  ( .A(\UART_RXFF/iFIFOMem[16][8] ), .B(
        \UART_RXFF/iFIFOMem[18][8] ), .C(\UART_RXFF/iFIFOMem[17][8] ), .D(
        \UART_RXFF/iFIFOMem[19][8] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n243 ) );
  notech_mux4 \UART_RXFF/U252  ( .A(\UART_RXFF/iFIFOMem[20][8] ), .B(
        \UART_RXFF/iFIFOMem[22][8] ), .C(\UART_RXFF/iFIFOMem[21][8] ), .D(
        \UART_RXFF/iFIFOMem[23][8] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n242 ) );
  notech_mux4 \UART_RXFF/U251  ( .A(\UART_RXFF/iFIFOMem[24][8] ), .B(
        \UART_RXFF/iFIFOMem[26][8] ), .C(\UART_RXFF/iFIFOMem[25][8] ), .D(
        \UART_RXFF/iFIFOMem[27][8] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n241 ) );
  notech_mux4 \UART_RXFF/U250  ( .A(\UART_RXFF/iFIFOMem[28][8] ), .B(
        \UART_RXFF/iFIFOMem[30][8] ), .C(\UART_RXFF/iFIFOMem[29][8] ), .D(
        \UART_RXFF/iFIFOMem[31][8] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n240 ) );
  notech_mux4 \UART_RXFF/U249  ( .A(\UART_RXFF/n238 ), .B(\UART_RXFF/n236 ), 
        .C(\UART_RXFF/n237 ), .D(\UART_RXFF/n235 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n239 ) );
  notech_mux4 \UART_RXFF/U248  ( .A(\UART_RXFF/iFIFOMem[32][8] ), .B(
        \UART_RXFF/iFIFOMem[34][8] ), .C(\UART_RXFF/iFIFOMem[33][8] ), .D(
        \UART_RXFF/iFIFOMem[35][8] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n238 ) );
  notech_mux4 \UART_RXFF/U247  ( .A(\UART_RXFF/iFIFOMem[36][8] ), .B(
        \UART_RXFF/iFIFOMem[38][8] ), .C(\UART_RXFF/iFIFOMem[37][8] ), .D(
        \UART_RXFF/iFIFOMem[39][8] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n237 ) );
  notech_mux4 \UART_RXFF/U246  ( .A(\UART_RXFF/iFIFOMem[40][8] ), .B(
        \UART_RXFF/iFIFOMem[42][8] ), .C(\UART_RXFF/iFIFOMem[41][8] ), .D(
        \UART_RXFF/iFIFOMem[43][8] ), .S0(\UART_RXFF/N13 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n236 ) );
  notech_mux4 \UART_RXFF/U245  ( .A(\UART_RXFF/iFIFOMem[44][8] ), .B(
        \UART_RXFF/iFIFOMem[46][8] ), .C(\UART_RXFF/iFIFOMem[45][8] ), .D(
        \UART_RXFF/iFIFOMem[47][8] ), .S0(\UART_RXFF/n59 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n235 ) );
  notech_mux4 \UART_RXFF/U244  ( .A(\UART_RXFF/n233 ), .B(\UART_RXFF/n231 ), 
        .C(\UART_RXFF/n232 ), .D(\UART_RXFF/n230 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n234 ) );
  notech_mux4 \UART_RXFF/U243  ( .A(\UART_RXFF/iFIFOMem[48][8] ), .B(
        \UART_RXFF/iFIFOMem[50][8] ), .C(\UART_RXFF/iFIFOMem[49][8] ), .D(
        \UART_RXFF/iFIFOMem[51][8] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n233 ) );
  notech_mux4 \UART_RXFF/U242  ( .A(\UART_RXFF/iFIFOMem[52][8] ), .B(
        \UART_RXFF/iFIFOMem[54][8] ), .C(\UART_RXFF/iFIFOMem[53][8] ), .D(
        \UART_RXFF/iFIFOMem[55][8] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n232 ) );
  notech_mux4 \UART_RXFF/U241  ( .A(\UART_RXFF/iFIFOMem[56][8] ), .B(
        \UART_RXFF/iFIFOMem[58][8] ), .C(\UART_RXFF/iFIFOMem[57][8] ), .D(
        \UART_RXFF/iFIFOMem[59][8] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n231 ) );
  notech_mux4 \UART_RXFF/U240  ( .A(\UART_RXFF/iFIFOMem[60][8] ), .B(
        \UART_RXFF/iFIFOMem[62][8] ), .C(\UART_RXFF/iFIFOMem[61][8] ), .D(
        \UART_RXFF/iFIFOMem[63][8] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n230 ) );
  notech_mux4 \UART_RXFF/U239  ( .A(\UART_RXFF/n229 ), .B(\UART_RXFF/n219 ), 
        .C(\UART_RXFF/n224 ), .D(\UART_RXFF/n214 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N126 ) );
  notech_mux4 \UART_RXFF/U238  ( .A(\UART_RXFF/n228 ), .B(\UART_RXFF/n226 ), 
        .C(\UART_RXFF/n227 ), .D(\UART_RXFF/n225 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n229 ) );
  notech_mux4 \UART_RXFF/U237  ( .A(\UART_RXFF/iFIFOMem[0][7] ), .B(
        \UART_RXFF/iFIFOMem[2][7] ), .C(\UART_RXFF/iFIFOMem[1][7] ), .D(
        \UART_RXFF/iFIFOMem[3][7] ), .S0(\UART_RXFF/n56 ), .S1(\UART_RXFF/n67 ), .Z(\UART_RXFF/n228 ) );
  notech_mux4 \UART_RXFF/U236  ( .A(\UART_RXFF/iFIFOMem[4][7] ), .B(
        \UART_RXFF/iFIFOMem[6][7] ), .C(\UART_RXFF/iFIFOMem[5][7] ), .D(
        \UART_RXFF/iFIFOMem[7][7] ), .S0(\UART_RXFF/n57 ), .S1(\UART_RXFF/n67 ), .Z(\UART_RXFF/n227 ) );
  notech_mux4 \UART_RXFF/U235  ( .A(\UART_RXFF/iFIFOMem[8][7] ), .B(
        \UART_RXFF/iFIFOMem[10][7] ), .C(\UART_RXFF/iFIFOMem[9][7] ), .D(
        \UART_RXFF/iFIFOMem[11][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n226 ) );
  notech_mux4 \UART_RXFF/U234  ( .A(\UART_RXFF/iFIFOMem[12][7] ), .B(
        \UART_RXFF/iFIFOMem[14][7] ), .C(\UART_RXFF/iFIFOMem[13][7] ), .D(
        \UART_RXFF/iFIFOMem[15][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n67 ), .Z(\UART_RXFF/n225 ) );
  notech_mux4 \UART_RXFF/U233  ( .A(\UART_RXFF/n223 ), .B(\UART_RXFF/n221 ), 
        .C(\UART_RXFF/n222 ), .D(\UART_RXFF/n220 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n224 ) );
  notech_mux4 \UART_RXFF/U232  ( .A(\UART_RXFF/iFIFOMem[16][7] ), .B(
        \UART_RXFF/iFIFOMem[18][7] ), .C(\UART_RXFF/iFIFOMem[17][7] ), .D(
        \UART_RXFF/iFIFOMem[19][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n223 ) );
  notech_mux4 \UART_RXFF/U231  ( .A(\UART_RXFF/iFIFOMem[20][7] ), .B(
        \UART_RXFF/iFIFOMem[22][7] ), .C(\UART_RXFF/iFIFOMem[21][7] ), .D(
        \UART_RXFF/iFIFOMem[23][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n222 ) );
  notech_mux4 \UART_RXFF/U230  ( .A(\UART_RXFF/iFIFOMem[24][7] ), .B(
        \UART_RXFF/iFIFOMem[26][7] ), .C(\UART_RXFF/iFIFOMem[25][7] ), .D(
        \UART_RXFF/iFIFOMem[27][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n221 ) );
  notech_mux4 \UART_RXFF/U229  ( .A(\UART_RXFF/iFIFOMem[28][7] ), .B(
        \UART_RXFF/iFIFOMem[30][7] ), .C(\UART_RXFF/iFIFOMem[29][7] ), .D(
        \UART_RXFF/iFIFOMem[31][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n220 ) );
  notech_mux4 \UART_RXFF/U228  ( .A(\UART_RXFF/n218 ), .B(\UART_RXFF/n216 ), 
        .C(\UART_RXFF/n217 ), .D(\UART_RXFF/n215 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n219 ) );
  notech_mux4 \UART_RXFF/U227  ( .A(\UART_RXFF/iFIFOMem[32][7] ), .B(
        \UART_RXFF/iFIFOMem[34][7] ), .C(\UART_RXFF/iFIFOMem[33][7] ), .D(
        \UART_RXFF/iFIFOMem[35][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n218 ) );
  notech_mux4 \UART_RXFF/U226  ( .A(\UART_RXFF/iFIFOMem[36][7] ), .B(
        \UART_RXFF/iFIFOMem[38][7] ), .C(\UART_RXFF/iFIFOMem[37][7] ), .D(
        \UART_RXFF/iFIFOMem[39][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n217 ) );
  notech_mux4 \UART_RXFF/U225  ( .A(\UART_RXFF/iFIFOMem[40][7] ), .B(
        \UART_RXFF/iFIFOMem[42][7] ), .C(\UART_RXFF/iFIFOMem[41][7] ), .D(
        \UART_RXFF/iFIFOMem[43][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n216 ) );
  notech_mux4 \UART_RXFF/U224  ( .A(\UART_RXFF/iFIFOMem[44][7] ), .B(
        \UART_RXFF/iFIFOMem[46][7] ), .C(\UART_RXFF/iFIFOMem[45][7] ), .D(
        \UART_RXFF/iFIFOMem[47][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n215 ) );
  notech_mux4 \UART_RXFF/U223  ( .A(\UART_RXFF/n213 ), .B(\UART_RXFF/n211 ), 
        .C(\UART_RXFF/n212 ), .D(\UART_RXFF/n210 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n214 ) );
  notech_mux4 \UART_RXFF/U222  ( .A(\UART_RXFF/iFIFOMem[48][7] ), .B(
        \UART_RXFF/iFIFOMem[50][7] ), .C(\UART_RXFF/iFIFOMem[49][7] ), .D(
        \UART_RXFF/iFIFOMem[51][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n213 ) );
  notech_mux4 \UART_RXFF/U221  ( .A(\UART_RXFF/iFIFOMem[52][7] ), .B(
        \UART_RXFF/iFIFOMem[54][7] ), .C(\UART_RXFF/iFIFOMem[53][7] ), .D(
        \UART_RXFF/iFIFOMem[55][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n212 ) );
  notech_mux4 \UART_RXFF/U220  ( .A(\UART_RXFF/iFIFOMem[56][7] ), .B(
        \UART_RXFF/iFIFOMem[58][7] ), .C(\UART_RXFF/iFIFOMem[57][7] ), .D(
        \UART_RXFF/iFIFOMem[59][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n211 ) );
  notech_mux4 \UART_RXFF/U219  ( .A(\UART_RXFF/iFIFOMem[60][7] ), .B(
        \UART_RXFF/iFIFOMem[62][7] ), .C(\UART_RXFF/iFIFOMem[61][7] ), .D(
        \UART_RXFF/iFIFOMem[63][7] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n210 ) );
  notech_mux4 \UART_RXFF/U218  ( .A(\UART_RXFF/n209 ), .B(\UART_RXFF/n199 ), 
        .C(\UART_RXFF/n204 ), .D(\UART_RXFF/n194 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N127 ) );
  notech_mux4 \UART_RXFF/U217  ( .A(\UART_RXFF/n208 ), .B(\UART_RXFF/n206 ), 
        .C(\UART_RXFF/n207 ), .D(\UART_RXFF/n205 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n209 ) );
  notech_mux4 \UART_RXFF/U216  ( .A(\UART_RXFF/iFIFOMem[0][6] ), .B(
        \UART_RXFF/iFIFOMem[2][6] ), .C(\UART_RXFF/iFIFOMem[1][6] ), .D(
        \UART_RXFF/iFIFOMem[3][6] ), .S0(\UART_RXFF/n58 ), .S1(\UART_RXFF/n66 ), .Z(\UART_RXFF/n208 ) );
  notech_mux4 \UART_RXFF/U215  ( .A(\UART_RXFF/iFIFOMem[4][6] ), .B(
        \UART_RXFF/iFIFOMem[6][6] ), .C(\UART_RXFF/iFIFOMem[5][6] ), .D(
        \UART_RXFF/iFIFOMem[7][6] ), .S0(\UART_RXFF/n58 ), .S1(\UART_RXFF/n66 ), .Z(\UART_RXFF/n207 ) );
  notech_mux4 \UART_RXFF/U214  ( .A(\UART_RXFF/iFIFOMem[8][6] ), .B(
        \UART_RXFF/iFIFOMem[10][6] ), .C(\UART_RXFF/iFIFOMem[9][6] ), .D(
        \UART_RXFF/iFIFOMem[11][6] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n206 ) );
  notech_mux4 \UART_RXFF/U213  ( .A(\UART_RXFF/iFIFOMem[12][6] ), .B(
        \UART_RXFF/iFIFOMem[14][6] ), .C(\UART_RXFF/iFIFOMem[13][6] ), .D(
        \UART_RXFF/iFIFOMem[15][6] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n205 ) );
  notech_mux4 \UART_RXFF/U212  ( .A(\UART_RXFF/n203 ), .B(\UART_RXFF/n201 ), 
        .C(\UART_RXFF/n202 ), .D(\UART_RXFF/n200 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n204 ) );
  notech_mux4 \UART_RXFF/U211  ( .A(\UART_RXFF/iFIFOMem[16][6] ), .B(
        \UART_RXFF/iFIFOMem[18][6] ), .C(\UART_RXFF/iFIFOMem[17][6] ), .D(
        \UART_RXFF/iFIFOMem[19][6] ), .S0(\UART_RXFF/n58 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n203 ) );
  notech_mux4 \UART_RXFF/U210  ( .A(\UART_RXFF/iFIFOMem[20][6] ), .B(
        \UART_RXFF/iFIFOMem[22][6] ), .C(\UART_RXFF/iFIFOMem[21][6] ), .D(
        \UART_RXFF/iFIFOMem[23][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n66 ), .Z(\UART_RXFF/n202 ) );
  notech_mux4 \UART_RXFF/U209  ( .A(\UART_RXFF/iFIFOMem[24][6] ), .B(
        \UART_RXFF/iFIFOMem[26][6] ), .C(\UART_RXFF/iFIFOMem[25][6] ), .D(
        \UART_RXFF/iFIFOMem[27][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n201 ) );
  notech_mux4 \UART_RXFF/U208  ( .A(\UART_RXFF/iFIFOMem[28][6] ), .B(
        \UART_RXFF/iFIFOMem[30][6] ), .C(\UART_RXFF/iFIFOMem[29][6] ), .D(
        \UART_RXFF/iFIFOMem[31][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n200 ) );
  notech_mux4 \UART_RXFF/U207  ( .A(\UART_RXFF/n198 ), .B(\UART_RXFF/n196 ), 
        .C(\UART_RXFF/n197 ), .D(\UART_RXFF/n195 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n199 ) );
  notech_mux4 \UART_RXFF/U206  ( .A(\UART_RXFF/iFIFOMem[32][6] ), .B(
        \UART_RXFF/iFIFOMem[34][6] ), .C(\UART_RXFF/iFIFOMem[33][6] ), .D(
        \UART_RXFF/iFIFOMem[35][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n198 ) );
  notech_mux4 \UART_RXFF/U205  ( .A(\UART_RXFF/iFIFOMem[36][6] ), .B(
        \UART_RXFF/iFIFOMem[38][6] ), .C(\UART_RXFF/iFIFOMem[37][6] ), .D(
        \UART_RXFF/iFIFOMem[39][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n197 ) );
  notech_mux4 \UART_RXFF/U204  ( .A(\UART_RXFF/iFIFOMem[40][6] ), .B(
        \UART_RXFF/iFIFOMem[42][6] ), .C(\UART_RXFF/iFIFOMem[41][6] ), .D(
        \UART_RXFF/iFIFOMem[43][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n196 ) );
  notech_mux4 \UART_RXFF/U203  ( .A(\UART_RXFF/iFIFOMem[44][6] ), .B(
        \UART_RXFF/iFIFOMem[46][6] ), .C(\UART_RXFF/iFIFOMem[45][6] ), .D(
        \UART_RXFF/iFIFOMem[47][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n195 ) );
  notech_mux4 \UART_RXFF/U202  ( .A(\UART_RXFF/n193 ), .B(\UART_RXFF/n191 ), 
        .C(\UART_RXFF/n192 ), .D(\UART_RXFF/n190 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n194 ) );
  notech_mux4 \UART_RXFF/U201  ( .A(\UART_RXFF/iFIFOMem[48][6] ), .B(
        \UART_RXFF/iFIFOMem[50][6] ), .C(\UART_RXFF/iFIFOMem[49][6] ), .D(
        \UART_RXFF/iFIFOMem[51][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n193 ) );
  notech_mux4 \UART_RXFF/U200  ( .A(\UART_RXFF/iFIFOMem[52][6] ), .B(
        \UART_RXFF/iFIFOMem[54][6] ), .C(\UART_RXFF/iFIFOMem[53][6] ), .D(
        \UART_RXFF/iFIFOMem[55][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n192 ) );
  notech_mux4 \UART_RXFF/U199  ( .A(\UART_RXFF/iFIFOMem[56][6] ), .B(
        \UART_RXFF/iFIFOMem[58][6] ), .C(\UART_RXFF/iFIFOMem[57][6] ), .D(
        \UART_RXFF/iFIFOMem[59][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n191 ) );
  notech_mux4 \UART_RXFF/U198  ( .A(\UART_RXFF/iFIFOMem[60][6] ), .B(
        \UART_RXFF/iFIFOMem[62][6] ), .C(\UART_RXFF/iFIFOMem[61][6] ), .D(
        \UART_RXFF/iFIFOMem[63][6] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n190 ) );
  notech_mux4 \UART_RXFF/U197  ( .A(\UART_RXFF/n189 ), .B(\UART_RXFF/n179 ), 
        .C(\UART_RXFF/n184 ), .D(\UART_RXFF/n174 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N128 ) );
  notech_mux4 \UART_RXFF/U196  ( .A(\UART_RXFF/n188 ), .B(\UART_RXFF/n186 ), 
        .C(\UART_RXFF/n187 ), .D(\UART_RXFF/n185 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n189 ) );
  notech_mux4 \UART_RXFF/U195  ( .A(\UART_RXFF/iFIFOMem[0][5] ), .B(
        \UART_RXFF/iFIFOMem[2][5] ), .C(\UART_RXFF/iFIFOMem[1][5] ), .D(
        \UART_RXFF/iFIFOMem[3][5] ), .S0(\UART_RXFF/n57 ), .S1(\UART_RXFF/n65 ), .Z(\UART_RXFF/n188 ) );
  notech_mux4 \UART_RXFF/U194  ( .A(\UART_RXFF/iFIFOMem[4][5] ), .B(
        \UART_RXFF/iFIFOMem[6][5] ), .C(\UART_RXFF/iFIFOMem[5][5] ), .D(
        \UART_RXFF/iFIFOMem[7][5] ), .S0(\UART_RXFF/n57 ), .S1(\UART_RXFF/n65 ), .Z(\UART_RXFF/n187 ) );
  notech_mux4 \UART_RXFF/U193  ( .A(\UART_RXFF/iFIFOMem[8][5] ), .B(
        \UART_RXFF/iFIFOMem[10][5] ), .C(\UART_RXFF/iFIFOMem[9][5] ), .D(
        \UART_RXFF/iFIFOMem[11][5] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n186 ) );
  notech_mux4 \UART_RXFF/U192  ( .A(\UART_RXFF/iFIFOMem[12][5] ), .B(
        \UART_RXFF/iFIFOMem[14][5] ), .C(\UART_RXFF/iFIFOMem[13][5] ), .D(
        \UART_RXFF/iFIFOMem[15][5] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n185 ) );
  notech_mux4 \UART_RXFF/U191  ( .A(\UART_RXFF/n183 ), .B(\UART_RXFF/n181 ), 
        .C(\UART_RXFF/n182 ), .D(\UART_RXFF/n180 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n184 ) );
  notech_mux4 \UART_RXFF/U190  ( .A(\UART_RXFF/iFIFOMem[16][5] ), .B(
        \UART_RXFF/iFIFOMem[18][5] ), .C(\UART_RXFF/iFIFOMem[17][5] ), .D(
        \UART_RXFF/iFIFOMem[19][5] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n183 ) );
  notech_mux4 \UART_RXFF/U189  ( .A(\UART_RXFF/iFIFOMem[20][5] ), .B(
        \UART_RXFF/iFIFOMem[22][5] ), .C(\UART_RXFF/iFIFOMem[21][5] ), .D(
        \UART_RXFF/iFIFOMem[23][5] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n182 ) );
  notech_mux4 \UART_RXFF/U188  ( .A(\UART_RXFF/iFIFOMem[24][5] ), .B(
        \UART_RXFF/iFIFOMem[26][5] ), .C(\UART_RXFF/iFIFOMem[25][5] ), .D(
        \UART_RXFF/iFIFOMem[27][5] ), .S0(\UART_RXFF/n57 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n181 ) );
  notech_mux4 \UART_RXFF/U187  ( .A(\UART_RXFF/iFIFOMem[28][5] ), .B(
        \UART_RXFF/iFIFOMem[30][5] ), .C(\UART_RXFF/iFIFOMem[29][5] ), .D(
        \UART_RXFF/iFIFOMem[31][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n65 ), .Z(\UART_RXFF/n180 ) );
  notech_mux4 \UART_RXFF/U186  ( .A(\UART_RXFF/n178 ), .B(\UART_RXFF/n176 ), 
        .C(\UART_RXFF/n177 ), .D(\UART_RXFF/n175 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n179 ) );
  notech_mux4 \UART_RXFF/U185  ( .A(\UART_RXFF/iFIFOMem[32][5] ), .B(
        \UART_RXFF/iFIFOMem[34][5] ), .C(\UART_RXFF/iFIFOMem[33][5] ), .D(
        \UART_RXFF/iFIFOMem[35][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n178 ) );
  notech_mux4 \UART_RXFF/U184  ( .A(\UART_RXFF/iFIFOMem[36][5] ), .B(
        \UART_RXFF/iFIFOMem[38][5] ), .C(\UART_RXFF/iFIFOMem[37][5] ), .D(
        \UART_RXFF/iFIFOMem[39][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n177 ) );
  notech_mux4 \UART_RXFF/U183  ( .A(\UART_RXFF/iFIFOMem[40][5] ), .B(
        \UART_RXFF/iFIFOMem[42][5] ), .C(\UART_RXFF/iFIFOMem[41][5] ), .D(
        \UART_RXFF/iFIFOMem[43][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n176 ) );
  notech_mux4 \UART_RXFF/U182  ( .A(\UART_RXFF/iFIFOMem[44][5] ), .B(
        \UART_RXFF/iFIFOMem[46][5] ), .C(\UART_RXFF/iFIFOMem[45][5] ), .D(
        \UART_RXFF/iFIFOMem[47][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n175 ) );
  notech_mux4 \UART_RXFF/U181  ( .A(\UART_RXFF/n173 ), .B(\UART_RXFF/n171 ), 
        .C(\UART_RXFF/n172 ), .D(\UART_RXFF/n170 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n174 ) );
  notech_mux4 \UART_RXFF/U180  ( .A(\UART_RXFF/iFIFOMem[48][5] ), .B(
        \UART_RXFF/iFIFOMem[50][5] ), .C(\UART_RXFF/iFIFOMem[49][5] ), .D(
        \UART_RXFF/iFIFOMem[51][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n173 ) );
  notech_mux4 \UART_RXFF/U179  ( .A(\UART_RXFF/iFIFOMem[52][5] ), .B(
        \UART_RXFF/iFIFOMem[54][5] ), .C(\UART_RXFF/iFIFOMem[53][5] ), .D(
        \UART_RXFF/iFIFOMem[55][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n172 ) );
  notech_mux4 \UART_RXFF/U178  ( .A(\UART_RXFF/iFIFOMem[56][5] ), .B(
        \UART_RXFF/iFIFOMem[58][5] ), .C(\UART_RXFF/iFIFOMem[57][5] ), .D(
        \UART_RXFF/iFIFOMem[59][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n171 ) );
  notech_mux4 \UART_RXFF/U177  ( .A(\UART_RXFF/iFIFOMem[60][5] ), .B(
        \UART_RXFF/iFIFOMem[62][5] ), .C(\UART_RXFF/iFIFOMem[61][5] ), .D(
        \UART_RXFF/iFIFOMem[63][5] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n170 ) );
  notech_mux4 \UART_RXFF/U176  ( .A(\UART_RXFF/n169 ), .B(\UART_RXFF/n159 ), 
        .C(\UART_RXFF/n164 ), .D(\UART_RXFF/n154 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N129 ) );
  notech_mux4 \UART_RXFF/U175  ( .A(\UART_RXFF/n168 ), .B(\UART_RXFF/n166 ), 
        .C(\UART_RXFF/n167 ), .D(\UART_RXFF/n165 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n169 ) );
  notech_mux4 \UART_RXFF/U174  ( .A(\UART_RXFF/iFIFOMem[0][4] ), .B(
        \UART_RXFF/iFIFOMem[2][4] ), .C(\UART_RXFF/iFIFOMem[1][4] ), .D(
        \UART_RXFF/iFIFOMem[3][4] ), .S0(\UART_RXFF/n56 ), .S1(\UART_RXFF/n64 ), .Z(\UART_RXFF/n168 ) );
  notech_mux4 \UART_RXFF/U173  ( .A(\UART_RXFF/iFIFOMem[4][4] ), .B(
        \UART_RXFF/iFIFOMem[6][4] ), .C(\UART_RXFF/iFIFOMem[5][4] ), .D(
        \UART_RXFF/iFIFOMem[7][4] ), .S0(\UART_RXFF/n56 ), .S1(\UART_RXFF/n64 ), .Z(\UART_RXFF/n167 ) );
  notech_mux4 \UART_RXFF/U172  ( .A(\UART_RXFF/iFIFOMem[8][4] ), .B(
        \UART_RXFF/iFIFOMem[10][4] ), .C(\UART_RXFF/iFIFOMem[9][4] ), .D(
        \UART_RXFF/iFIFOMem[11][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n166 ) );
  notech_mux4 \UART_RXFF/U171  ( .A(\UART_RXFF/iFIFOMem[12][4] ), .B(
        \UART_RXFF/iFIFOMem[14][4] ), .C(\UART_RXFF/iFIFOMem[13][4] ), .D(
        \UART_RXFF/iFIFOMem[15][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n165 ) );
  notech_mux4 \UART_RXFF/U170  ( .A(\UART_RXFF/n163 ), .B(\UART_RXFF/n161 ), 
        .C(\UART_RXFF/n162 ), .D(\UART_RXFF/n160 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n164 ) );
  notech_mux4 \UART_RXFF/U169  ( .A(\UART_RXFF/iFIFOMem[16][4] ), .B(
        \UART_RXFF/iFIFOMem[18][4] ), .C(\UART_RXFF/iFIFOMem[17][4] ), .D(
        \UART_RXFF/iFIFOMem[19][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n163 ) );
  notech_mux4 \UART_RXFF/U168  ( .A(\UART_RXFF/iFIFOMem[20][4] ), .B(
        \UART_RXFF/iFIFOMem[22][4] ), .C(\UART_RXFF/iFIFOMem[21][4] ), .D(
        \UART_RXFF/iFIFOMem[23][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n162 ) );
  notech_mux4 \UART_RXFF/U167  ( .A(\UART_RXFF/iFIFOMem[24][4] ), .B(
        \UART_RXFF/iFIFOMem[26][4] ), .C(\UART_RXFF/iFIFOMem[25][4] ), .D(
        \UART_RXFF/iFIFOMem[27][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n161 ) );
  notech_mux4 \UART_RXFF/U166  ( .A(\UART_RXFF/iFIFOMem[28][4] ), .B(
        \UART_RXFF/iFIFOMem[30][4] ), .C(\UART_RXFF/iFIFOMem[29][4] ), .D(
        \UART_RXFF/iFIFOMem[31][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n160 ) );
  notech_mux4 \UART_RXFF/U165  ( .A(\UART_RXFF/n158 ), .B(\UART_RXFF/n156 ), 
        .C(\UART_RXFF/n157 ), .D(\UART_RXFF/n155 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n159 ) );
  notech_mux4 \UART_RXFF/U164  ( .A(\UART_RXFF/iFIFOMem[32][4] ), .B(
        \UART_RXFF/iFIFOMem[34][4] ), .C(\UART_RXFF/iFIFOMem[33][4] ), .D(
        \UART_RXFF/iFIFOMem[35][4] ), .S0(\UART_RXFF/n56 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n158 ) );
  notech_mux4 \UART_RXFF/U163  ( .A(\UART_RXFF/iFIFOMem[36][4] ), .B(
        \UART_RXFF/iFIFOMem[38][4] ), .C(\UART_RXFF/iFIFOMem[37][4] ), .D(
        \UART_RXFF/iFIFOMem[39][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n64 ), .Z(\UART_RXFF/n157 ) );
  notech_mux4 \UART_RXFF/U162  ( .A(\UART_RXFF/iFIFOMem[40][4] ), .B(
        \UART_RXFF/iFIFOMem[42][4] ), .C(\UART_RXFF/iFIFOMem[41][4] ), .D(
        \UART_RXFF/iFIFOMem[43][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n156 ) );
  notech_mux4 \UART_RXFF/U161  ( .A(\UART_RXFF/iFIFOMem[44][4] ), .B(
        \UART_RXFF/iFIFOMem[46][4] ), .C(\UART_RXFF/iFIFOMem[45][4] ), .D(
        \UART_RXFF/iFIFOMem[47][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n155 ) );
  notech_mux4 \UART_RXFF/U160  ( .A(\UART_RXFF/n153 ), .B(\UART_RXFF/n151 ), 
        .C(\UART_RXFF/n152 ), .D(\UART_RXFF/n150 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n154 ) );
  notech_mux4 \UART_RXFF/U159  ( .A(\UART_RXFF/iFIFOMem[48][4] ), .B(
        \UART_RXFF/iFIFOMem[50][4] ), .C(\UART_RXFF/iFIFOMem[49][4] ), .D(
        \UART_RXFF/iFIFOMem[51][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n153 ) );
  notech_mux4 \UART_RXFF/U158  ( .A(\UART_RXFF/iFIFOMem[52][4] ), .B(
        \UART_RXFF/iFIFOMem[54][4] ), .C(\UART_RXFF/iFIFOMem[53][4] ), .D(
        \UART_RXFF/iFIFOMem[55][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n152 ) );
  notech_mux4 \UART_RXFF/U157  ( .A(\UART_RXFF/iFIFOMem[56][4] ), .B(
        \UART_RXFF/iFIFOMem[58][4] ), .C(\UART_RXFF/iFIFOMem[57][4] ), .D(
        \UART_RXFF/iFIFOMem[59][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n151 ) );
  notech_mux4 \UART_RXFF/U156  ( .A(\UART_RXFF/iFIFOMem[60][4] ), .B(
        \UART_RXFF/iFIFOMem[62][4] ), .C(\UART_RXFF/iFIFOMem[61][4] ), .D(
        \UART_RXFF/iFIFOMem[63][4] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n150 ) );
  notech_mux4 \UART_RXFF/U155  ( .A(\UART_RXFF/n149 ), .B(\UART_RXFF/n139 ), 
        .C(\UART_RXFF/n144 ), .D(\UART_RXFF/n134 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N130 ) );
  notech_mux4 \UART_RXFF/U154  ( .A(\UART_RXFF/n148 ), .B(\UART_RXFF/n146 ), 
        .C(\UART_RXFF/n147 ), .D(\UART_RXFF/n145 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n149 ) );
  notech_mux4 \UART_RXFF/U153  ( .A(\UART_RXFF/iFIFOMem[0][3] ), .B(
        \UART_RXFF/iFIFOMem[2][3] ), .C(\UART_RXFF/iFIFOMem[1][3] ), .D(
        \UART_RXFF/iFIFOMem[3][3] ), .S0(\UART_RXFF/n55 ), .S1(\UART_RXFF/n63 ), .Z(\UART_RXFF/n148 ) );
  notech_mux4 \UART_RXFF/U152  ( .A(\UART_RXFF/iFIFOMem[4][3] ), .B(
        \UART_RXFF/iFIFOMem[6][3] ), .C(\UART_RXFF/iFIFOMem[5][3] ), .D(
        \UART_RXFF/iFIFOMem[7][3] ), .S0(\UART_RXFF/n55 ), .S1(\UART_RXFF/n63 ), .Z(\UART_RXFF/n147 ) );
  notech_mux4 \UART_RXFF/U151  ( .A(\UART_RXFF/iFIFOMem[8][3] ), .B(
        \UART_RXFF/iFIFOMem[10][3] ), .C(\UART_RXFF/iFIFOMem[9][3] ), .D(
        \UART_RXFF/iFIFOMem[11][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n146 ) );
  notech_mux4 \UART_RXFF/U150  ( .A(\UART_RXFF/iFIFOMem[12][3] ), .B(
        \UART_RXFF/iFIFOMem[14][3] ), .C(\UART_RXFF/iFIFOMem[13][3] ), .D(
        \UART_RXFF/iFIFOMem[15][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n145 ) );
  notech_mux4 \UART_RXFF/U149  ( .A(\UART_RXFF/n143 ), .B(\UART_RXFF/n141 ), 
        .C(\UART_RXFF/n142 ), .D(\UART_RXFF/n140 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n144 ) );
  notech_mux4 \UART_RXFF/U148  ( .A(\UART_RXFF/iFIFOMem[16][3] ), .B(
        \UART_RXFF/iFIFOMem[18][3] ), .C(\UART_RXFF/iFIFOMem[17][3] ), .D(
        \UART_RXFF/iFIFOMem[19][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n143 ) );
  notech_mux4 \UART_RXFF/U147  ( .A(\UART_RXFF/iFIFOMem[20][3] ), .B(
        \UART_RXFF/iFIFOMem[22][3] ), .C(\UART_RXFF/iFIFOMem[21][3] ), .D(
        \UART_RXFF/iFIFOMem[23][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n142 ) );
  notech_mux4 \UART_RXFF/U146  ( .A(\UART_RXFF/iFIFOMem[24][3] ), .B(
        \UART_RXFF/iFIFOMem[26][3] ), .C(\UART_RXFF/iFIFOMem[25][3] ), .D(
        \UART_RXFF/iFIFOMem[27][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n141 ) );
  notech_mux4 \UART_RXFF/U145  ( .A(\UART_RXFF/iFIFOMem[28][3] ), .B(
        \UART_RXFF/iFIFOMem[30][3] ), .C(\UART_RXFF/iFIFOMem[29][3] ), .D(
        \UART_RXFF/iFIFOMem[31][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n140 ) );
  notech_mux4 \UART_RXFF/U144  ( .A(\UART_RXFF/n138 ), .B(\UART_RXFF/n136 ), 
        .C(\UART_RXFF/n137 ), .D(\UART_RXFF/n135 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n139 ) );
  notech_mux4 \UART_RXFF/U143  ( .A(\UART_RXFF/iFIFOMem[32][3] ), .B(
        \UART_RXFF/iFIFOMem[34][3] ), .C(\UART_RXFF/iFIFOMem[33][3] ), .D(
        \UART_RXFF/iFIFOMem[35][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n138 ) );
  notech_mux4 \UART_RXFF/U142  ( .A(\UART_RXFF/iFIFOMem[36][3] ), .B(
        \UART_RXFF/iFIFOMem[38][3] ), .C(\UART_RXFF/iFIFOMem[37][3] ), .D(
        \UART_RXFF/iFIFOMem[39][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n137 ) );
  notech_mux4 \UART_RXFF/U141  ( .A(\UART_RXFF/iFIFOMem[40][3] ), .B(
        \UART_RXFF/iFIFOMem[42][3] ), .C(\UART_RXFF/iFIFOMem[41][3] ), .D(
        \UART_RXFF/iFIFOMem[43][3] ), .S0(\UART_RXFF/n55 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n136 ) );
  notech_mux4 \UART_RXFF/U140  ( .A(\UART_RXFF/iFIFOMem[44][3] ), .B(
        \UART_RXFF/iFIFOMem[46][3] ), .C(\UART_RXFF/iFIFOMem[45][3] ), .D(
        \UART_RXFF/iFIFOMem[47][3] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n63 ), .Z(\UART_RXFF/n135 ) );
  notech_mux4 \UART_RXFF/U139  ( .A(\UART_RXFF/n133 ), .B(\UART_RXFF/n131 ), 
        .C(\UART_RXFF/n132 ), .D(\UART_RXFF/n130 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n134 ) );
  notech_mux4 \UART_RXFF/U138  ( .A(\UART_RXFF/iFIFOMem[48][3] ), .B(
        \UART_RXFF/iFIFOMem[50][3] ), .C(\UART_RXFF/iFIFOMem[49][3] ), .D(
        \UART_RXFF/iFIFOMem[51][3] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n133 ) );
  notech_mux4 \UART_RXFF/U137  ( .A(\UART_RXFF/iFIFOMem[52][3] ), .B(
        \UART_RXFF/iFIFOMem[54][3] ), .C(\UART_RXFF/iFIFOMem[53][3] ), .D(
        \UART_RXFF/iFIFOMem[55][3] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n132 ) );
  notech_mux4 \UART_RXFF/U136  ( .A(\UART_RXFF/iFIFOMem[56][3] ), .B(
        \UART_RXFF/iFIFOMem[58][3] ), .C(\UART_RXFF/iFIFOMem[57][3] ), .D(
        \UART_RXFF/iFIFOMem[59][3] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n131 ) );
  notech_mux4 \UART_RXFF/U135  ( .A(\UART_RXFF/iFIFOMem[60][3] ), .B(
        \UART_RXFF/iFIFOMem[62][3] ), .C(\UART_RXFF/iFIFOMem[61][3] ), .D(
        \UART_RXFF/iFIFOMem[63][3] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n130 ) );
  notech_mux4 \UART_RXFF/U134  ( .A(\UART_RXFF/n129 ), .B(\UART_RXFF/n119 ), 
        .C(\UART_RXFF/n124 ), .D(\UART_RXFF/n114 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N131 ) );
  notech_mux4 \UART_RXFF/U133  ( .A(\UART_RXFF/n128 ), .B(\UART_RXFF/n126 ), 
        .C(\UART_RXFF/n127 ), .D(\UART_RXFF/n125 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n129 ) );
  notech_mux4 \UART_RXFF/U132  ( .A(\UART_RXFF/iFIFOMem[0][2] ), .B(
        \UART_RXFF/iFIFOMem[2][2] ), .C(\UART_RXFF/iFIFOMem[1][2] ), .D(
        \UART_RXFF/iFIFOMem[3][2] ), .S0(\UART_RXFF/n54 ), .S1(\UART_RXFF/n62 ), .Z(\UART_RXFF/n128 ) );
  notech_mux4 \UART_RXFF/U131  ( .A(\UART_RXFF/iFIFOMem[4][2] ), .B(
        \UART_RXFF/iFIFOMem[6][2] ), .C(\UART_RXFF/iFIFOMem[5][2] ), .D(
        \UART_RXFF/iFIFOMem[7][2] ), .S0(\UART_RXFF/n54 ), .S1(\UART_RXFF/n62 ), .Z(\UART_RXFF/n127 ) );
  notech_mux4 \UART_RXFF/U130  ( .A(\UART_RXFF/iFIFOMem[8][2] ), .B(
        \UART_RXFF/iFIFOMem[10][2] ), .C(\UART_RXFF/iFIFOMem[9][2] ), .D(
        \UART_RXFF/iFIFOMem[11][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n126 ) );
  notech_mux4 \UART_RXFF/U129  ( .A(\UART_RXFF/iFIFOMem[12][2] ), .B(
        \UART_RXFF/iFIFOMem[14][2] ), .C(\UART_RXFF/iFIFOMem[13][2] ), .D(
        \UART_RXFF/iFIFOMem[15][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n125 ) );
  notech_mux4 \UART_RXFF/U128  ( .A(\UART_RXFF/n123 ), .B(\UART_RXFF/n121 ), 
        .C(\UART_RXFF/n122 ), .D(\UART_RXFF/n120 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n124 ) );
  notech_mux4 \UART_RXFF/U127  ( .A(\UART_RXFF/iFIFOMem[16][2] ), .B(
        \UART_RXFF/iFIFOMem[18][2] ), .C(\UART_RXFF/iFIFOMem[17][2] ), .D(
        \UART_RXFF/iFIFOMem[19][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n123 ) );
  notech_mux4 \UART_RXFF/U126  ( .A(\UART_RXFF/iFIFOMem[20][2] ), .B(
        \UART_RXFF/iFIFOMem[22][2] ), .C(\UART_RXFF/iFIFOMem[21][2] ), .D(
        \UART_RXFF/iFIFOMem[23][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n122 ) );
  notech_mux4 \UART_RXFF/U125  ( .A(\UART_RXFF/iFIFOMem[24][2] ), .B(
        \UART_RXFF/iFIFOMem[26][2] ), .C(\UART_RXFF/iFIFOMem[25][2] ), .D(
        \UART_RXFF/iFIFOMem[27][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n121 ) );
  notech_mux4 \UART_RXFF/U124  ( .A(\UART_RXFF/iFIFOMem[28][2] ), .B(
        \UART_RXFF/iFIFOMem[30][2] ), .C(\UART_RXFF/iFIFOMem[29][2] ), .D(
        \UART_RXFF/iFIFOMem[31][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n120 ) );
  notech_mux4 \UART_RXFF/U123  ( .A(\UART_RXFF/n118 ), .B(\UART_RXFF/n116 ), 
        .C(\UART_RXFF/n117 ), .D(\UART_RXFF/n115 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n119 ) );
  notech_mux4 \UART_RXFF/U122  ( .A(\UART_RXFF/iFIFOMem[32][2] ), .B(
        \UART_RXFF/iFIFOMem[34][2] ), .C(\UART_RXFF/iFIFOMem[33][2] ), .D(
        \UART_RXFF/iFIFOMem[35][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n118 ) );
  notech_mux4 \UART_RXFF/U121  ( .A(\UART_RXFF/iFIFOMem[36][2] ), .B(
        \UART_RXFF/iFIFOMem[38][2] ), .C(\UART_RXFF/iFIFOMem[37][2] ), .D(
        \UART_RXFF/iFIFOMem[39][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n117 ) );
  notech_mux4 \UART_RXFF/U120  ( .A(\UART_RXFF/iFIFOMem[40][2] ), .B(
        \UART_RXFF/iFIFOMem[42][2] ), .C(\UART_RXFF/iFIFOMem[41][2] ), .D(
        \UART_RXFF/iFIFOMem[43][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n116 ) );
  notech_mux4 \UART_RXFF/U119  ( .A(\UART_RXFF/iFIFOMem[44][2] ), .B(
        \UART_RXFF/iFIFOMem[46][2] ), .C(\UART_RXFF/iFIFOMem[45][2] ), .D(
        \UART_RXFF/iFIFOMem[47][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n115 ) );
  notech_mux4 \UART_RXFF/U118  ( .A(\UART_RXFF/n113 ), .B(\UART_RXFF/n111 ), 
        .C(\UART_RXFF/n112 ), .D(\UART_RXFF/n110 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n114 ) );
  notech_mux4 \UART_RXFF/U117  ( .A(\UART_RXFF/iFIFOMem[48][2] ), .B(
        \UART_RXFF/iFIFOMem[50][2] ), .C(\UART_RXFF/iFIFOMem[49][2] ), .D(
        \UART_RXFF/iFIFOMem[51][2] ), .S0(\UART_RXFF/n54 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n113 ) );
  notech_mux4 \UART_RXFF/U116  ( .A(\UART_RXFF/iFIFOMem[52][2] ), .B(
        \UART_RXFF/iFIFOMem[54][2] ), .C(\UART_RXFF/iFIFOMem[53][2] ), .D(
        \UART_RXFF/iFIFOMem[55][2] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n62 ), .Z(\UART_RXFF/n112 ) );
  notech_mux4 \UART_RXFF/U115  ( .A(\UART_RXFF/iFIFOMem[56][2] ), .B(
        \UART_RXFF/iFIFOMem[58][2] ), .C(\UART_RXFF/iFIFOMem[57][2] ), .D(
        \UART_RXFF/iFIFOMem[59][2] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n111 ) );
  notech_mux4 \UART_RXFF/U114  ( .A(\UART_RXFF/iFIFOMem[60][2] ), .B(
        \UART_RXFF/iFIFOMem[62][2] ), .C(\UART_RXFF/iFIFOMem[61][2] ), .D(
        \UART_RXFF/iFIFOMem[63][2] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n110 ) );
  notech_mux4 \UART_RXFF/U113  ( .A(\UART_RXFF/n109 ), .B(\UART_RXFF/n99 ), 
        .C(\UART_RXFF/n104 ), .D(\UART_RXFF/n94 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N132 ) );
  notech_mux4 \UART_RXFF/U112  ( .A(\UART_RXFF/n108 ), .B(\UART_RXFF/n106 ), 
        .C(\UART_RXFF/n107 ), .D(\UART_RXFF/n105 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n109 ) );
  notech_mux4 \UART_RXFF/U111  ( .A(\UART_RXFF/iFIFOMem[0][1] ), .B(
        \UART_RXFF/iFIFOMem[2][1] ), .C(\UART_RXFF/iFIFOMem[1][1] ), .D(
        \UART_RXFF/iFIFOMem[3][1] ), .S0(\UART_RXFF/n53 ), .S1(\UART_RXFF/n61 ), .Z(\UART_RXFF/n108 ) );
  notech_mux4 \UART_RXFF/U110  ( .A(\UART_RXFF/iFIFOMem[4][1] ), .B(
        \UART_RXFF/iFIFOMem[6][1] ), .C(\UART_RXFF/iFIFOMem[5][1] ), .D(
        \UART_RXFF/iFIFOMem[7][1] ), .S0(\UART_RXFF/n53 ), .S1(\UART_RXFF/n61 ), .Z(\UART_RXFF/n107 ) );
  notech_mux4 \UART_RXFF/U109  ( .A(\UART_RXFF/iFIFOMem[8][1] ), .B(
        \UART_RXFF/iFIFOMem[10][1] ), .C(\UART_RXFF/iFIFOMem[9][1] ), .D(
        \UART_RXFF/iFIFOMem[11][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n106 ) );
  notech_mux4 \UART_RXFF/U108  ( .A(\UART_RXFF/iFIFOMem[12][1] ), .B(
        \UART_RXFF/iFIFOMem[14][1] ), .C(\UART_RXFF/iFIFOMem[13][1] ), .D(
        \UART_RXFF/iFIFOMem[15][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n105 ) );
  notech_mux4 \UART_RXFF/U107  ( .A(\UART_RXFF/n103 ), .B(\UART_RXFF/n101 ), 
        .C(\UART_RXFF/n102 ), .D(\UART_RXFF/n100 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n104 ) );
  notech_mux4 \UART_RXFF/U106  ( .A(\UART_RXFF/iFIFOMem[16][1] ), .B(
        \UART_RXFF/iFIFOMem[18][1] ), .C(\UART_RXFF/iFIFOMem[17][1] ), .D(
        \UART_RXFF/iFIFOMem[19][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n103 ) );
  notech_mux4 \UART_RXFF/U105  ( .A(\UART_RXFF/iFIFOMem[20][1] ), .B(
        \UART_RXFF/iFIFOMem[22][1] ), .C(\UART_RXFF/iFIFOMem[21][1] ), .D(
        \UART_RXFF/iFIFOMem[23][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n102 ) );
  notech_mux4 \UART_RXFF/U104  ( .A(\UART_RXFF/iFIFOMem[24][1] ), .B(
        \UART_RXFF/iFIFOMem[26][1] ), .C(\UART_RXFF/iFIFOMem[25][1] ), .D(
        \UART_RXFF/iFIFOMem[27][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n101 ) );
  notech_mux4 \UART_RXFF/U103  ( .A(\UART_RXFF/iFIFOMem[28][1] ), .B(
        \UART_RXFF/iFIFOMem[30][1] ), .C(\UART_RXFF/iFIFOMem[29][1] ), .D(
        \UART_RXFF/iFIFOMem[31][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n100 ) );
  notech_mux4 \UART_RXFF/U102  ( .A(\UART_RXFF/n98 ), .B(\UART_RXFF/n96 ), .C(
        \UART_RXFF/n97 ), .D(\UART_RXFF/n95 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n99 ) );
  notech_mux4 \UART_RXFF/U101  ( .A(\UART_RXFF/iFIFOMem[32][1] ), .B(
        \UART_RXFF/iFIFOMem[34][1] ), .C(\UART_RXFF/iFIFOMem[33][1] ), .D(
        \UART_RXFF/iFIFOMem[35][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n98 ) );
  notech_mux4 \UART_RXFF/U100  ( .A(\UART_RXFF/iFIFOMem[36][1] ), .B(
        \UART_RXFF/iFIFOMem[38][1] ), .C(\UART_RXFF/iFIFOMem[37][1] ), .D(
        \UART_RXFF/iFIFOMem[39][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n97 ) );
  notech_mux4 \UART_RXFF/U99  ( .A(\UART_RXFF/iFIFOMem[40][1] ), .B(
        \UART_RXFF/iFIFOMem[42][1] ), .C(\UART_RXFF/iFIFOMem[41][1] ), .D(
        \UART_RXFF/iFIFOMem[43][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n96 ) );
  notech_mux4 \UART_RXFF/U98  ( .A(\UART_RXFF/iFIFOMem[44][1] ), .B(
        \UART_RXFF/iFIFOMem[46][1] ), .C(\UART_RXFF/iFIFOMem[45][1] ), .D(
        \UART_RXFF/iFIFOMem[47][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n95 ) );
  notech_mux4 \UART_RXFF/U97  ( .A(\UART_RXFF/n93 ), .B(\UART_RXFF/n91 ), .C(
        \UART_RXFF/n92 ), .D(\UART_RXFF/n90 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n94 ) );
  notech_mux4 \UART_RXFF/U96  ( .A(\UART_RXFF/iFIFOMem[48][1] ), .B(
        \UART_RXFF/iFIFOMem[50][1] ), .C(\UART_RXFF/iFIFOMem[49][1] ), .D(
        \UART_RXFF/iFIFOMem[51][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n93 ) );
  notech_mux4 \UART_RXFF/U95  ( .A(\UART_RXFF/iFIFOMem[52][1] ), .B(
        \UART_RXFF/iFIFOMem[54][1] ), .C(\UART_RXFF/iFIFOMem[53][1] ), .D(
        \UART_RXFF/iFIFOMem[55][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n92 ) );
  notech_mux4 \UART_RXFF/U94  ( .A(\UART_RXFF/iFIFOMem[56][1] ), .B(
        \UART_RXFF/iFIFOMem[58][1] ), .C(\UART_RXFF/iFIFOMem[57][1] ), .D(
        \UART_RXFF/iFIFOMem[59][1] ), .S0(\UART_RXFF/n53 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n91 ) );
  notech_mux4 \UART_RXFF/U93  ( .A(\UART_RXFF/iFIFOMem[60][1] ), .B(
        \UART_RXFF/iFIFOMem[62][1] ), .C(\UART_RXFF/iFIFOMem[61][1] ), .D(
        \UART_RXFF/iFIFOMem[63][1] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/n61 ), .Z(\UART_RXFF/n90 ) );
  notech_mux4 \UART_RXFF/U92  ( .A(\UART_RXFF/n89 ), .B(\UART_RXFF/n79 ), .C(
        \UART_RXFF/n84 ), .D(\UART_RXFF/n74 ), .S0(\UART_RXFF/N17 ), .S1(
        \UART_RXFF/N16 ), .Z(\UART_RXFF/N133 ) );
  notech_mux4 \UART_RXFF/U91  ( .A(\UART_RXFF/n88 ), .B(\UART_RXFF/n86 ), .C(
        \UART_RXFF/n87 ), .D(\UART_RXFF/n85 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n89 ) );
  notech_mux4 \UART_RXFF/U90  ( .A(\UART_RXFF/iFIFOMem[0][0] ), .B(
        \UART_RXFF/iFIFOMem[2][0] ), .C(\UART_RXFF/iFIFOMem[1][0] ), .D(
        \UART_RXFF/iFIFOMem[3][0] ), .S0(\UART_RXFF/n52 ), .S1(\UART_RXFF/N12 ), .Z(\UART_RXFF/n88 ) );
  notech_mux4 \UART_RXFF/U89  ( .A(\UART_RXFF/iFIFOMem[4][0] ), .B(
        \UART_RXFF/iFIFOMem[6][0] ), .C(\UART_RXFF/iFIFOMem[5][0] ), .D(
        \UART_RXFF/iFIFOMem[7][0] ), .S0(\UART_RXFF/n52 ), .S1(\UART_RXFF/N12 ), .Z(\UART_RXFF/n87 ) );
  notech_mux4 \UART_RXFF/U88  ( .A(\UART_RXFF/iFIFOMem[8][0] ), .B(
        \UART_RXFF/iFIFOMem[10][0] ), .C(\UART_RXFF/iFIFOMem[9][0] ), .D(
        \UART_RXFF/iFIFOMem[11][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n86 ) );
  notech_mux4 \UART_RXFF/U87  ( .A(\UART_RXFF/iFIFOMem[12][0] ), .B(
        \UART_RXFF/iFIFOMem[14][0] ), .C(\UART_RXFF/iFIFOMem[13][0] ), .D(
        \UART_RXFF/iFIFOMem[15][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n85 ) );
  notech_mux4 \UART_RXFF/U86  ( .A(\UART_RXFF/n83 ), .B(\UART_RXFF/n81 ), .C(
        \UART_RXFF/n82 ), .D(\UART_RXFF/n80 ), .S0(\UART_RXFF/n50 ), .S1(
        \UART_RXFF/n48 ), .Z(\UART_RXFF/n84 ) );
  notech_mux4 \UART_RXFF/U85  ( .A(\UART_RXFF/iFIFOMem[16][0] ), .B(
        \UART_RXFF/iFIFOMem[18][0] ), .C(\UART_RXFF/iFIFOMem[17][0] ), .D(
        \UART_RXFF/iFIFOMem[19][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n83 ) );
  notech_mux4 \UART_RXFF/U84  ( .A(\UART_RXFF/iFIFOMem[20][0] ), .B(
        \UART_RXFF/iFIFOMem[22][0] ), .C(\UART_RXFF/iFIFOMem[21][0] ), .D(
        \UART_RXFF/iFIFOMem[23][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n82 ) );
  notech_mux4 \UART_RXFF/U83  ( .A(\UART_RXFF/iFIFOMem[24][0] ), .B(
        \UART_RXFF/iFIFOMem[26][0] ), .C(\UART_RXFF/iFIFOMem[25][0] ), .D(
        \UART_RXFF/iFIFOMem[27][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n81 ) );
  notech_mux4 \UART_RXFF/U82  ( .A(\UART_RXFF/iFIFOMem[28][0] ), .B(
        \UART_RXFF/iFIFOMem[30][0] ), .C(\UART_RXFF/iFIFOMem[29][0] ), .D(
        \UART_RXFF/iFIFOMem[31][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n80 ) );
  notech_mux4 \UART_RXFF/U81  ( .A(\UART_RXFF/n78 ), .B(\UART_RXFF/n76 ), .C(
        \UART_RXFF/n77 ), .D(\UART_RXFF/n75 ), .S0(\UART_RXFF/N15 ), .S1(
        \UART_RXFF/n47 ), .Z(\UART_RXFF/n79 ) );
  notech_mux4 \UART_RXFF/U80  ( .A(\UART_RXFF/iFIFOMem[32][0] ), .B(
        \UART_RXFF/iFIFOMem[34][0] ), .C(\UART_RXFF/iFIFOMem[33][0] ), .D(
        \UART_RXFF/iFIFOMem[35][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n78 ) );
  notech_mux4 \UART_RXFF/U79  ( .A(\UART_RXFF/iFIFOMem[36][0] ), .B(
        \UART_RXFF/iFIFOMem[38][0] ), .C(\UART_RXFF/iFIFOMem[37][0] ), .D(
        \UART_RXFF/iFIFOMem[39][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n77 ) );
  notech_mux4 \UART_RXFF/U78  ( .A(\UART_RXFF/iFIFOMem[40][0] ), .B(
        \UART_RXFF/iFIFOMem[42][0] ), .C(\UART_RXFF/iFIFOMem[41][0] ), .D(
        \UART_RXFF/iFIFOMem[43][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n76 ) );
  notech_mux4 \UART_RXFF/U77  ( .A(\UART_RXFF/iFIFOMem[44][0] ), .B(
        \UART_RXFF/iFIFOMem[46][0] ), .C(\UART_RXFF/iFIFOMem[45][0] ), .D(
        \UART_RXFF/iFIFOMem[47][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n75 ) );
  notech_mux4 \UART_RXFF/U76  ( .A(\UART_RXFF/n73 ), .B(\UART_RXFF/n71 ), .C(
        \UART_RXFF/n72 ), .D(\UART_RXFF/n70 ), .S0(\UART_RXFF/n51 ), .S1(
        \UART_RXFF/N14 ), .Z(\UART_RXFF/n74 ) );
  notech_mux4 \UART_RXFF/U75  ( .A(\UART_RXFF/iFIFOMem[48][0] ), .B(
        \UART_RXFF/iFIFOMem[50][0] ), .C(\UART_RXFF/iFIFOMem[49][0] ), .D(
        \UART_RXFF/iFIFOMem[51][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n73 ) );
  notech_mux4 \UART_RXFF/U74  ( .A(\UART_RXFF/iFIFOMem[52][0] ), .B(
        \UART_RXFF/iFIFOMem[54][0] ), .C(\UART_RXFF/iFIFOMem[53][0] ), .D(
        \UART_RXFF/iFIFOMem[55][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n72 ) );
  notech_mux4 \UART_RXFF/U73  ( .A(\UART_RXFF/iFIFOMem[56][0] ), .B(
        \UART_RXFF/iFIFOMem[58][0] ), .C(\UART_RXFF/iFIFOMem[57][0] ), .D(
        \UART_RXFF/iFIFOMem[59][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n71 ) );
  notech_mux4 \UART_RXFF/U72  ( .A(\UART_RXFF/iFIFOMem[60][0] ), .B(
        \UART_RXFF/iFIFOMem[62][0] ), .C(\UART_RXFF/iFIFOMem[61][0] ), .D(
        \UART_RXFF/iFIFOMem[63][0] ), .S0(\UART_RXFF/n52 ), .S1(
        \UART_RXFF/N12 ), .Z(\UART_RXFF/n70 ) );
  notech_inv \UART_RXFF/U71  ( .A(\UART_RXFF/N12 ), .Z(\UART_RXFF/n69 ) );
  notech_inv \UART_RXFF/U70  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n68 ) );
  notech_inv \UART_RXFF/U69  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n67 ) );
  notech_inv \UART_RXFF/U68  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n66 ) );
  notech_inv \UART_RXFF/U67  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n65 ) );
  notech_inv \UART_RXFF/U66  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n64 ) );
  notech_inv \UART_RXFF/U65  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n63 ) );
  notech_inv \UART_RXFF/U64  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n62 ) );
  notech_inv \UART_RXFF/U63  ( .A(\UART_RXFF/n69 ), .Z(\UART_RXFF/n61 ) );
  notech_inv \UART_RXFF/U62  ( .A(\UART_RXFF/N13 ), .Z(\UART_RXFF/n60 ) );
  notech_inv \UART_RXFF/U61  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n59 ) );
  notech_inv \UART_RXFF/U60  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n58 ) );
  notech_inv \UART_RXFF/U59  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n57 ) );
  notech_inv \UART_RXFF/U58  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n56 ) );
  notech_inv \UART_RXFF/U57  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n55 ) );
  notech_inv \UART_RXFF/U56  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n54 ) );
  notech_inv \UART_RXFF/U55  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n53 ) );
  notech_inv \UART_RXFF/U54  ( .A(\UART_RXFF/n60 ), .Z(\UART_RXFF/n52 ) );
  notech_inv \UART_RXFF/U53  ( .A(\UART_RXFF/n49 ), .Z(\UART_RXFF/n51 ) );
  notech_inv \UART_RXFF/U52  ( .A(\UART_RXFF/n49 ), .Z(\UART_RXFF/n50 ) );
  notech_inv \UART_RXFF/U51  ( .A(\UART_RXFF/N15 ), .Z(\UART_RXFF/n49 ) );
  notech_inv \UART_RXFF/U50  ( .A(\UART_RXFF/n46 ), .Z(\UART_RXFF/n48 ) );
  notech_inv \UART_RXFF/U49  ( .A(\UART_RXFF/n46 ), .Z(\UART_RXFF/n47 ) );
  notech_inv \UART_RXFF/U48  ( .A(\UART_RXFF/N14 ), .Z(\UART_RXFF/n46 ) );
  notech_inv \UART_RXFF/U46  ( .A(n535), .Z(\UART_RXFF/n44 ) );
  notech_inv \UART_RXFF/U45  ( .A(n535), .Z(\UART_RXFF/n43 ) );
  notech_inv \UART_RXFF/U44  ( .A(n535), .Z(\UART_RXFF/n42 ) );
  notech_inv \UART_RXFF/U42  ( .A(\UART_RXFF/n37 ), .Z(\UART_RXFF/n40 ) );
  notech_inv \UART_RXFF/U41  ( .A(\UART_RXFF/n37 ), .Z(\UART_RXFF/n39 ) );
  notech_inv \UART_RXFF/U40  ( .A(\UART_RXFF/n37 ), .Z(\UART_RXFF/n38 ) );
  notech_inv \UART_RXFF/U39  ( .A(iRXFIFOD[9]), .Z(\UART_RXFF/n37 ) );
  notech_inv \UART_RXFF/U38  ( .A(\UART_RXFF/n33 ), .Z(\UART_RXFF/n36 ) );
  notech_inv \UART_RXFF/U37  ( .A(\UART_RXFF/n33 ), .Z(\UART_RXFF/n35 ) );
  notech_inv \UART_RXFF/U36  ( .A(\UART_RXFF/n33 ), .Z(\UART_RXFF/n34 ) );
  notech_inv \UART_RXFF/U35  ( .A(iRXFIFOD[8]), .Z(\UART_RXFF/n33 ) );
  notech_inv \UART_RXFF/U34  ( .A(\UART_RXFF/n29 ), .Z(\UART_RXFF/n32 ) );
  notech_inv \UART_RXFF/U33  ( .A(\UART_RXFF/n29 ), .Z(\UART_RXFF/n31 ) );
  notech_inv \UART_RXFF/U32  ( .A(\UART_RXFF/n29 ), .Z(\UART_RXFF/n30 ) );
  notech_inv \UART_RXFF/U31  ( .A(iRXFIFOD[7]), .Z(\UART_RXFF/n29 ) );
  notech_inv \UART_RXFF/U30  ( .A(\UART_RXFF/n25 ), .Z(\UART_RXFF/n28 ) );
  notech_inv \UART_RXFF/U29  ( .A(\UART_RXFF/n25 ), .Z(\UART_RXFF/n27 ) );
  notech_inv \UART_RXFF/U28  ( .A(\UART_RXFF/n25 ), .Z(\UART_RXFF/n26 ) );
  notech_inv \UART_RXFF/U27  ( .A(iRXFIFOD[6]), .Z(\UART_RXFF/n25 ) );
  notech_inv \UART_RXFF/U26  ( .A(\UART_RXFF/n21 ), .Z(\UART_RXFF/n24 ) );
  notech_inv \UART_RXFF/U25  ( .A(\UART_RXFF/n21 ), .Z(\UART_RXFF/n23 ) );
  notech_inv \UART_RXFF/U24  ( .A(\UART_RXFF/n21 ), .Z(\UART_RXFF/n22 ) );
  notech_inv \UART_RXFF/U23  ( .A(iRXFIFOD[5]), .Z(\UART_RXFF/n21 ) );
  notech_inv \UART_RXFF/U22  ( .A(\UART_RXFF/n17 ), .Z(\UART_RXFF/n20 ) );
  notech_inv \UART_RXFF/U21  ( .A(\UART_RXFF/n17 ), .Z(\UART_RXFF/n19 ) );
  notech_inv \UART_RXFF/U20  ( .A(\UART_RXFF/n17 ), .Z(\UART_RXFF/n18 ) );
  notech_inv \UART_RXFF/U19  ( .A(iRXFIFOD[4]), .Z(\UART_RXFF/n17 ) );
  notech_inv \UART_RXFF/U18  ( .A(\UART_RXFF/n13 ), .Z(\UART_RXFF/n16 ) );
  notech_inv \UART_RXFF/U17  ( .A(\UART_RXFF/n13 ), .Z(\UART_RXFF/n15 ) );
  notech_inv \UART_RXFF/U16  ( .A(\UART_RXFF/n13 ), .Z(\UART_RXFF/n14 ) );
  notech_inv \UART_RXFF/U15  ( .A(iRXFIFOD[3]), .Z(\UART_RXFF/n13 ) );
  notech_inv \UART_RXFF/U14  ( .A(\UART_RXFF/n9 ), .Z(\UART_RXFF/n12 ) );
  notech_inv \UART_RXFF/U13  ( .A(\UART_RXFF/n9 ), .Z(\UART_RXFF/n11 ) );
  notech_inv \UART_RXFF/U12  ( .A(\UART_RXFF/n9 ), .Z(\UART_RXFF/n10 ) );
  notech_inv \UART_RXFF/U11  ( .A(iRXFIFOD[2]), .Z(\UART_RXFF/n9 ) );
  notech_inv \UART_RXFF/U10  ( .A(\UART_RXFF/n5 ), .Z(\UART_RXFF/n8 ) );
  notech_inv \UART_RXFF/U9  ( .A(\UART_RXFF/n5 ), .Z(\UART_RXFF/n7 ) );
  notech_inv \UART_RXFF/U8  ( .A(\UART_RXFF/n5 ), .Z(\UART_RXFF/n6 ) );
  notech_inv \UART_RXFF/U7  ( .A(iRXFIFOD[1]), .Z(\UART_RXFF/n5 ) );
  notech_inv \UART_RXFF/U6  ( .A(\UART_RXFF/n1 ), .Z(\UART_RXFF/n4 ) );
  notech_inv \UART_RXFF/U5  ( .A(\UART_RXFF/n1 ), .Z(\UART_RXFF/n3 ) );
  notech_inv \UART_RXFF/U4  ( .A(\UART_RXFF/n1 ), .Z(\UART_RXFF/n2 ) );
  notech_inv \UART_RXFF/U3  ( .A(iRXFIFOD[0]), .Z(\UART_RXFF/n1 ) );
  notech_reg \UART_RXFF/iUSAGE_reg[4]  ( .D(\UART_RXFF/n1686 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(iRXFIFOUsage[4]) );
  notech_reg \UART_RXFF/iUSAGE_reg[3]  ( .D(\UART_RXFF/n1687 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(iRXFIFOUsage[3]) );
  notech_reg \UART_RXFF/iUSAGE_reg[2]  ( .D(\UART_RXFF/n1688 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(iRXFIFOUsage[2]) );
  notech_reg \UART_RXFF/iUSAGE_reg[1]  ( .D(\UART_RXFF/n1689 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(iRXFIFOUsage[1]) );
  notech_reg \UART_RXFF/iUSAGE_reg[5]  ( .D(\UART_RXFF/n1685 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(iRXFIFOUsage[5]) );
  notech_reg \UART_RXFF/iUSAGE_reg[0]  ( .D(\UART_RXFF/n1690 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(\UART_RXFF/USAGE[0] ) );
  notech_reg \UART_RXFF/Q_reg[0]  ( .D(\UART_RXFF/n959 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[0]) );
  notech_reg \UART_RXFF/Q_reg[1]  ( .D(\UART_RXFF/n961 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[1]) );
  notech_reg \UART_RXFF/Q_reg[2]  ( .D(\UART_RXFF/n963 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[2]) );
  notech_reg \UART_RXFF/Q_reg[3]  ( .D(\UART_RXFF/n965 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[3]) );
  notech_reg \UART_RXFF/Q_reg[4]  ( .D(\UART_RXFF/n967 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[4]) );
  notech_reg \UART_RXFF/Q_reg[5]  ( .D(\UART_RXFF/n969 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[5]) );
  notech_reg \UART_RXFF/Q_reg[6]  ( .D(\UART_RXFF/n971 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[6]) );
  notech_reg \UART_RXFF/Q_reg[7]  ( .D(\UART_RXFF/n973 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[7]) );
  notech_reg \UART_RXFF/Q_reg[8]  ( .D(\UART_RXFF/n975 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[8]) );
  notech_reg \UART_RXFF/Q_reg[9]  ( .D(\UART_RXFF/n977 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[9]) );
  notech_reg \UART_RXFF/Q_reg[10]  ( .D(\UART_RXFF/n979 ), .CP(CLK), .CD(1'b1), 
        .Q(iRXFIFOQ[10]) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][0]  ( .D(\UART_RXFF/n1691 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][1]  ( .D(\UART_RXFF/n1692 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][2]  ( .D(\UART_RXFF/n1693 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][3]  ( .D(\UART_RXFF/n1694 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][4]  ( .D(\UART_RXFF/n1695 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][5]  ( .D(\UART_RXFF/n1696 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][6]  ( .D(\UART_RXFF/n1697 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][7]  ( .D(\UART_RXFF/n1698 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][8]  ( .D(\UART_RXFF/n1699 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][9]  ( .D(\UART_RXFF/n1700 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[0][10]  ( .D(\UART_RXFF/n1701 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[0][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][0]  ( .D(\UART_RXFF/n1702 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][1]  ( .D(\UART_RXFF/n1703 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][2]  ( .D(\UART_RXFF/n1704 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][3]  ( .D(\UART_RXFF/n1705 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][4]  ( .D(\UART_RXFF/n1706 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][5]  ( .D(\UART_RXFF/n1707 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][6]  ( .D(\UART_RXFF/n1708 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][7]  ( .D(\UART_RXFF/n1709 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][8]  ( .D(\UART_RXFF/n1710 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][9]  ( .D(\UART_RXFF/n1711 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[1][10]  ( .D(\UART_RXFF/n1712 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[1][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][0]  ( .D(\UART_RXFF/n1713 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][1]  ( .D(\UART_RXFF/n1714 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][2]  ( .D(\UART_RXFF/n1715 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][3]  ( .D(\UART_RXFF/n1716 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][4]  ( .D(\UART_RXFF/n1717 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][5]  ( .D(\UART_RXFF/n1718 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][6]  ( .D(\UART_RXFF/n1719 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][7]  ( .D(\UART_RXFF/n1720 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][8]  ( .D(\UART_RXFF/n1721 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][9]  ( .D(\UART_RXFF/n1722 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[2][10]  ( .D(\UART_RXFF/n1723 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[2][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][0]  ( .D(\UART_RXFF/n1724 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][1]  ( .D(\UART_RXFF/n1725 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][2]  ( .D(\UART_RXFF/n1726 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][3]  ( .D(\UART_RXFF/n1727 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][4]  ( .D(\UART_RXFF/n1728 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][5]  ( .D(\UART_RXFF/n1729 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][6]  ( .D(\UART_RXFF/n1730 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][7]  ( .D(\UART_RXFF/n1731 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][8]  ( .D(\UART_RXFF/n1732 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][9]  ( .D(\UART_RXFF/n1733 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[3][10]  ( .D(\UART_RXFF/n1734 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[3][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][0]  ( .D(\UART_RXFF/n1735 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][1]  ( .D(\UART_RXFF/n1736 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][2]  ( .D(\UART_RXFF/n1737 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][3]  ( .D(\UART_RXFF/n1738 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][4]  ( .D(\UART_RXFF/n1739 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][5]  ( .D(\UART_RXFF/n1740 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][6]  ( .D(\UART_RXFF/n1741 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][7]  ( .D(\UART_RXFF/n1742 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][8]  ( .D(\UART_RXFF/n1743 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][9]  ( .D(\UART_RXFF/n1744 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[4][10]  ( .D(\UART_RXFF/n1745 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[4][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][0]  ( .D(\UART_RXFF/n1746 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][1]  ( .D(\UART_RXFF/n1747 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][2]  ( .D(\UART_RXFF/n1748 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][3]  ( .D(\UART_RXFF/n1749 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][4]  ( .D(\UART_RXFF/n1750 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][5]  ( .D(\UART_RXFF/n1751 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][6]  ( .D(\UART_RXFF/n1752 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][7]  ( .D(\UART_RXFF/n1753 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][8]  ( .D(\UART_RXFF/n1754 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][9]  ( .D(\UART_RXFF/n1755 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[5][10]  ( .D(\UART_RXFF/n1756 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[5][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][0]  ( .D(\UART_RXFF/n1757 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][1]  ( .D(\UART_RXFF/n1758 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][2]  ( .D(\UART_RXFF/n1759 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][3]  ( .D(\UART_RXFF/n1760 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][4]  ( .D(\UART_RXFF/n1761 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][5]  ( .D(\UART_RXFF/n1762 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][6]  ( .D(\UART_RXFF/n1763 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][7]  ( .D(\UART_RXFF/n1764 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][8]  ( .D(\UART_RXFF/n1765 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][9]  ( .D(\UART_RXFF/n1766 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[6][10]  ( .D(\UART_RXFF/n1767 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[6][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][0]  ( .D(\UART_RXFF/n1768 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][1]  ( .D(\UART_RXFF/n1769 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][2]  ( .D(\UART_RXFF/n1770 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][3]  ( .D(\UART_RXFF/n1771 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][4]  ( .D(\UART_RXFF/n1772 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][5]  ( .D(\UART_RXFF/n1773 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][6]  ( .D(\UART_RXFF/n1774 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][7]  ( .D(\UART_RXFF/n1775 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][8]  ( .D(\UART_RXFF/n1776 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][9]  ( .D(\UART_RXFF/n1777 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[7][10]  ( .D(\UART_RXFF/n1778 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[7][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][0]  ( .D(\UART_RXFF/n1779 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][1]  ( .D(\UART_RXFF/n1780 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][2]  ( .D(\UART_RXFF/n1781 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][3]  ( .D(\UART_RXFF/n1782 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][4]  ( .D(\UART_RXFF/n1783 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][5]  ( .D(\UART_RXFF/n1784 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][6]  ( .D(\UART_RXFF/n1785 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][7]  ( .D(\UART_RXFF/n1786 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][8]  ( .D(\UART_RXFF/n1787 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][9]  ( .D(\UART_RXFF/n1788 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[8][10]  ( .D(\UART_RXFF/n1789 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[8][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][0]  ( .D(\UART_RXFF/n1790 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][1]  ( .D(\UART_RXFF/n1791 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][2]  ( .D(\UART_RXFF/n1792 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][3]  ( .D(\UART_RXFF/n1793 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][4]  ( .D(\UART_RXFF/n1794 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][5]  ( .D(\UART_RXFF/n1795 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][6]  ( .D(\UART_RXFF/n1796 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][7]  ( .D(\UART_RXFF/n1797 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][8]  ( .D(\UART_RXFF/n1798 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][9]  ( .D(\UART_RXFF/n1799 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[9][10]  ( .D(\UART_RXFF/n1800 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[9][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][0]  ( .D(\UART_RXFF/n1801 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][1]  ( .D(\UART_RXFF/n1802 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][2]  ( .D(\UART_RXFF/n1803 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][3]  ( .D(\UART_RXFF/n1804 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][4]  ( .D(\UART_RXFF/n1805 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][5]  ( .D(\UART_RXFF/n1806 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][6]  ( .D(\UART_RXFF/n1807 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][7]  ( .D(\UART_RXFF/n1808 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][8]  ( .D(\UART_RXFF/n1809 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][9]  ( .D(\UART_RXFF/n1810 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[10][10]  ( .D(\UART_RXFF/n1811 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[10][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][0]  ( .D(\UART_RXFF/n1812 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][1]  ( .D(\UART_RXFF/n1813 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][2]  ( .D(\UART_RXFF/n1814 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][3]  ( .D(\UART_RXFF/n1815 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][4]  ( .D(\UART_RXFF/n1816 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][5]  ( .D(\UART_RXFF/n1817 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][6]  ( .D(\UART_RXFF/n1818 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][7]  ( .D(\UART_RXFF/n1819 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][8]  ( .D(\UART_RXFF/n1820 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][9]  ( .D(\UART_RXFF/n1821 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[11][10]  ( .D(\UART_RXFF/n1822 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[11][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][0]  ( .D(\UART_RXFF/n1823 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][1]  ( .D(\UART_RXFF/n1824 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][2]  ( .D(\UART_RXFF/n1825 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][3]  ( .D(\UART_RXFF/n1826 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][4]  ( .D(\UART_RXFF/n1827 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][5]  ( .D(\UART_RXFF/n1828 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][6]  ( .D(\UART_RXFF/n1829 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][7]  ( .D(\UART_RXFF/n1830 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][8]  ( .D(\UART_RXFF/n1831 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][9]  ( .D(\UART_RXFF/n1832 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[12][10]  ( .D(\UART_RXFF/n1833 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[12][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][0]  ( .D(\UART_RXFF/n1834 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][1]  ( .D(\UART_RXFF/n1835 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][2]  ( .D(\UART_RXFF/n1836 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][3]  ( .D(\UART_RXFF/n1837 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][4]  ( .D(\UART_RXFF/n1838 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][5]  ( .D(\UART_RXFF/n1839 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][6]  ( .D(\UART_RXFF/n1840 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][7]  ( .D(\UART_RXFF/n1841 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][8]  ( .D(\UART_RXFF/n1842 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][9]  ( .D(\UART_RXFF/n1843 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[13][10]  ( .D(\UART_RXFF/n1844 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[13][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][0]  ( .D(\UART_RXFF/n1845 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][1]  ( .D(\UART_RXFF/n1846 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][2]  ( .D(\UART_RXFF/n1847 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][3]  ( .D(\UART_RXFF/n1848 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][4]  ( .D(\UART_RXFF/n1849 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][5]  ( .D(\UART_RXFF/n1850 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][6]  ( .D(\UART_RXFF/n1851 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][7]  ( .D(\UART_RXFF/n1852 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][8]  ( .D(\UART_RXFF/n1853 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][9]  ( .D(\UART_RXFF/n1854 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[14][10]  ( .D(\UART_RXFF/n1855 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[14][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][0]  ( .D(\UART_RXFF/n1856 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][1]  ( .D(\UART_RXFF/n1857 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][2]  ( .D(\UART_RXFF/n1858 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][3]  ( .D(\UART_RXFF/n1859 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][4]  ( .D(\UART_RXFF/n1860 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][5]  ( .D(\UART_RXFF/n1861 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][6]  ( .D(\UART_RXFF/n1862 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][7]  ( .D(\UART_RXFF/n1863 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][8]  ( .D(\UART_RXFF/n1864 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][9]  ( .D(\UART_RXFF/n1865 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[15][10]  ( .D(\UART_RXFF/n1866 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[15][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][0]  ( .D(\UART_RXFF/n1867 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][1]  ( .D(\UART_RXFF/n1868 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][2]  ( .D(\UART_RXFF/n1869 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][3]  ( .D(\UART_RXFF/n1870 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][4]  ( .D(\UART_RXFF/n1871 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][5]  ( .D(\UART_RXFF/n1872 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][6]  ( .D(\UART_RXFF/n1873 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][7]  ( .D(\UART_RXFF/n1874 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][8]  ( .D(\UART_RXFF/n1875 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][9]  ( .D(\UART_RXFF/n1876 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[16][10]  ( .D(\UART_RXFF/n1877 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[16][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][0]  ( .D(\UART_RXFF/n1878 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][1]  ( .D(\UART_RXFF/n1879 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][2]  ( .D(\UART_RXFF/n1880 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][3]  ( .D(\UART_RXFF/n1881 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][4]  ( .D(\UART_RXFF/n1882 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][5]  ( .D(\UART_RXFF/n1883 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][6]  ( .D(\UART_RXFF/n1884 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][7]  ( .D(\UART_RXFF/n1885 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][8]  ( .D(\UART_RXFF/n1886 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][9]  ( .D(\UART_RXFF/n1887 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[17][10]  ( .D(\UART_RXFF/n1888 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[17][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][0]  ( .D(\UART_RXFF/n1889 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][1]  ( .D(\UART_RXFF/n1890 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][2]  ( .D(\UART_RXFF/n1891 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][3]  ( .D(\UART_RXFF/n1892 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][4]  ( .D(\UART_RXFF/n1893 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][5]  ( .D(\UART_RXFF/n1894 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][6]  ( .D(\UART_RXFF/n1895 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][7]  ( .D(\UART_RXFF/n1896 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][8]  ( .D(\UART_RXFF/n1897 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][9]  ( .D(\UART_RXFF/n1898 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[18][10]  ( .D(\UART_RXFF/n1899 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[18][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][0]  ( .D(\UART_RXFF/n1900 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][1]  ( .D(\UART_RXFF/n1901 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][2]  ( .D(\UART_RXFF/n1902 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][3]  ( .D(\UART_RXFF/n1903 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][4]  ( .D(\UART_RXFF/n1904 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][5]  ( .D(\UART_RXFF/n1905 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][6]  ( .D(\UART_RXFF/n1906 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][7]  ( .D(\UART_RXFF/n1907 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][8]  ( .D(\UART_RXFF/n1908 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][9]  ( .D(\UART_RXFF/n1909 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[19][10]  ( .D(\UART_RXFF/n1910 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[19][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][0]  ( .D(\UART_RXFF/n1911 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][1]  ( .D(\UART_RXFF/n1912 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][2]  ( .D(\UART_RXFF/n1913 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][3]  ( .D(\UART_RXFF/n1914 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][4]  ( .D(\UART_RXFF/n1915 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][5]  ( .D(\UART_RXFF/n1916 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][6]  ( .D(\UART_RXFF/n1917 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][7]  ( .D(\UART_RXFF/n1918 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][8]  ( .D(\UART_RXFF/n1919 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][9]  ( .D(\UART_RXFF/n1920 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[20][10]  ( .D(\UART_RXFF/n1921 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[20][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][0]  ( .D(\UART_RXFF/n1922 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][1]  ( .D(\UART_RXFF/n1923 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][2]  ( .D(\UART_RXFF/n1924 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][3]  ( .D(\UART_RXFF/n1925 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][4]  ( .D(\UART_RXFF/n1926 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][5]  ( .D(\UART_RXFF/n1927 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][6]  ( .D(\UART_RXFF/n1928 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][7]  ( .D(\UART_RXFF/n1929 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][8]  ( .D(\UART_RXFF/n1930 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][9]  ( .D(\UART_RXFF/n1931 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[21][10]  ( .D(\UART_RXFF/n1932 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[21][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][0]  ( .D(\UART_RXFF/n1933 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][1]  ( .D(\UART_RXFF/n1934 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][2]  ( .D(\UART_RXFF/n1935 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][3]  ( .D(\UART_RXFF/n1936 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][4]  ( .D(\UART_RXFF/n1937 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][5]  ( .D(\UART_RXFF/n1938 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][6]  ( .D(\UART_RXFF/n1939 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][7]  ( .D(\UART_RXFF/n1940 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][8]  ( .D(\UART_RXFF/n1941 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][9]  ( .D(\UART_RXFF/n1942 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[22][10]  ( .D(\UART_RXFF/n1943 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[22][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][0]  ( .D(\UART_RXFF/n1944 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][1]  ( .D(\UART_RXFF/n1945 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][2]  ( .D(\UART_RXFF/n1946 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][3]  ( .D(\UART_RXFF/n1947 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][4]  ( .D(\UART_RXFF/n1948 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][5]  ( .D(\UART_RXFF/n1949 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][6]  ( .D(\UART_RXFF/n1950 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][7]  ( .D(\UART_RXFF/n1951 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][8]  ( .D(\UART_RXFF/n1952 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][9]  ( .D(\UART_RXFF/n1953 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[23][10]  ( .D(\UART_RXFF/n1954 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[23][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][0]  ( .D(\UART_RXFF/n1955 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][1]  ( .D(\UART_RXFF/n1956 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][2]  ( .D(\UART_RXFF/n1957 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][3]  ( .D(\UART_RXFF/n1958 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][4]  ( .D(\UART_RXFF/n1959 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][5]  ( .D(\UART_RXFF/n1960 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][6]  ( .D(\UART_RXFF/n1961 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][7]  ( .D(\UART_RXFF/n1962 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][8]  ( .D(\UART_RXFF/n1963 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][9]  ( .D(\UART_RXFF/n1964 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[24][10]  ( .D(\UART_RXFF/n1965 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[24][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][0]  ( .D(\UART_RXFF/n1966 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][1]  ( .D(\UART_RXFF/n1967 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][2]  ( .D(\UART_RXFF/n1968 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][3]  ( .D(\UART_RXFF/n1969 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][4]  ( .D(\UART_RXFF/n1970 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][5]  ( .D(\UART_RXFF/n1971 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][6]  ( .D(\UART_RXFF/n1972 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][7]  ( .D(\UART_RXFF/n1973 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][8]  ( .D(\UART_RXFF/n1974 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][9]  ( .D(\UART_RXFF/n1975 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[25][10]  ( .D(\UART_RXFF/n1976 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[25][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][0]  ( .D(\UART_RXFF/n1977 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][1]  ( .D(\UART_RXFF/n1978 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][2]  ( .D(\UART_RXFF/n1979 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][3]  ( .D(\UART_RXFF/n1980 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][4]  ( .D(\UART_RXFF/n1981 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][5]  ( .D(\UART_RXFF/n1982 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][6]  ( .D(\UART_RXFF/n1983 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][7]  ( .D(\UART_RXFF/n1984 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][8]  ( .D(\UART_RXFF/n1985 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][9]  ( .D(\UART_RXFF/n1986 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[26][10]  ( .D(\UART_RXFF/n1987 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[26][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][0]  ( .D(\UART_RXFF/n1988 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][1]  ( .D(\UART_RXFF/n1989 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][2]  ( .D(\UART_RXFF/n1990 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][3]  ( .D(\UART_RXFF/n1991 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][4]  ( .D(\UART_RXFF/n1992 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][5]  ( .D(\UART_RXFF/n1993 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][6]  ( .D(\UART_RXFF/n1994 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][7]  ( .D(\UART_RXFF/n1995 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][8]  ( .D(\UART_RXFF/n1996 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][9]  ( .D(\UART_RXFF/n1997 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[27][10]  ( .D(\UART_RXFF/n1998 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[27][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][0]  ( .D(\UART_RXFF/n1999 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][1]  ( .D(\UART_RXFF/n2000 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][2]  ( .D(\UART_RXFF/n2001 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][3]  ( .D(\UART_RXFF/n2002 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][4]  ( .D(\UART_RXFF/n2003 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][5]  ( .D(\UART_RXFF/n2004 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][6]  ( .D(\UART_RXFF/n2005 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][7]  ( .D(\UART_RXFF/n2006 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][8]  ( .D(\UART_RXFF/n2007 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][9]  ( .D(\UART_RXFF/n2008 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[28][10]  ( .D(\UART_RXFF/n2009 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[28][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][0]  ( .D(\UART_RXFF/n2010 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][1]  ( .D(\UART_RXFF/n2011 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][2]  ( .D(\UART_RXFF/n2012 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][3]  ( .D(\UART_RXFF/n2013 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][4]  ( .D(\UART_RXFF/n2014 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][5]  ( .D(\UART_RXFF/n2015 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][6]  ( .D(\UART_RXFF/n2016 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][7]  ( .D(\UART_RXFF/n2017 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][8]  ( .D(\UART_RXFF/n2018 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][9]  ( .D(\UART_RXFF/n2019 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[29][10]  ( .D(\UART_RXFF/n2020 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[29][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][0]  ( .D(\UART_RXFF/n2021 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][1]  ( .D(\UART_RXFF/n2022 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][2]  ( .D(\UART_RXFF/n2023 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][3]  ( .D(\UART_RXFF/n2024 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][4]  ( .D(\UART_RXFF/n2025 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][5]  ( .D(\UART_RXFF/n2026 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][6]  ( .D(\UART_RXFF/n2027 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][7]  ( .D(\UART_RXFF/n2028 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][8]  ( .D(\UART_RXFF/n2029 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][9]  ( .D(\UART_RXFF/n2030 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[30][10]  ( .D(\UART_RXFF/n2031 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[30][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][0]  ( .D(\UART_RXFF/n2032 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][1]  ( .D(\UART_RXFF/n2033 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][2]  ( .D(\UART_RXFF/n2034 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][3]  ( .D(\UART_RXFF/n2035 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][4]  ( .D(\UART_RXFF/n2036 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][5]  ( .D(\UART_RXFF/n2037 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][6]  ( .D(\UART_RXFF/n2038 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][7]  ( .D(\UART_RXFF/n2039 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][8]  ( .D(\UART_RXFF/n2040 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][9]  ( .D(\UART_RXFF/n2041 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[31][10]  ( .D(\UART_RXFF/n2042 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[31][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][0]  ( .D(\UART_RXFF/n2043 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][1]  ( .D(\UART_RXFF/n2044 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][2]  ( .D(\UART_RXFF/n2045 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][3]  ( .D(\UART_RXFF/n2046 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][4]  ( .D(\UART_RXFF/n2047 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][5]  ( .D(\UART_RXFF/n2048 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][6]  ( .D(\UART_RXFF/n2049 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][7]  ( .D(\UART_RXFF/n2050 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][8]  ( .D(\UART_RXFF/n2051 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][9]  ( .D(\UART_RXFF/n2052 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[32][10]  ( .D(\UART_RXFF/n2053 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[32][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][0]  ( .D(\UART_RXFF/n2054 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][1]  ( .D(\UART_RXFF/n2055 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][2]  ( .D(\UART_RXFF/n2056 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][3]  ( .D(\UART_RXFF/n2057 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][4]  ( .D(\UART_RXFF/n2058 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][5]  ( .D(\UART_RXFF/n2059 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][6]  ( .D(\UART_RXFF/n2060 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][7]  ( .D(\UART_RXFF/n2061 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][8]  ( .D(\UART_RXFF/n2062 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][9]  ( .D(\UART_RXFF/n2063 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[33][10]  ( .D(\UART_RXFF/n2064 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[33][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][0]  ( .D(\UART_RXFF/n2065 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][1]  ( .D(\UART_RXFF/n2066 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][2]  ( .D(\UART_RXFF/n2067 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][3]  ( .D(\UART_RXFF/n2068 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][4]  ( .D(\UART_RXFF/n2069 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][5]  ( .D(\UART_RXFF/n2070 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][6]  ( .D(\UART_RXFF/n2071 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][7]  ( .D(\UART_RXFF/n2072 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][8]  ( .D(\UART_RXFF/n2073 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][9]  ( .D(\UART_RXFF/n2074 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[34][10]  ( .D(\UART_RXFF/n2075 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[34][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][0]  ( .D(\UART_RXFF/n2076 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][1]  ( .D(\UART_RXFF/n2077 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][2]  ( .D(\UART_RXFF/n2078 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][3]  ( .D(\UART_RXFF/n2079 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][4]  ( .D(\UART_RXFF/n2080 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][5]  ( .D(\UART_RXFF/n2081 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][6]  ( .D(\UART_RXFF/n2082 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][7]  ( .D(\UART_RXFF/n2083 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][8]  ( .D(\UART_RXFF/n2084 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][9]  ( .D(\UART_RXFF/n2085 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[35][10]  ( .D(\UART_RXFF/n2086 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[35][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][0]  ( .D(\UART_RXFF/n2087 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][1]  ( .D(\UART_RXFF/n2088 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][2]  ( .D(\UART_RXFF/n2089 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][3]  ( .D(\UART_RXFF/n2090 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][4]  ( .D(\UART_RXFF/n2091 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][5]  ( .D(\UART_RXFF/n2092 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][6]  ( .D(\UART_RXFF/n2093 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][7]  ( .D(\UART_RXFF/n2094 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][8]  ( .D(\UART_RXFF/n2095 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][9]  ( .D(\UART_RXFF/n2096 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[36][10]  ( .D(\UART_RXFF/n2097 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[36][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][0]  ( .D(\UART_RXFF/n2098 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][1]  ( .D(\UART_RXFF/n2099 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][2]  ( .D(\UART_RXFF/n2100 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][3]  ( .D(\UART_RXFF/n2101 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][4]  ( .D(\UART_RXFF/n2102 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][5]  ( .D(\UART_RXFF/n2103 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][6]  ( .D(\UART_RXFF/n2104 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][7]  ( .D(\UART_RXFF/n2105 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][8]  ( .D(\UART_RXFF/n2106 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][9]  ( .D(\UART_RXFF/n2107 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[37][10]  ( .D(\UART_RXFF/n2108 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[37][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][0]  ( .D(\UART_RXFF/n2109 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][1]  ( .D(\UART_RXFF/n2110 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][2]  ( .D(\UART_RXFF/n2111 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][3]  ( .D(\UART_RXFF/n2112 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][4]  ( .D(\UART_RXFF/n2113 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][5]  ( .D(\UART_RXFF/n2114 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][6]  ( .D(\UART_RXFF/n2115 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][7]  ( .D(\UART_RXFF/n2116 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][8]  ( .D(\UART_RXFF/n2117 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][9]  ( .D(\UART_RXFF/n2118 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[38][10]  ( .D(\UART_RXFF/n2119 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[38][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][0]  ( .D(\UART_RXFF/n2120 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][1]  ( .D(\UART_RXFF/n2121 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][2]  ( .D(\UART_RXFF/n2122 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][3]  ( .D(\UART_RXFF/n2123 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][4]  ( .D(\UART_RXFF/n2124 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][5]  ( .D(\UART_RXFF/n2125 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][6]  ( .D(\UART_RXFF/n2126 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][7]  ( .D(\UART_RXFF/n2127 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][8]  ( .D(\UART_RXFF/n2128 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][9]  ( .D(\UART_RXFF/n2129 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[39][10]  ( .D(\UART_RXFF/n2130 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[39][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][0]  ( .D(\UART_RXFF/n2131 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][1]  ( .D(\UART_RXFF/n2132 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][2]  ( .D(\UART_RXFF/n2133 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][3]  ( .D(\UART_RXFF/n2134 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][4]  ( .D(\UART_RXFF/n2135 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][5]  ( .D(\UART_RXFF/n2136 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][6]  ( .D(\UART_RXFF/n2137 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][7]  ( .D(\UART_RXFF/n2138 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][8]  ( .D(\UART_RXFF/n2139 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][9]  ( .D(\UART_RXFF/n2140 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[40][10]  ( .D(\UART_RXFF/n2141 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[40][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][0]  ( .D(\UART_RXFF/n2142 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][1]  ( .D(\UART_RXFF/n2143 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][2]  ( .D(\UART_RXFF/n2144 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][3]  ( .D(\UART_RXFF/n2145 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][4]  ( .D(\UART_RXFF/n2146 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][5]  ( .D(\UART_RXFF/n2147 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][6]  ( .D(\UART_RXFF/n2148 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][7]  ( .D(\UART_RXFF/n2149 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][8]  ( .D(\UART_RXFF/n2150 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][9]  ( .D(\UART_RXFF/n2151 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[41][10]  ( .D(\UART_RXFF/n2152 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[41][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][0]  ( .D(\UART_RXFF/n2153 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][1]  ( .D(\UART_RXFF/n2154 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][2]  ( .D(\UART_RXFF/n2155 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][3]  ( .D(\UART_RXFF/n2156 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][4]  ( .D(\UART_RXFF/n2157 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][5]  ( .D(\UART_RXFF/n2158 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][6]  ( .D(\UART_RXFF/n2159 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][7]  ( .D(\UART_RXFF/n2160 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][8]  ( .D(\UART_RXFF/n2161 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][9]  ( .D(\UART_RXFF/n2162 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[42][10]  ( .D(\UART_RXFF/n2163 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[42][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][0]  ( .D(\UART_RXFF/n2164 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][1]  ( .D(\UART_RXFF/n2165 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][2]  ( .D(\UART_RXFF/n2166 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][3]  ( .D(\UART_RXFF/n2167 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][4]  ( .D(\UART_RXFF/n2168 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][5]  ( .D(\UART_RXFF/n2169 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][6]  ( .D(\UART_RXFF/n2170 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][7]  ( .D(\UART_RXFF/n2171 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][8]  ( .D(\UART_RXFF/n2172 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][9]  ( .D(\UART_RXFF/n2173 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[43][10]  ( .D(\UART_RXFF/n2174 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[43][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][0]  ( .D(\UART_RXFF/n2175 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][1]  ( .D(\UART_RXFF/n2176 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][2]  ( .D(\UART_RXFF/n2177 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][3]  ( .D(\UART_RXFF/n2178 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][4]  ( .D(\UART_RXFF/n2179 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][5]  ( .D(\UART_RXFF/n2180 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][6]  ( .D(\UART_RXFF/n2181 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][7]  ( .D(\UART_RXFF/n2182 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][8]  ( .D(\UART_RXFF/n2183 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][9]  ( .D(\UART_RXFF/n2184 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[44][10]  ( .D(\UART_RXFF/n2185 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[44][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][0]  ( .D(\UART_RXFF/n2186 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][1]  ( .D(\UART_RXFF/n2187 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][2]  ( .D(\UART_RXFF/n2188 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][3]  ( .D(\UART_RXFF/n2189 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][4]  ( .D(\UART_RXFF/n2190 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][5]  ( .D(\UART_RXFF/n2191 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][6]  ( .D(\UART_RXFF/n2192 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][7]  ( .D(\UART_RXFF/n2193 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][8]  ( .D(\UART_RXFF/n2194 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][9]  ( .D(\UART_RXFF/n2195 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[45][10]  ( .D(\UART_RXFF/n2196 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[45][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][0]  ( .D(\UART_RXFF/n2197 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][1]  ( .D(\UART_RXFF/n2198 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][2]  ( .D(\UART_RXFF/n2199 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][3]  ( .D(\UART_RXFF/n2200 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][4]  ( .D(\UART_RXFF/n2201 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][5]  ( .D(\UART_RXFF/n2202 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][6]  ( .D(\UART_RXFF/n2203 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][7]  ( .D(\UART_RXFF/n2204 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][8]  ( .D(\UART_RXFF/n2205 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][9]  ( .D(\UART_RXFF/n2206 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[46][10]  ( .D(\UART_RXFF/n2207 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[46][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][0]  ( .D(\UART_RXFF/n2208 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][1]  ( .D(\UART_RXFF/n2209 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][2]  ( .D(\UART_RXFF/n2210 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][3]  ( .D(\UART_RXFF/n2211 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][4]  ( .D(\UART_RXFF/n2212 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][5]  ( .D(\UART_RXFF/n2213 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][6]  ( .D(\UART_RXFF/n2214 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][7]  ( .D(\UART_RXFF/n2215 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][8]  ( .D(\UART_RXFF/n2216 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][9]  ( .D(\UART_RXFF/n2217 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[47][10]  ( .D(\UART_RXFF/n2218 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[47][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][0]  ( .D(\UART_RXFF/n2219 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][1]  ( .D(\UART_RXFF/n2220 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][2]  ( .D(\UART_RXFF/n2221 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][3]  ( .D(\UART_RXFF/n2222 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][4]  ( .D(\UART_RXFF/n2223 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][5]  ( .D(\UART_RXFF/n2224 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][6]  ( .D(\UART_RXFF/n2225 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][7]  ( .D(\UART_RXFF/n2226 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][8]  ( .D(\UART_RXFF/n2227 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][9]  ( .D(\UART_RXFF/n2228 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[48][10]  ( .D(\UART_RXFF/n2229 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[48][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][0]  ( .D(\UART_RXFF/n2230 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][1]  ( .D(\UART_RXFF/n2231 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][2]  ( .D(\UART_RXFF/n2232 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][3]  ( .D(\UART_RXFF/n2233 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][4]  ( .D(\UART_RXFF/n2234 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][5]  ( .D(\UART_RXFF/n2235 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][6]  ( .D(\UART_RXFF/n2236 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][7]  ( .D(\UART_RXFF/n2237 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][8]  ( .D(\UART_RXFF/n2238 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][9]  ( .D(\UART_RXFF/n2239 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[49][10]  ( .D(\UART_RXFF/n2240 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[49][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][0]  ( .D(\UART_RXFF/n2241 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][1]  ( .D(\UART_RXFF/n2242 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][2]  ( .D(\UART_RXFF/n2243 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][3]  ( .D(\UART_RXFF/n2244 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][4]  ( .D(\UART_RXFF/n2245 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][5]  ( .D(\UART_RXFF/n2246 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][6]  ( .D(\UART_RXFF/n2247 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][7]  ( .D(\UART_RXFF/n2248 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][8]  ( .D(\UART_RXFF/n2249 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][9]  ( .D(\UART_RXFF/n2250 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[50][10]  ( .D(\UART_RXFF/n2251 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[50][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][0]  ( .D(\UART_RXFF/n2252 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][1]  ( .D(\UART_RXFF/n2253 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][2]  ( .D(\UART_RXFF/n2254 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][3]  ( .D(\UART_RXFF/n2255 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][4]  ( .D(\UART_RXFF/n2256 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][5]  ( .D(\UART_RXFF/n2257 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][6]  ( .D(\UART_RXFF/n2258 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][7]  ( .D(\UART_RXFF/n2259 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][8]  ( .D(\UART_RXFF/n2260 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][9]  ( .D(\UART_RXFF/n2261 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[51][10]  ( .D(\UART_RXFF/n2262 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[51][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][0]  ( .D(\UART_RXFF/n2263 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][1]  ( .D(\UART_RXFF/n2264 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][2]  ( .D(\UART_RXFF/n2265 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][3]  ( .D(\UART_RXFF/n2266 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][4]  ( .D(\UART_RXFF/n2267 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][5]  ( .D(\UART_RXFF/n2268 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][6]  ( .D(\UART_RXFF/n2269 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][7]  ( .D(\UART_RXFF/n2270 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][8]  ( .D(\UART_RXFF/n2271 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][9]  ( .D(\UART_RXFF/n2272 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[52][10]  ( .D(\UART_RXFF/n2273 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[52][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][0]  ( .D(\UART_RXFF/n2274 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][1]  ( .D(\UART_RXFF/n2275 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][2]  ( .D(\UART_RXFF/n2276 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][3]  ( .D(\UART_RXFF/n2277 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][4]  ( .D(\UART_RXFF/n2278 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][5]  ( .D(\UART_RXFF/n2279 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][6]  ( .D(\UART_RXFF/n2280 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][7]  ( .D(\UART_RXFF/n2281 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][8]  ( .D(\UART_RXFF/n2282 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][9]  ( .D(\UART_RXFF/n2283 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[53][10]  ( .D(\UART_RXFF/n2284 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[53][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][0]  ( .D(\UART_RXFF/n2285 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][1]  ( .D(\UART_RXFF/n2286 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][2]  ( .D(\UART_RXFF/n2287 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][3]  ( .D(\UART_RXFF/n2288 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][4]  ( .D(\UART_RXFF/n2289 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][5]  ( .D(\UART_RXFF/n2290 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][6]  ( .D(\UART_RXFF/n2291 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][7]  ( .D(\UART_RXFF/n2292 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][8]  ( .D(\UART_RXFF/n2293 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][9]  ( .D(\UART_RXFF/n2294 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[54][10]  ( .D(\UART_RXFF/n2295 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[54][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][0]  ( .D(\UART_RXFF/n2296 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][1]  ( .D(\UART_RXFF/n2297 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][2]  ( .D(\UART_RXFF/n2298 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][3]  ( .D(\UART_RXFF/n2299 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][4]  ( .D(\UART_RXFF/n2300 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][5]  ( .D(\UART_RXFF/n2301 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][6]  ( .D(\UART_RXFF/n2302 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][7]  ( .D(\UART_RXFF/n2303 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][8]  ( .D(\UART_RXFF/n2304 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][9]  ( .D(\UART_RXFF/n2305 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[55][10]  ( .D(\UART_RXFF/n2306 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[55][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][0]  ( .D(\UART_RXFF/n2307 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][1]  ( .D(\UART_RXFF/n2308 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][2]  ( .D(\UART_RXFF/n2309 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][3]  ( .D(\UART_RXFF/n2310 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][4]  ( .D(\UART_RXFF/n2311 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][5]  ( .D(\UART_RXFF/n2312 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][6]  ( .D(\UART_RXFF/n2313 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][7]  ( .D(\UART_RXFF/n2314 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][8]  ( .D(\UART_RXFF/n2315 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][9]  ( .D(\UART_RXFF/n2316 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[56][10]  ( .D(\UART_RXFF/n2317 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[56][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][0]  ( .D(\UART_RXFF/n2318 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][1]  ( .D(\UART_RXFF/n2319 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][2]  ( .D(\UART_RXFF/n2320 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][3]  ( .D(\UART_RXFF/n2321 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][4]  ( .D(\UART_RXFF/n2322 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][5]  ( .D(\UART_RXFF/n2323 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][6]  ( .D(\UART_RXFF/n2324 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][7]  ( .D(\UART_RXFF/n2325 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][8]  ( .D(\UART_RXFF/n2326 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][9]  ( .D(\UART_RXFF/n2327 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[57][10]  ( .D(\UART_RXFF/n2328 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[57][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][0]  ( .D(\UART_RXFF/n2329 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][1]  ( .D(\UART_RXFF/n2330 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][2]  ( .D(\UART_RXFF/n2331 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][3]  ( .D(\UART_RXFF/n2332 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][4]  ( .D(\UART_RXFF/n2333 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][5]  ( .D(\UART_RXFF/n2334 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][6]  ( .D(\UART_RXFF/n2335 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][7]  ( .D(\UART_RXFF/n2336 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][8]  ( .D(\UART_RXFF/n2337 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][9]  ( .D(\UART_RXFF/n2338 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[58][10]  ( .D(\UART_RXFF/n2339 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[58][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][0]  ( .D(\UART_RXFF/n2340 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][1]  ( .D(\UART_RXFF/n2341 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][2]  ( .D(\UART_RXFF/n2342 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][3]  ( .D(\UART_RXFF/n2343 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][4]  ( .D(\UART_RXFF/n2344 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][5]  ( .D(\UART_RXFF/n2345 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][6]  ( .D(\UART_RXFF/n2346 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][7]  ( .D(\UART_RXFF/n2347 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][8]  ( .D(\UART_RXFF/n2348 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][9]  ( .D(\UART_RXFF/n2349 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[59][10]  ( .D(\UART_RXFF/n2350 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[59][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][0]  ( .D(\UART_RXFF/n2351 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][1]  ( .D(\UART_RXFF/n2352 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][2]  ( .D(\UART_RXFF/n2353 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][3]  ( .D(\UART_RXFF/n2354 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][4]  ( .D(\UART_RXFF/n2355 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][5]  ( .D(\UART_RXFF/n2356 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][6]  ( .D(\UART_RXFF/n2357 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][7]  ( .D(\UART_RXFF/n2358 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][8]  ( .D(\UART_RXFF/n2359 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][9]  ( .D(\UART_RXFF/n2360 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[60][10]  ( .D(\UART_RXFF/n2361 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[60][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][0]  ( .D(\UART_RXFF/n2362 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][1]  ( .D(\UART_RXFF/n2363 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][2]  ( .D(\UART_RXFF/n2364 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][3]  ( .D(\UART_RXFF/n2365 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][4]  ( .D(\UART_RXFF/n2366 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][5]  ( .D(\UART_RXFF/n2367 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][6]  ( .D(\UART_RXFF/n2368 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][7]  ( .D(\UART_RXFF/n2369 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][8]  ( .D(\UART_RXFF/n2370 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][9]  ( .D(\UART_RXFF/n2371 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[61][10]  ( .D(\UART_RXFF/n2372 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[61][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][0]  ( .D(\UART_RXFF/n2373 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][1]  ( .D(\UART_RXFF/n2374 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][2]  ( .D(\UART_RXFF/n2375 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][3]  ( .D(\UART_RXFF/n2376 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][4]  ( .D(\UART_RXFF/n2377 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][5]  ( .D(\UART_RXFF/n2378 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][6]  ( .D(\UART_RXFF/n2379 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][7]  ( .D(\UART_RXFF/n2380 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][8]  ( .D(\UART_RXFF/n2381 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][9]  ( .D(\UART_RXFF/n2382 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[62][10]  ( .D(\UART_RXFF/n2383 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[62][10] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][0]  ( .D(\UART_RXFF/n2384 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][0] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][1]  ( .D(\UART_RXFF/n2385 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][1] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][2]  ( .D(\UART_RXFF/n2386 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][2] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][3]  ( .D(\UART_RXFF/n2387 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][3] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][4]  ( .D(\UART_RXFF/n2388 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][4] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][5]  ( .D(\UART_RXFF/n2389 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][5] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][6]  ( .D(\UART_RXFF/n2390 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][6] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][7]  ( .D(\UART_RXFF/n2391 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][7] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][8]  ( .D(\UART_RXFF/n2392 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][8] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][9]  ( .D(\UART_RXFF/n2393 ), .CP(CLK), 
        .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][9] ) );
  notech_reg \UART_RXFF/iFIFOMem_reg[63][10]  ( .D(\UART_RXFF/n2394 ), .CP(CLK), .CD(1'b1), .Q(\UART_RXFF/iFIFOMem[63][10] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[5]  ( .D(\UART_RXFF/n2401 ), .CP(CLK), 
        .CD(\UART_IS_DSR/n1 ), .Q(\UART_RXFF/iWRAddr[5] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[4]  ( .D(\UART_RXFF/n2402 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_RXFF/iWRAddr[4] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[3]  ( .D(\UART_RXFF/n2403 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_RXFF/iWRAddr[3] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[2]  ( .D(\UART_RXFF/n2404 ), .CP(CLK), 
        .CD(\UART_IS_SIN/n1 ), .Q(\UART_RXFF/iWRAddr[2] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[1]  ( .D(\UART_RXFF/n2405 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_RXFF/iWRAddr[1] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[0]  ( .D(\UART_RXFF/n2406 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_RXFF/iWRAddr[0] ) );
  notech_reg \UART_RXFF/iWRAddr_reg[6]  ( .D(\UART_RXFF/n2407 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_RXFF/iWRAddr[6] ) );
  notech_reg \UART_RXFF/iRDAddr_reg[5]  ( .D(\UART_RXFF/n2395 ), .CP(CLK), 
        .CD(\UART_IS_DSR/n1 ), .Q(\UART_RXFF/N17 ) );
  notech_reg \UART_RXFF/iRDAddr_reg[4]  ( .D(\UART_RXFF/n2396 ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_RXFF/N16 ) );
  notech_reg \UART_RXFF/iRDAddr_reg[3]  ( .D(\UART_RXFF/n2397 ), .CP(CLK), 
        .CD(\UART_IS_SIN/n1 ), .Q(\UART_RXFF/N15 ) );
  notech_reg \UART_RXFF/iRDAddr_reg[2]  ( .D(\UART_RXFF/n2398 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_RXFF/N14 ) );
  notech_reg \UART_RXFF/iRDAddr_reg[1]  ( .D(\UART_RXFF/n2399 ), .CP(CLK), 
        .CD(\UART_IS_DSR/n1 ), .Q(\UART_RXFF/N13 ) );
  notech_reg \UART_RXFF/iRDAddr_reg[6]  ( .D(\UART_RXFF/n2400 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_RXFF/iRDAddr[6] ) );
  notech_reg_set \UART_RXFF/iEMPTY_reg  ( .D(\UART_RXFF/N56 ), .CP(CLK), .SD(
        \UART_IS_DCD/n1 ), .Q(iRXFIFOEmpty) );
  notech_reg \UART_RXFF/iRDAddr_reg[0]  ( .D(\UART_RXFF/n2408 ), .CP(CLK), 
        .CD(\UART_IS_RI/n1 ), .Q(\UART_RXFF/N12 ) );
  notech_xor2 \UART_RXFF/add_73/U1  ( .A(\UART_RXFF/add_73/carry [6]), .B(
        \UART_RXFF/iWRAddr[6] ), .Z(\UART_RXFF/N30 ) );
  notech_ha2 \UART_RXFF/add_73/U1_1_1  ( .A(\UART_RXFF/iWRAddr[1] ), .B(
        \UART_RXFF/iWRAddr[0] ), .CO(\UART_RXFF/add_73/carry [2]), .Z(
        \UART_RXFF/N25 ) );
  notech_ha2 \UART_RXFF/add_73/U1_1_2  ( .A(\UART_RXFF/iWRAddr[2] ), .B(
        \UART_RXFF/add_73/carry [2]), .CO(\UART_RXFF/add_73/carry [3]), .Z(
        \UART_RXFF/N26 ) );
  notech_ha2 \UART_RXFF/add_73/U1_1_3  ( .A(\UART_RXFF/iWRAddr[3] ), .B(
        \UART_RXFF/add_73/carry [3]), .CO(\UART_RXFF/add_73/carry [4]), .Z(
        \UART_RXFF/N27 ) );
  notech_ha2 \UART_RXFF/add_73/U1_1_4  ( .A(\UART_RXFF/iWRAddr[4] ), .B(
        \UART_RXFF/add_73/carry [4]), .CO(\UART_RXFF/add_73/carry [5]), .Z(
        \UART_RXFF/N28 ) );
  notech_ha2 \UART_RXFF/add_73/U1_1_5  ( .A(\UART_RXFF/iWRAddr[5] ), .B(
        \UART_RXFF/add_73/carry [5]), .CO(\UART_RXFF/add_73/carry [6]), .Z(
        \UART_RXFF/N29 ) );
  notech_xor2 \UART_RXFF/add_77/U1  ( .A(\UART_RXFF/add_77/carry [6]), .B(
        \UART_RXFF/iRDAddr[6] ), .Z(\UART_RXFF/N38 ) );
  notech_ha2 \UART_RXFF/add_77/U1_1_1  ( .A(\UART_RXFF/n52 ), .B(
        \UART_RXFF/N12 ), .CO(\UART_RXFF/add_77/carry [2]), .Z(\UART_RXFF/N33 ) );
  notech_ha2 \UART_RXFF/add_77/U1_1_2  ( .A(\UART_RXFF/n48 ), .B(
        \UART_RXFF/add_77/carry [2]), .CO(\UART_RXFF/add_77/carry [3]), .Z(
        \UART_RXFF/N34 ) );
  notech_ha2 \UART_RXFF/add_77/U1_1_3  ( .A(\UART_RXFF/n50 ), .B(
        \UART_RXFF/add_77/carry [3]), .CO(\UART_RXFF/add_77/carry [4]), .Z(
        \UART_RXFF/N35 ) );
  notech_ha2 \UART_RXFF/add_77/U1_1_4  ( .A(\UART_RXFF/N16 ), .B(
        \UART_RXFF/add_77/carry [4]), .CO(\UART_RXFF/add_77/carry [5]), .Z(
        \UART_RXFF/N36 ) );
  notech_ha2 \UART_RXFF/add_77/U1_1_5  ( .A(\UART_RXFF/N17 ), .B(
        \UART_RXFF/add_77/carry [5]), .CO(\UART_RXFF/add_77/carry [6]), .Z(
        \UART_RXFF/N37 ) );
  notech_inv \UART_TX/U95  ( .A(\UART_TX/CState[1] ), .Z(\UART_TX/n28 ) );
  notech_nor2 \UART_TX/U94  ( .A(\UART_TX/n28 ), .B(\UART_TX/CState[2] ), .Z(
        \UART_TX/n15 ) );
  notech_nand2 \UART_TX/U93  ( .A(\UART_TX/n15 ), .B(\UART_TX/CState[0] ), .Z(
        \UART_TX/n40 ) );
  notech_inv \UART_TX/U92  ( .A(\UART_TX/CState[3] ), .Z(\UART_TX/n20 ) );
  notech_or2 \UART_TX/U91  ( .A(\UART_TX/n40 ), .B(\UART_TX/n20 ), .Z(
        \UART_TX/n25 ) );
  notech_nor2 \UART_TX/U90  ( .A(\UART_TX/iLast ), .B(\UART_TX/n25 ), .Z(
        \UART_TX/N127 ) );
  notech_inv \UART_TX/U89  ( .A(\UART_TX/CState[2] ), .Z(\UART_TX/n21 ) );
  notech_inv \UART_TX/U88  ( .A(iTSR[1]), .Z(\UART_TX/n83 ) );
  notech_ao4 \UART_TX/U87  ( .A(\UART_TX/n20 ), .B(\UART_TX/n21 ), .C(
        \UART_TX/n40 ), .D(\UART_TX/n83 ), .Z(\UART_TX/n59 ) );
  notech_nor2 \UART_TX/U86  ( .A(\UART_TX/n21 ), .B(\UART_TX/CState[3] ), .Z(
        \UART_TX/n43 ) );
  notech_and2 \UART_TX/U85  ( .A(\UART_TX/n43 ), .B(\UART_TX/n28 ), .Z(
        \UART_TX/n44 ) );
  notech_nand2 \UART_TX/U84  ( .A(\UART_TX/n44 ), .B(iTSR[3]), .Z(
        \UART_TX/n67 ) );
  notech_inv \UART_TX/U83  ( .A(iTSR[6]), .Z(\UART_TX/n64 ) );
  notech_fa2 \UART_TX/U82  ( .A(iTSR[4]), .B(iTSR[3]), .CI(iTSR[2]), .Z(
        \UART_TX/n84 ) );
  notech_fa2 \UART_TX/U81  ( .A(\UART_TX/n83 ), .B(\UART_TX/n84 ), .CI(iTSR[0]), .Z(\UART_TX/n81 ) );
  notech_xor2 \UART_TX/U80  ( .A(\UART_TX/n81 ), .B(iTSR[5]), .Z(\UART_TX/n80 ) );
  notech_nand2 \UART_TX/U79  ( .A(iTSR[7]), .B(iLCR[0]), .Z(\UART_TX/n82 ) );
  notech_fa2 \UART_TX/U78  ( .A(\UART_TX/n64 ), .B(\UART_TX/n80 ), .CI(
        \UART_TX/n82 ), .Z(\UART_TX/n78 ) );
  notech_inv \UART_TX/U77  ( .A(iLCR[0]), .Z(\UART_TX/n24 ) );
  notech_mux2 \UART_TX/U76  ( .A(\UART_TX/n80 ), .B(\UART_TX/n81 ), .S(
        \UART_TX/n24 ), .Z(\UART_TX/n79 ) );
  notech_inv \UART_TX/U75  ( .A(iLCR[1]), .Z(\UART_TX/n37 ) );
  notech_mux2 \UART_TX/U74  ( .A(\UART_TX/n78 ), .B(\UART_TX/n79 ), .S(
        \UART_TX/n37 ), .Z(\UART_TX/n77 ) );
  notech_nor2 \UART_TX/U73  ( .A(iLCR[5]), .B(\UART_TX/n77 ), .Z(\UART_TX/n76 ) );
  notech_xor2 \UART_TX/U72  ( .A(iLCR[4]), .B(\UART_TX/n76 ), .Z(\UART_TX/n74 ) );
  notech_inv \UART_TX/U71  ( .A(\UART_TX/n43 ), .Z(\UART_TX/n18 ) );
  notech_inv \UART_TX/U70  ( .A(iTSR[4]), .Z(\UART_TX/n75 ) );
  notech_ao4 \UART_TX/U69  ( .A(\UART_TX/n20 ), .B(\UART_TX/n74 ), .C(
        \UART_TX/n18 ), .D(\UART_TX/n75 ), .Z(\UART_TX/n73 ) );
  notech_or2 \UART_TX/U68  ( .A(\UART_TX/n73 ), .B(\UART_TX/n28 ), .Z(
        \UART_TX/n69 ) );
  notech_or2 \UART_TX/U67  ( .A(\UART_TX/n28 ), .B(iTSR[0]), .Z(\UART_TX/n72 )
         );
  notech_nao3 \UART_TX/U66  ( .C(\UART_TX/CState[2] ), .A(\UART_TX/n20 ), .B(
        \UART_TX/n72 ), .Z(\UART_TX/n70 ) );
  notech_nand2 \UART_TX/U65  ( .A(\UART_TX/n44 ), .B(iTSR[2]), .Z(
        \UART_TX/n71 ) );
  notech_and3 \UART_TX/U64  ( .A(\UART_TX/n69 ), .B(\UART_TX/n70 ), .C(
        \UART_TX/n71 ), .Z(\UART_TX/n68 ) );
  notech_inv \UART_TX/U63  ( .A(\UART_TX/CState[0] ), .Z(\UART_TX/n5 ) );
  notech_mux2 \UART_TX/U62  ( .A(\UART_TX/n67 ), .B(\UART_TX/n68 ), .S(
        \UART_TX/n5 ), .Z(\UART_TX/n60 ) );
  notech_and3 \UART_TX/U61  ( .A(\UART_TX/n28 ), .B(\UART_TX/n21 ), .C(
        \UART_TX/CState[3] ), .Z(\UART_TX/n66 ) );
  notech_and2 \UART_TX/U60  ( .A(\UART_TX/n66 ), .B(\UART_TX/CState[0] ), .Z(
        \UART_TX/n51 ) );
  notech_nand2 \UART_TX/U59  ( .A(\UART_TX/n51 ), .B(iTSR[7]), .Z(
        \UART_TX/n62 ) );
  notech_and2 \UART_TX/U58  ( .A(\UART_TX/n66 ), .B(\UART_TX/n5 ), .Z(
        \UART_TX/n22 ) );
  notech_inv \UART_TX/U57  ( .A(\UART_TX/n22 ), .Z(\UART_TX/n50 ) );
  notech_nao3 \UART_TX/U56  ( .C(\UART_TX/n18 ), .A(\UART_TX/CState[1] ), .B(
        \UART_TX/CState[0] ), .Z(\UART_TX/n36 ) );
  notech_inv \UART_TX/U55  ( .A(iTSR[5]), .Z(\UART_TX/n65 ) );
  notech_ao4 \UART_TX/U54  ( .A(\UART_TX/n50 ), .B(\UART_TX/n64 ), .C(
        \UART_TX/n36 ), .D(\UART_TX/n65 ), .Z(\UART_TX/n63 ) );
  notech_and3 \UART_TX/U53  ( .A(\UART_TX/n62 ), .B(\UART_TX/n63 ), .C(
        \UART_TX/n25 ), .Z(\UART_TX/n61 ) );
  notech_and3 \UART_TX/U52  ( .A(\UART_TX/n59 ), .B(\UART_TX/n60 ), .C(
        \UART_TX/n61 ), .Z(\UART_TX/n58 ) );
  notech_nor2 \UART_TX/U51  ( .A(iLCR[6]), .B(\UART_TX/n58 ), .Z(iSOUT) );
  notech_and4 \UART_TX/U50  ( .A(\UART_TX/n37 ), .B(\UART_TX/n24 ), .C(
        \UART_TX/n28 ), .D(\UART_TX/n5 ), .Z(\UART_TX/n57 ) );
  notech_and4 \UART_TX/U49  ( .A(\UART_TX/CState[2] ), .B(\UART_TX/CState[3] ), 
        .C(iLCR[2]), .D(\UART_TX/n57 ), .Z(\UART_TX/n56 ) );
  notech_inv \UART_TX/U48  ( .A(\UART_TX/iTx2 ), .Z(\UART_TX/n53 ) );
  notech_nor2 \UART_TX/U47  ( .A(\UART_TX/n56 ), .B(\UART_TX/n53 ), .Z(
        \UART_TX/n54 ) );
  notech_nor2 \UART_TX/U45  ( .A(\UART_TX/n54 ), .B(\UART_IF_RI/n3 ), .Z(
        \UART_TX/n29 ) );
  notech_inv \UART_TX/U44  ( .A(\UART_TX/n29 ), .Z(\UART_TX/n6 ) );
  notech_or2 \UART_TX/U43  ( .A(\UART_TX/n53 ), .B(iBaudtick2x), .Z(
        \UART_TX/n52 ) );
  notech_nand2 \UART_TX/U42  ( .A(\UART_TX/n6 ), .B(\UART_TX/n52 ), .Z(
        \UART_TX/n87 ) );
  notech_or4 \UART_TX/U41  ( .A(\UART_TX/n28 ), .B(\UART_TX/n18 ), .C(iLCR[1]), 
        .D(iLCR[0]), .Z(\UART_TX/n49 ) );
  notech_inv \UART_TX/U40  ( .A(\UART_TX/n51 ), .Z(\UART_TX/n3 ) );
  notech_and4 \UART_TX/U39  ( .A(\UART_TX/n49 ), .B(\UART_TX/n36 ), .C(
        \UART_TX/n50 ), .D(\UART_TX/n3 ), .Z(\UART_TX/n45 ) );
  notech_or2 \UART_TX/U38  ( .A(\UART_TX/n5 ), .B(iLCR[2]), .Z(\UART_TX/n48 )
         );
  notech_nand2 \UART_TX/U37  ( .A(\UART_TX/n15 ), .B(\UART_TX/n48 ), .Z(
        \UART_TX/n47 ) );
  notech_and2 \UART_TX/U36  ( .A(\UART_TX/n29 ), .B(\UART_TX/n47 ), .Z(
        \UART_TX/n46 ) );
  notech_nao4 \UART_TX/U35  ( .A(\UART_TX/n45 ), .B(\UART_TX/n6 ), .C(
        \UART_TX/n46 ), .D(\UART_TX/n20 ), .Z(\UART_TX/n88 ) );
  notech_inv \UART_TX/U34  ( .A(\UART_TX/n44 ), .Z(\UART_TX/n13 ) );
  notech_nand2 \UART_TX/U33  ( .A(\UART_TX/n37 ), .B(\UART_TX/n24 ), .Z(
        \UART_TX/n42 ) );
  notech_nao3 \UART_TX/U32  ( .C(\UART_TX/CState[0] ), .A(\UART_TX/n42 ), .B(
        \UART_TX/n43 ), .Z(\UART_TX/n8 ) );
  notech_nor2 \UART_TX/U31  ( .A(\UART_TX/n20 ), .B(iLCR[2]), .Z(\UART_TX/n41 ) );
  notech_or2 \UART_TX/U30  ( .A(\UART_TX/n40 ), .B(\UART_TX/n41 ), .Z(
        \UART_TX/n39 ) );
  notech_nand3 \UART_TX/U29  ( .A(\UART_TX/n13 ), .B(\UART_TX/n8 ), .C(
        \UART_TX/n39 ), .Z(\UART_TX/n38 ) );
  notech_mux2 \UART_TX/U28  ( .A(\UART_TX/n38 ), .B(\UART_TX/CState[2] ), .S(
        \UART_TX/n6 ), .Z(\UART_TX/n89 ) );
  notech_nao3 \UART_TX/U27  ( .C(\UART_TX/n37 ), .A(\UART_TX/n24 ), .B(
        \UART_TX/n22 ), .Z(\UART_TX/n32 ) );
  notech_nao3 \UART_TX/U26  ( .C(\UART_TX/n36 ), .A(\UART_TX/n37 ), .B(iLCR[0]), .Z(\UART_TX/n11 ) );
  notech_nand2 \UART_TX/U25  ( .A(\UART_TX/n21 ), .B(\UART_TX/n28 ), .Z(
        \UART_TX/n35 ) );
  notech_and2 \UART_TX/U24  ( .A(\UART_TX/n13 ), .B(\UART_TX/n35 ), .Z(
        \UART_TX/n34 ) );
  notech_or2 \UART_TX/U23  ( .A(\UART_TX/n34 ), .B(\UART_TX/n5 ), .Z(
        \UART_TX/n33 ) );
  notech_and3 \UART_TX/U22  ( .A(\UART_TX/n32 ), .B(\UART_TX/n11 ), .C(
        \UART_TX/n33 ), .Z(\UART_TX/n26 ) );
  notech_nand2 \UART_TX/U21  ( .A(\UART_TX/n18 ), .B(\UART_TX/CState[2] ), .Z(
        \UART_TX/n31 ) );
  notech_nand2 \UART_TX/U20  ( .A(\UART_TX/n31 ), .B(\UART_TX/n5 ), .Z(
        \UART_TX/n30 ) );
  notech_and2 \UART_TX/U19  ( .A(\UART_TX/n29 ), .B(\UART_TX/n30 ), .Z(
        \UART_TX/n27 ) );
  notech_nao4 \UART_TX/U18  ( .A(\UART_TX/n26 ), .B(\UART_TX/n6 ), .C(
        \UART_TX/n27 ), .D(\UART_TX/n28 ), .Z(\UART_TX/n90 ) );
  notech_inv \UART_TX/U17  ( .A(\UART_TX/n25 ), .Z(\UART_TX/n93 ) );
  notech_nao3 \UART_TX/U16  ( .C(iLCR[2]), .A(\UART_TX/n93 ), .B(iTXStart), 
        .Z(\UART_TX/n7 ) );
  notech_nand3 \UART_TX/U15  ( .A(\UART_TX/n24 ), .B(iLCR[3]), .C(iLCR[1]), 
        .Z(\UART_TX/n23 ) );
  notech_nand2 \UART_TX/U14  ( .A(\UART_TX/n22 ), .B(\UART_TX/n23 ), .Z(
        \UART_TX/n9 ) );
  notech_inv \UART_TX/U13  ( .A(iTXStart), .Z(\UART_TX/n16 ) );
  notech_or2 \UART_TX/U12  ( .A(\UART_TX/n21 ), .B(\UART_TX/CState[1] ), .Z(
        \UART_TX/n19 ) );
  notech_mux2 \UART_TX/U11  ( .A(\UART_TX/n19 ), .B(\UART_TX/CState[2] ), .S(
        \UART_TX/n20 ), .Z(\UART_TX/n17 ) );
  notech_ao4 \UART_TX/U10  ( .A(\UART_TX/n16 ), .B(\UART_TX/n17 ), .C(iLCR[3]), 
        .D(\UART_TX/n18 ), .Z(\UART_TX/n14 ) );
  notech_ao3 \UART_TX/U9  ( .A(\UART_TX/n13 ), .B(\UART_TX/n14 ), .C(
        \UART_TX/n15 ), .Z(\UART_TX/n12 ) );
  notech_ao4 \UART_TX/U8  ( .A(iLCR[3]), .B(\UART_TX/n11 ), .C(
        \UART_TX/CState[0] ), .D(\UART_TX/n12 ), .Z(\UART_TX/n10 ) );
  notech_and4 \UART_TX/U7  ( .A(\UART_TX/n7 ), .B(\UART_TX/n8 ), .C(
        \UART_TX/n9 ), .D(\UART_TX/n10 ), .Z(\UART_TX/n4 ) );
  notech_mux2 \UART_TX/U6  ( .A(\UART_TX/n4 ), .B(\UART_TX/n5 ), .S(
        \UART_TX/n6 ), .Z(\UART_TX/n1 ) );
  notech_or2 \UART_TX/U5  ( .A(\UART_TX/n3 ), .B(iLCR[3]), .Z(\UART_TX/n2 ) );
  notech_nand2 \UART_TX/U4  ( .A(\UART_TX/n1 ), .B(\UART_TX/n2 ), .Z(
        \UART_TX/n92 ) );
  notech_reg \UART_TX/iFinished_reg  ( .D(\UART_TX/N127 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(iTXFinished) );
  notech_reg \UART_TX/iLast_reg  ( .D(\UART_TX/n93 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_TX/iLast ) );
  notech_reg \UART_TX/iTx2_reg  ( .D(\UART_TX/n87 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(\UART_TX/iTx2 ) );
  notech_reg \UART_TX/CState_reg[3]  ( .D(\UART_TX/n88 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_TX/CState[3] ) );
  notech_reg \UART_TX/CState_reg[2]  ( .D(\UART_TX/n89 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(\UART_TX/CState[2] ) );
  notech_reg \UART_TX/CState_reg[1]  ( .D(\UART_TX/n90 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_TX/CState[1] ) );
  notech_reg \UART_TX/CState_reg[0]  ( .D(\UART_TX/n92 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(\UART_TX/CState[0] ) );
  notech_inv \UART_RX/U110  ( .A(iRXData[2]), .Z(\UART_RX/n78 ) );
  notech_xor2 \UART_RX/U109  ( .A(iRXData[3]), .B(\UART_RX/n78 ), .Z(
        \UART_RX/n82 ) );
  notech_inv \UART_RX/U108  ( .A(iRXData[1]), .Z(\UART_RX/n77 ) );
  notech_inv \UART_RX/U107  ( .A(iRXData[0]), .Z(\UART_RX/n73 ) );
  notech_xor2 \UART_RX/U106  ( .A(\UART_RX/n77 ), .B(\UART_RX/n73 ), .Z(
        \UART_RX/n83 ) );
  notech_xor2 \UART_RX/U105  ( .A(iRXData[7]), .B(iRXData[6]), .Z(
        \UART_RX/n85 ) );
  notech_fa2 \UART_RX/U104  ( .A(iRXData[5]), .B(\UART_RX/n85 ), .CI(
        iRXData[4]), .Z(\UART_RX/n84 ) );
  notech_fa2 \UART_RX/U103  ( .A(\UART_RX/n82 ), .B(\UART_RX/n83 ), .CI(
        \UART_RX/n84 ), .Z(\UART_RX/n81 ) );
  notech_nor2 \UART_RX/U102  ( .A(iLCR[5]), .B(\UART_RX/n81 ), .Z(
        \UART_RX/n80 ) );
  notech_fa2 \UART_RX/U101  ( .A(iLCR[4]), .B(\UART_RX/n80 ), .CI(
        \UART_RX/iParityReceived ), .Z(\UART_RX/n79 ) );
  notech_inv \UART_RX/U100  ( .A(iLCR[3]), .Z(\UART_RX/n47 ) );
  notech_nor2 \UART_RX/U99  ( .A(\UART_RX/n79 ), .B(\UART_RX/n47 ), .Z(
        \UART_RX/N106 ) );
  notech_inv \UART_RX/U98  ( .A(\UART_RX/CState[0] ), .Z(\UART_RX/n63 ) );
  notech_nao3 \UART_RX/U97  ( .C(\UART_RX/CState[1] ), .A(\UART_RX/CState[2] ), 
        .B(\UART_RX/n63 ), .Z(\UART_RX/n50 ) );
  notech_nor2 \UART_RX/U96  ( .A(\UART_RX/n50 ), .B(\UART_RX/iFStopBit ), .Z(
        iRXFE) );
  notech_ao3 \UART_RX/U95  ( .A(\UART_RX/n77 ), .B(\UART_RX/n78 ), .C(
        iRXData[3]), .Z(\UART_RX/n74 ) );
  notech_or2 \UART_RX/U94  ( .A(\UART_RX/iParityReceived ), .B(iRXData[7]), 
        .Z(\UART_RX/n76 ) );
  notech_nor4 \UART_RX/U93  ( .A(iRXData[4]), .B(iRXData[5]), .C(\UART_RX/n76 ), .D(iRXData[6]), .Z(\UART_RX/n75 ) );
  notech_and4 \UART_RX/U92  ( .A(iRXFE), .B(\UART_RX/n73 ), .C(\UART_RX/n74 ), 
        .D(\UART_RX/n75 ), .Z(iRXBI) );
  notech_nor2 \UART_RX/U91  ( .A(\UART_RX/CState[2] ), .B(\UART_RX/CState[1] ), 
        .Z(\UART_RX/n5 ) );
  notech_nand2 \UART_RX/U90  ( .A(\UART_RX/n5 ), .B(\UART_RX/n63 ), .Z(
        \UART_RX/n61 ) );
  notech_inv \UART_RX/U89  ( .A(\UART_RX/n61 ), .Z(\UART_RX/N75 ) );
  notech_inv \UART_RX/U88  ( .A(\UART_RX/CState[2] ), .Z(\UART_RX/n72 ) );
  notech_nor4 \UART_RX/U87  ( .A(\UART_RX/n72 ), .B(\UART_RX/n63 ), .C(iSIN), 
        .D(\UART_RX/CState[1] ), .Z(\UART_RX/n48 ) );
  notech_inv \UART_RX/U86  ( .A(\UART_RX/iBaudStep ), .Z(\UART_RX/n42 ) );
  notech_and3 \UART_RX/U85  ( .A(\UART_RX/n72 ), .B(\UART_RX/n42 ), .C(
        \UART_RX/CState[0] ), .Z(\UART_RX/n57 ) );
  notech_nand2 \UART_RX/U84  ( .A(\UART_RX/CState[1] ), .B(\UART_RX/n72 ), .Z(
        \UART_RX/n52 ) );
  notech_and2 \UART_RX/U83  ( .A(\UART_RX/iDataCount[1] ), .B(
        \UART_RX/iDataCount[0] ), .Z(\UART_RX/n6 ) );
  notech_and2 \UART_RX/U81  ( .A(\UART_RX/n6 ), .B(\UART_TX/n37 ), .Z(
        \UART_RX/n67 ) );
  notech_inv \UART_RX/U80  ( .A(\UART_RX/iDataCount[0] ), .Z(\UART_RX/n22 ) );
  notech_mux2 \UART_RX/U79  ( .A(\UART_RX/n22 ), .B(iLCR[1]), .S(iLCR[0]), .Z(
        \UART_RX/n68 ) );
  notech_or2 \UART_RX/U78  ( .A(iLCR[0]), .B(iLCR[1]), .Z(\UART_RX/n70 ) );
  notech_inv \UART_RX/U77  ( .A(\UART_RX/iDataCount[1] ), .Z(\UART_RX/n24 ) );
  notech_and2 \UART_RX/U76  ( .A(\UART_RX/n70 ), .B(\UART_RX/n24 ), .Z(
        \UART_RX/n69 ) );
  notech_nor4 \UART_RX/U75  ( .A(\UART_RX/n67 ), .B(\UART_RX/n68 ), .C(
        \UART_RX/iDataCount[3] ), .D(\UART_RX/n69 ), .Z(\UART_RX/n64 ) );
  notech_and2 \UART_RX/U74  ( .A(\UART_RX/n24 ), .B(\UART_RX/n22 ), .Z(
        \UART_RX/n66 ) );
  notech_and4 \UART_RX/U73  ( .A(iLCR[1]), .B(\UART_RX/iDataCount[3] ), .C(
        iLCR[0]), .D(\UART_RX/n66 ), .Z(\UART_RX/n65 ) );
  notech_inv \UART_RX/U72  ( .A(\UART_RX/iDataCount[2] ), .Z(\UART_RX/n31 ) );
  notech_mux2 \UART_RX/U71  ( .A(\UART_RX/n64 ), .B(\UART_RX/n65 ), .S(
        \UART_RX/n31 ), .Z(\UART_RX/n41 ) );
  notech_nao3 \UART_RX/U70  ( .C(\UART_RX/n52 ), .A(\UART_RX/n41 ), .B(
        \UART_RX/n63 ), .Z(\UART_RX/n51 ) );
  notech_nor2 \UART_RX/U69  ( .A(\UART_RX/n51 ), .B(\UART_RX/n47 ), .Z(
        \UART_RX/n58 ) );
  notech_inv \UART_RX/U68  ( .A(\UART_RX/n50 ), .Z(\UART_RX/n62 ) );
  notech_nao4 \UART_RX/U65  ( .A(\UART_RX/iFStopBit ), .B(n680), .C(iSIN), .D(
        \UART_RX/n61 ), .Z(\UART_RX/n59 ) );
  notech_or4 \UART_RX/U64  ( .A(\UART_RX/n48 ), .B(\UART_RX/n57 ), .C(
        \UART_RX/n58 ), .D(\UART_RX/n59 ), .Z(\UART_RX/NState [0]) );
  notech_and2 \UART_RX/U63  ( .A(\UART_RX/n41 ), .B(\UART_RX/n47 ), .Z(
        \UART_RX/n56 ) );
  notech_mux2 \UART_RX/U62  ( .A(\UART_RX/n56 ), .B(\UART_RX/iBaudStep ), .S(
        \UART_RX/CState[0] ), .Z(\UART_RX/n53 ) );
  notech_inv \UART_RX/U61  ( .A(\UART_RX/iFSIN ), .Z(\UART_RX/n43 ) );
  notech_nand2 \UART_RX/U60  ( .A(\UART_RX/iBaudStep ), .B(\UART_RX/n43 ), .Z(
        \UART_RX/n54 ) );
  notech_nand2 \UART_RX/U59  ( .A(\UART_RX/n5 ), .B(\UART_RX/CState[0] ), .Z(
        \UART_RX/n55 ) );
  notech_nao4 \UART_RX/U58  ( .A(\UART_RX/n52 ), .B(\UART_RX/n53 ), .C(
        \UART_RX/n54 ), .D(\UART_RX/n55 ), .Z(\UART_RX/NState [1]) );
  notech_ao3 \UART_RX/U57  ( .A(\UART_RX/CState[0] ), .B(\UART_RX/iBaudStep ), 
        .C(\UART_RX/n52 ), .Z(\UART_RX/n46 ) );
  notech_nao4 \UART_RX/U56  ( .A(\UART_RX/iBaudCount[3] ), .B(\UART_RX/n50 ), 
        .C(iLCR[3]), .D(\UART_RX/n51 ), .Z(\UART_RX/n49 ) );
  notech_or4 \UART_RX/U55  ( .A(iRXFE), .B(\UART_RX/n46 ), .C(\UART_RX/n48 ), 
        .D(\UART_RX/n49 ), .Z(\UART_RX/NState [2]) );
  notech_or2 \UART_RX/U54  ( .A(\UART_RX/N75 ), .B(\UART_RX/iBaudStepD ), .Z(
        \UART_RX/iFilterClear ) );
  notech_and2 \UART_RX/U53  ( .A(iLCR[3]), .B(\UART_RX/iFSIN ), .Z(
        \UART_RX/n44 ) );
  notech_nor2 \UART_RX/U52  ( .A(\UART_RX/n46 ), .B(\UART_RX/n47 ), .Z(
        \UART_RX/n45 ) );
  notech_mux2 \UART_RX/U51  ( .A(\UART_RX/n44 ), .B(\UART_RX/iParityReceived ), 
        .S(\UART_RX/n45 ), .Z(\UART_RX/n105 ) );
  notech_nor2 \UART_RX/U50  ( .A(\UART_RX/n5 ), .B(\UART_RX/n43 ), .Z(
        \UART_RX/n19 ) );
  notech_nor2 \UART_RX/U49  ( .A(\UART_RX/n41 ), .B(\UART_RX/n42 ), .Z(
        \UART_RX/n18 ) );
  notech_and2 \UART_RX/U48  ( .A(\UART_RX/n18 ), .B(\UART_RX/iDataCount[2] ), 
        .Z(\UART_RX/n34 ) );
  notech_and2 \UART_RX/U47  ( .A(\UART_RX/n34 ), .B(\UART_RX/n6 ), .Z(
        \UART_RX/n40 ) );
  notech_nor2 \UART_RX/U46  ( .A(\UART_RX/n40 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n39 ) );
  notech_mux2 \UART_RX/U45  ( .A(\UART_RX/n19 ), .B(iRXData[7]), .S(
        \UART_RX/n39 ), .Z(\UART_RX/n106 ) );
  notech_and2 \UART_RX/U44  ( .A(\UART_RX/iDataCount[1] ), .B(\UART_RX/n22 ), 
        .Z(\UART_RX/n14 ) );
  notech_and2 \UART_RX/U43  ( .A(\UART_RX/n34 ), .B(\UART_RX/n14 ), .Z(
        \UART_RX/n38 ) );
  notech_nor2 \UART_RX/U42  ( .A(\UART_RX/n38 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n37 ) );
  notech_mux2 \UART_RX/U41  ( .A(\UART_RX/n19 ), .B(iRXData[6]), .S(
        \UART_RX/n37 ), .Z(\UART_RX/n107 ) );
  notech_and2 \UART_RX/U40  ( .A(\UART_RX/iDataCount[0] ), .B(\UART_RX/n24 ), 
        .Z(\UART_RX/n15 ) );
  notech_and2 \UART_RX/U39  ( .A(\UART_RX/n34 ), .B(\UART_RX/n15 ), .Z(
        \UART_RX/n36 ) );
  notech_nor2 \UART_RX/U38  ( .A(\UART_RX/n36 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n35 ) );
  notech_mux2 \UART_RX/U37  ( .A(\UART_RX/n19 ), .B(iRXData[5]), .S(
        \UART_RX/n35 ), .Z(\UART_RX/n108 ) );
  notech_and3 \UART_RX/U36  ( .A(\UART_RX/n22 ), .B(\UART_RX/n34 ), .C(
        \UART_RX/n24 ), .Z(\UART_RX/n33 ) );
  notech_nor2 \UART_RX/U35  ( .A(\UART_RX/n33 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n32 ) );
  notech_mux2 \UART_RX/U34  ( .A(\UART_RX/n19 ), .B(iRXData[4]), .S(
        \UART_RX/n32 ), .Z(\UART_RX/n109 ) );
  notech_and2 \UART_RX/U33  ( .A(\UART_RX/n18 ), .B(\UART_RX/n31 ), .Z(
        \UART_RX/n23 ) );
  notech_and2 \UART_RX/U32  ( .A(\UART_RX/n23 ), .B(\UART_RX/n6 ), .Z(
        \UART_RX/n30 ) );
  notech_nor2 \UART_RX/U31  ( .A(\UART_RX/n30 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n29 ) );
  notech_mux2 \UART_RX/U30  ( .A(\UART_RX/n19 ), .B(iRXData[3]), .S(
        \UART_RX/n29 ), .Z(\UART_RX/n110 ) );
  notech_and2 \UART_RX/U29  ( .A(\UART_RX/n23 ), .B(\UART_RX/n14 ), .Z(
        \UART_RX/n28 ) );
  notech_nor2 \UART_RX/U28  ( .A(\UART_RX/n28 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n27 ) );
  notech_mux2 \UART_RX/U27  ( .A(\UART_RX/n19 ), .B(iRXData[2]), .S(
        \UART_RX/n27 ), .Z(\UART_RX/n111 ) );
  notech_and2 \UART_RX/U26  ( .A(\UART_RX/n23 ), .B(\UART_RX/n15 ), .Z(
        \UART_RX/n26 ) );
  notech_nor2 \UART_RX/U25  ( .A(\UART_RX/n26 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n25 ) );
  notech_mux2 \UART_RX/U24  ( .A(\UART_RX/n19 ), .B(iRXData[1]), .S(
        \UART_RX/n25 ), .Z(\UART_RX/n112 ) );
  notech_and3 \UART_RX/U23  ( .A(\UART_RX/n22 ), .B(\UART_RX/n23 ), .C(
        \UART_RX/n24 ), .Z(\UART_RX/n21 ) );
  notech_nor2 \UART_RX/U22  ( .A(\UART_RX/n21 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n20 ) );
  notech_mux2 \UART_RX/U21  ( .A(\UART_RX/n19 ), .B(iRXData[0]), .S(
        \UART_RX/n20 ), .Z(\UART_RX/n113 ) );
  notech_nor2 \UART_RX/U20  ( .A(\UART_RX/n18 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n8 ) );
  notech_or2 \UART_RX/U19  ( .A(\UART_RX/n8 ), .B(\UART_RX/n5 ), .Z(
        \UART_RX/n11 ) );
  notech_inv \UART_RX/U18  ( .A(\UART_RX/n11 ), .Z(\UART_RX/n7 ) );
  notech_and2 \UART_RX/U17  ( .A(\UART_RX/n7 ), .B(\UART_RX/n6 ), .Z(
        \UART_RX/n16 ) );
  notech_nor2 \UART_RX/U16  ( .A(\UART_RX/n5 ), .B(\UART_RX/n6 ), .Z(
        \UART_RX/n17 ) );
  notech_or2 \UART_RX/U15  ( .A(\UART_RX/n8 ), .B(\UART_RX/n17 ), .Z(
        \UART_RX/n3 ) );
  notech_mux2 \UART_RX/U14  ( .A(\UART_RX/n16 ), .B(\UART_RX/n3 ), .S(
        \UART_RX/iDataCount[2] ), .Z(\UART_RX/n114 ) );
  notech_inv \UART_RX/U13  ( .A(\UART_RX/n15 ), .Z(\UART_RX/n12 ) );
  notech_inv \UART_RX/U12  ( .A(\UART_RX/n14 ), .Z(\UART_RX/n13 ) );
  notech_ao4 \UART_RX/U11  ( .A(\UART_RX/n11 ), .B(\UART_RX/n12 ), .C(
        \UART_RX/n5 ), .D(\UART_RX/n13 ), .Z(\UART_RX/n9 ) );
  notech_nand2 \UART_RX/U10  ( .A(\UART_RX/n8 ), .B(\UART_RX/iDataCount[1] ), 
        .Z(\UART_RX/n10 ) );
  notech_nand2 \UART_RX/U9  ( .A(\UART_RX/n9 ), .B(\UART_RX/n10 ), .Z(
        \UART_RX/n115 ) );
  notech_mux2 \UART_RX/U8  ( .A(\UART_RX/n7 ), .B(\UART_RX/n8 ), .S(
        \UART_RX/iDataCount[0] ), .Z(\UART_RX/n116 ) );
  notech_and3 \UART_RX/U7  ( .A(\UART_RX/iDataCount[2] ), .B(\UART_RX/n6 ), 
        .C(\UART_RX/n7 ), .Z(\UART_RX/n1 ) );
  notech_nor2 \UART_RX/U6  ( .A(\UART_RX/n5 ), .B(\UART_RX/iDataCount[2] ), 
        .Z(\UART_RX/n4 ) );
  notech_or2 \UART_RX/U5  ( .A(\UART_RX/n3 ), .B(\UART_RX/n4 ), .Z(
        \UART_RX/n2 ) );
  notech_mux2 \UART_RX/U4  ( .A(\UART_RX/n1 ), .B(\UART_RX/n2 ), .S(
        \UART_RX/iDataCount[3] ), .Z(\UART_RX/n117 ) );
  notech_reg \UART_RX/PE_reg  ( .D(\UART_RX/N106 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(iRXPE) );
  notech_reg \UART_RX/iParityReceived_reg  ( .D(\UART_RX/n105 ), .CP(CLK), 
        .CD(\UART_IF_CTS/n8 ), .Q(\UART_RX/iParityReceived ) );
  notech_reg \UART_RX/iDOUT_reg[7]  ( .D(\UART_RX/n106 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(iRXData[7]) );
  notech_reg \UART_RX/iDOUT_reg[6]  ( .D(\UART_RX/n107 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(iRXData[6]) );
  notech_reg \UART_RX/iDOUT_reg[5]  ( .D(\UART_RX/n108 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(iRXData[5]) );
  notech_reg \UART_RX/iDOUT_reg[4]  ( .D(\UART_RX/n109 ), .CP(CLK), .CD(
        \UART_IS_CTS/n1 ), .Q(iRXData[4]) );
  notech_reg \UART_RX/iDOUT_reg[3]  ( .D(\UART_RX/n110 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(iRXData[3]) );
  notech_reg \UART_RX/iDOUT_reg[2]  ( .D(\UART_RX/n111 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(iRXData[2]) );
  notech_reg \UART_RX/iDOUT_reg[1]  ( .D(\UART_RX/n112 ), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(iRXData[1]) );
  notech_reg \UART_RX/iDOUT_reg[0]  ( .D(\UART_RX/n113 ), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(iRXData[0]) );
  notech_reg \UART_RX/CState_reg[2]  ( .D(\UART_RX/NState [2]), .CP(CLK), .CD(
        \UART_IS_RI/n1 ), .Q(\UART_RX/CState[2] ) );
  notech_reg \UART_RX/iDataCount_reg[2]  ( .D(\UART_RX/n114 ), .CP(CLK), .CD(
        \UART_IS_DCD/n1 ), .Q(\UART_RX/iDataCount[2] ) );
  notech_reg \UART_RX/iDataCount_reg[1]  ( .D(\UART_RX/n115 ), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_RX/iDataCount[1] ) );
  notech_reg \UART_RX/iDataCount_reg[0]  ( .D(\UART_RX/n116 ), .CP(CLK), .CD(
        \UART_IS_SIN/n1 ), .Q(\UART_RX/iDataCount[0] ) );
  notech_reg \UART_RX/iDataCount_reg[3]  ( .D(\UART_RX/n117 ), .CP(CLK), .CD(
        \UART_IF_DSR/n8 ), .Q(\UART_RX/iDataCount[3] ) );
  notech_reg \UART_RX/iBaudStepD_reg  ( .D(\UART_RX/iBaudStep ), .CP(CLK), 
        .CD(\UART_IS_DCD/n1 ), .Q(\UART_RX/iBaudStepD ) );
  notech_reg \UART_RX/CState_reg[1]  ( .D(\UART_RX/NState [1]), .CP(CLK), .CD(
        \UART_IS_DSR/n1 ), .Q(\UART_RX/CState[1] ) );
  notech_reg \UART_RX/CState_reg[0]  ( .D(\UART_RX/NState [0]), .CP(CLK), .CD(
        \UART_IF_CTS/n8 ), .Q(\UART_RX/CState[0] ) );
  notech_inv \UART_RX/RX_BRC/U33  ( .A(\UART_RX/RX_BRC/Q[2] ), .Z(
        \UART_RX/RX_BRC/n12 ) );
  notech_inv \UART_RX/RX_BRC/U29  ( .A(\UART_RX/iBaudCount[3] ), .Z(
        \UART_RX/RX_BRC/n17 ) );
  notech_and3 \UART_RX/RX_BRC/U22  ( .A(\UART_RX/RX_BRC/n22 ), .B(iRCLK), .C(
        \UART_RX/RX_BRC/n23 ), .Z(\UART_RX/RX_BRC/n26 ) );
  notech_nand2 \UART_RX/RX_BRC/U20  ( .A(\UART_RX/RX_BRC/n6 ), .B(
        \UART_RX/n61 ), .Z(\UART_RX/RX_BRC/n7 ) );
  notech_nao4 \UART_RX/RX_BRC/U16  ( .A(\UART_RX/RX_BRC/n6 ), .B(
        \UART_RX/RX_BRC/n17 ), .C(\UART_RX/RX_BRC/n7 ), .D(
        \UART_RX/RX_BRC/n18 ), .Z(\UART_RX/RX_BRC/n27 ) );
  notech_nao4 \UART_RX/RX_BRC/U12  ( .A(\UART_RX/RX_BRC/n6 ), .B(
        \UART_RX/RX_BRC/n12 ), .C(\UART_RX/RX_BRC/n7 ), .D(
        \UART_RX/RX_BRC/n13 ), .Z(\UART_RX/RX_BRC/n28 ) );
  notech_inv \UART_RX/RX_BRC/U11  ( .A(\UART_RX/RX_BRC/Q[1] ), .Z(
        \UART_RX/RX_BRC/n5 ) );
  notech_inv \UART_RX/RX_BRC/U8  ( .A(\UART_RX/RX_BRC/n9 ), .Z(
        \UART_RX/RX_BRC/n8 ) );
  notech_nao4 \UART_RX/RX_BRC/U7  ( .A(\UART_RX/RX_BRC/n5 ), .B(
        \UART_RX/RX_BRC/n6 ), .C(\UART_RX/RX_BRC/n7 ), .D(\UART_RX/RX_BRC/n8 ), 
        .Z(\UART_RX/RX_BRC/n29 ) );
  notech_xor2 \UART_RX/RX_BRC/U6  ( .A(\UART_RX/RX_BRC/Q[0] ), .B(iRCLK), .Z(
        \UART_RX/RX_BRC/n1 ) );
  notech_and2 \UART_RX/RX_BRC/U4  ( .A(\UART_RX/RX_BRC/n1 ), .B(\UART_RX/n61 ), 
        .Z(\UART_RX/RX_BRC/n30 ) );
  notech_reg \UART_RX/RX_BRC/iCounter_reg[4]  ( .D(\UART_RX/RX_BRC/n26 ), .CP(
        CLK), .CD(\UART_IS_DSR/n1 ), .Q(\UART_RX/iBaudStep ) );
  notech_reg \UART_RX/RX_BRC/iCounter_reg[3]  ( .D(\UART_RX/RX_BRC/n27 ), .CP(
        CLK), .CD(\UART_IF_DSR/n8 ), .Q(\UART_RX/iBaudCount[3] ) );
  notech_reg \UART_RX/RX_BRC/iCounter_reg[2]  ( .D(\UART_RX/RX_BRC/n28 ), .CP(
        CLK), .CD(\UART_IF_CTS/n8 ), .Q(\UART_RX/RX_BRC/Q[2] ) );
  notech_reg \UART_RX/RX_BRC/iCounter_reg[1]  ( .D(\UART_RX/RX_BRC/n29 ), .CP(
        CLK), .CD(\UART_IS_RI/n1 ), .Q(\UART_RX/RX_BRC/Q[1] ) );
  notech_reg \UART_RX/RX_BRC/iCounter_reg[0]  ( .D(\UART_RX/RX_BRC/n30 ), .CP(
        CLK), .CD(\UART_IS_DCD/n1 ), .Q(\UART_RX/RX_BRC/Q[0] ) );
  notech_nor2 \UART_RX/RX_MVF/U26  ( .A(\UART_RX/RX_MVF/iCounter[2] ), .B(
        \UART_RX/RX_MVF/iCounter[1] ), .Z(\UART_RX/RX_MVF/n18 ) );
  notech_inv \UART_RX/RX_MVF/U25  ( .A(\UART_RX/RX_MVF/iCounter[3] ), .Z(
        \UART_RX/RX_MVF/n12 ) );
  notech_or2 \UART_RX/RX_MVF/U24  ( .A(\UART_RX/RX_MVF/n18 ), .B(
        \UART_RX/RX_MVF/n12 ), .Z(\UART_RX/RX_MVF/n16 ) );
  notech_nor2 \UART_RX/RX_MVF/U23  ( .A(\UART_RX/RX_MVF/n17 ), .B(
        \UART_RX/iFilterClear ), .Z(\UART_RX/RX_MVF/n21 ) );
  notech_nor2 \UART_RX/RX_MVF/U22  ( .A(\UART_RX/RX_MVF/n15 ), .B(
        \UART_RX/iFilterClear ), .Z(\UART_RX/RX_MVF/n2 ) );
  notech_or2 \UART_RX/RX_MVF/U21  ( .A(\UART_RX/RX_MVF/n2 ), .B(
        \UART_RX/iFilterClear ), .Z(\UART_RX/RX_MVF/n10 ) );
  notech_inv \UART_RX/RX_MVF/U20  ( .A(\UART_RX/RX_MVF/n10 ), .Z(
        \UART_RX/RX_MVF/n1 ) );
  notech_nor2 \UART_RX/RX_MVF/U19  ( .A(\UART_RX/RX_MVF/n1 ), .B(
        \UART_RX/RX_MVF/n2 ), .Z(\UART_RX/RX_MVF/n3 ) );
  notech_nand2 \UART_RX/RX_MVF/U18  ( .A(\UART_RX/RX_MVF/n1 ), .B(
        \UART_RX/RX_MVF/iCounter[0] ), .Z(\UART_RX/RX_MVF/n13 ) );
  notech_nand2 \UART_RX/RX_MVF/U17  ( .A(\UART_RX/RX_MVF/iCounter[2] ), .B(
        \UART_RX/RX_MVF/iCounter[1] ), .Z(\UART_RX/RX_MVF/n14 ) );
  notech_nao4 \UART_RX/RX_MVF/U16  ( .A(\UART_RX/RX_MVF/n3 ), .B(
        \UART_RX/RX_MVF/n12 ), .C(\UART_RX/RX_MVF/n13 ), .D(
        \UART_RX/RX_MVF/n14 ), .Z(\UART_RX/RX_MVF/n22 ) );
  notech_ao3 \UART_RX/RX_MVF/U15  ( .A(\UART_RX/RX_MVF/iCounter[1] ), .B(
        \UART_RX/RX_MVF/iCounter[0] ), .C(\UART_RX/RX_MVF/n10 ), .Z(
        \UART_RX/RX_MVF/n7 ) );
  notech_nor2 \UART_RX/RX_MVF/U14  ( .A(\UART_RX/RX_MVF/n10 ), .B(
        \UART_RX/RX_MVF/iCounter[0] ), .Z(\UART_RX/RX_MVF/n11 ) );
  notech_or2 \UART_RX/RX_MVF/U13  ( .A(\UART_RX/RX_MVF/n11 ), .B(
        \UART_RX/RX_MVF/n2 ), .Z(\UART_RX/RX_MVF/n6 ) );
  notech_nor2 \UART_RX/RX_MVF/U12  ( .A(\UART_RX/RX_MVF/n10 ), .B(
        \UART_RX/RX_MVF/iCounter[1] ), .Z(\UART_RX/RX_MVF/n9 ) );
  notech_or2 \UART_RX/RX_MVF/U11  ( .A(\UART_RX/RX_MVF/n6 ), .B(
        \UART_RX/RX_MVF/n9 ), .Z(\UART_RX/RX_MVF/n8 ) );
  notech_mux2 \UART_RX/RX_MVF/U10  ( .A(\UART_RX/RX_MVF/n7 ), .B(
        \UART_RX/RX_MVF/n8 ), .S(\UART_RX/RX_MVF/iCounter[2] ), .Z(
        \UART_RX/RX_MVF/n23 ) );
  notech_and2 \UART_RX/RX_MVF/U9  ( .A(\UART_RX/RX_MVF/n1 ), .B(
        \UART_RX/RX_MVF/iCounter[0] ), .Z(\UART_RX/RX_MVF/n5 ) );
  notech_mux2 \UART_RX/RX_MVF/U8  ( .A(\UART_RX/RX_MVF/n5 ), .B(
        \UART_RX/RX_MVF/n6 ), .S(\UART_RX/RX_MVF/iCounter[1] ), .Z(
        \UART_RX/RX_MVF/n24 ) );
  notech_mux2 \UART_RX/RX_MVF/U7  ( .A(\UART_RX/RX_MVF/n1 ), .B(
        \UART_RX/RX_MVF/n2 ), .S(\UART_RX/RX_MVF/iCounter[0] ), .Z(
        \UART_RX/RX_MVF/n26 ) );
  notech_and3 \UART_RX/RX_MVF/U3  ( .A(iSIN), .B(\UART_RX/RX_MVF/n16 ), .C(
        iRCLK), .Z(\UART_RX/RX_MVF/n15 ) );
  notech_reg \UART_RX/RX_MVF/iQ_reg  ( .D(\UART_RX/RX_MVF/n21 ), .CP(CLK), 
        .CD(\UART_IS_CTS/n1 ), .Q(\UART_RX/iFSIN ) );
  notech_reg \UART_RX/RX_MVF/iCounter_reg[1]  ( .D(\UART_RX/RX_MVF/n24 ), .CP(
        CLK), .CD(\UART_IF_CTS/n8 ), .Q(\UART_RX/RX_MVF/iCounter[1] ) );
  notech_reg \UART_RX/RX_MVF/iCounter_reg[2]  ( .D(\UART_RX/RX_MVF/n23 ), .CP(
        CLK), .CD(\UART_IS_SIN/n1 ), .Q(\UART_RX/RX_MVF/iCounter[2] ) );
  notech_reg \UART_RX/RX_MVF/iCounter_reg[3]  ( .D(\UART_RX/RX_MVF/n22 ), .CP(
        CLK), .CD(\UART_IS_SIN/n1 ), .Q(\UART_RX/RX_MVF/iCounter[3] ) );
  notech_reg \UART_RX/RX_MVF/iCounter_reg[0]  ( .D(\UART_RX/RX_MVF/n26 ), .CP(
        CLK), .CD(\UART_IF_DSR/n8 ), .Q(\UART_RX/RX_MVF/iCounter[0] ) );
  notech_nor2 \UART_RX/RX_IFSB/U25  ( .A(\UART_RX/RX_IFSB/iCount[0] ), .B(
        \UART_RX/RX_IFSB/iCount[1] ), .Z(\UART_RX/RX_IFSB/n18 ) );
  notech_inv \UART_RX/RX_IFSB/U24  ( .A(\UART_RX/RX_IFSB/n18 ), .Z(
        \UART_RX/RX_IFSB/n15 ) );
  notech_and2 \UART_RX/RX_IFSB/U23  ( .A(\UART_RX/iFStopBit ), .B(
        \UART_RX/RX_IFSB/n15 ), .Z(\UART_RX/RX_IFSB/n17 ) );
  notech_and2 \UART_RX/RX_IFSB/U22  ( .A(\UART_RX/RX_IFSB/n18 ), .B(
        \UART_RX/RX_IFSB/iCount[2] ), .Z(\UART_RX/RX_IFSB/n16 ) );
  notech_or2 \UART_RX/RX_IFSB/U21  ( .A(\UART_RX/RX_IFSB/n17 ), .B(
        \UART_RX/RX_IFSB/n16 ), .Z(\UART_RX/RX_IFSB/n30 ) );
  notech_inv \UART_RX/RX_IFSB/U20  ( .A(iSIN), .Z(\UART_RX/RX_IFSB/n8 ) );
  notech_nor2 \UART_RX/RX_IFSB/U19  ( .A(\UART_RX/RX_IFSB/n16 ), .B(
        \UART_RX/RX_IFSB/n8 ), .Z(\UART_RX/RX_IFSB/n11 ) );
  notech_or2 \UART_RX/RX_IFSB/U18  ( .A(\UART_RX/RX_IFSB/n15 ), .B(
        \UART_RX/RX_IFSB/iCount[2] ), .Z(\UART_RX/RX_IFSB/n14 ) );
  notech_and2 \UART_RX/RX_IFSB/U17  ( .A(\UART_RX/RX_IFSB/n14 ), .B(
        \UART_RX/RX_IFSB/n8 ), .Z(\UART_RX/RX_IFSB/n13 ) );
  notech_or2 \UART_RX/RX_IFSB/U16  ( .A(\UART_RX/RX_IFSB/n11 ), .B(
        \UART_RX/RX_IFSB/n13 ), .Z(\UART_RX/RX_IFSB/n12 ) );
  notech_nand2 \UART_RX/RX_IFSB/U15  ( .A(\UART_RX/RX_IFSB/n12 ), .B(iRCLK), 
        .Z(\UART_RX/RX_IFSB/n2 ) );
  notech_xor2 \UART_RX/RX_IFSB/U14  ( .A(\UART_RX/RX_IFSB/iCount[0] ), .B(
        \UART_RX/RX_IFSB/n11 ), .Z(\UART_RX/RX_IFSB/n10 ) );
  notech_nor2 \UART_RX/RX_IFSB/U13  ( .A(\UART_RX/RX_IFSB/n2 ), .B(
        \UART_RX/RX_IFSB/n10 ), .Z(\UART_RX/RX_IFSB/n9 ) );
  notech_xor2 \UART_RX/RX_IFSB/U12  ( .A(\UART_RX/RX_IFSB/iCount[1] ), .B(
        \UART_RX/RX_IFSB/n9 ), .Z(\UART_RX/RX_IFSB/n31 ) );
  notech_and4 \UART_RX/RX_IFSB/U11  ( .A(\UART_RX/RX_IFSB/iCount[1] ), .B(
        \UART_RX/RX_IFSB/iCount[0] ), .C(iRCLK), .D(iSIN), .Z(
        \UART_RX/RX_IFSB/n3 ) );
  notech_inv \UART_RX/RX_IFSB/U10  ( .A(\UART_RX/RX_IFSB/iCount[1] ), .Z(
        \UART_RX/RX_IFSB/n7 ) );
  notech_nand2 \UART_RX/RX_IFSB/U9  ( .A(\UART_RX/RX_IFSB/iCount[0] ), .B(
        \UART_RX/RX_IFSB/n7 ), .Z(\UART_RX/RX_IFSB/n5 ) );
  notech_mux2 \UART_RX/RX_IFSB/U8  ( .A(\UART_RX/RX_IFSB/iCount[0] ), .B(
        \UART_RX/RX_IFSB/n7 ), .S(\UART_RX/RX_IFSB/n8 ), .Z(
        \UART_RX/RX_IFSB/n6 ) );
  notech_nand3 \UART_RX/RX_IFSB/U7  ( .A(iRCLK), .B(\UART_RX/RX_IFSB/n5 ), .C(
        \UART_RX/RX_IFSB/n6 ), .Z(\UART_RX/RX_IFSB/n4 ) );
  notech_mux2 \UART_RX/RX_IFSB/U6  ( .A(\UART_RX/RX_IFSB/n3 ), .B(
        \UART_RX/RX_IFSB/n4 ), .S(\UART_RX/RX_IFSB/iCount[2] ), .Z(
        \UART_RX/RX_IFSB/n32 ) );
  notech_xor2 \UART_RX/RX_IFSB/U5  ( .A(\UART_RX/RX_IFSB/iCount[0] ), .B(
        \UART_RX/RX_IFSB/n2 ), .Z(\UART_RX/RX_IFSB/n1 ) );
  notech_inv \UART_RX/RX_IFSB/U4  ( .A(\UART_RX/RX_IFSB/n1 ), .Z(
        \UART_RX/RX_IFSB/n33 ) );
  notech_reg \UART_RX/RX_IFSB/Q_reg  ( .D(\UART_RX/RX_IFSB/n30 ), .CP(CLK), 
        .CD(\UART_IF_DSR/n8 ), .Q(\UART_RX/iFStopBit ) );
  notech_reg \UART_RX/RX_IFSB/iCount_reg[2]  ( .D(\UART_RX/RX_IFSB/n32 ), .CP(
        CLK), .CD(\UART_IF_DSR/n8 ), .Q(\UART_RX/RX_IFSB/iCount[2] ) );
  notech_reg \UART_RX/RX_IFSB/iCount_reg[1]  ( .D(\UART_RX/RX_IFSB/n31 ), .CP(
        CLK), .CD(\UART_IS_DCD/n1 ), .Q(\UART_RX/RX_IFSB/iCount[1] ) );
  notech_reg \UART_RX/RX_IFSB/iCount_reg[0]  ( .D(\UART_RX/RX_IFSB/n33 ), .CP(
        CLK), .CD(\UART_IS_SIN/n1 ), .Q(\UART_RX/RX_IFSB/iCount[0] ) );
  notech_inv \r108/U1  ( .A(\U3/U1/Z_0 ), .Z(\r108/n1 ) );
  notech_fa2 \r108/U1_0  ( .A(iFECounter[0]), .B(\U3/U1/Z_0 ), .CI(\r108/n1 ), 
        .CO(\r108/carry [1]) );
  notech_fa2 \r108/U1_1  ( .A(iFECounter[1]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [1]), .CO(\r108/carry [2]), .Z(N130) );
  notech_fa2 \r108/U1_2  ( .A(iFECounter[2]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [2]), .CO(\r108/carry [3]), .Z(N131) );
  notech_fa2 \r108/U1_3  ( .A(iFECounter[3]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [3]), .CO(\r108/carry [4]), .Z(N132) );
  notech_fa2 \r108/U1_4  ( .A(iFECounter[4]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [4]), .CO(\r108/carry [5]), .Z(N133) );
  notech_fa2 \r108/U1_5  ( .A(iFECounter[5]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [5]), .CO(\r108/carry [6]), .Z(N134) );
  notech_fa2 \r108/U1_6  ( .A(iFECounter[6]), .B(\U3/U1/Z_0 ), .CI(
        \r108/carry [6]), .Z(N135) );
  notech_nand2 U458 ( .A(\UART_RX/n62 ), .B(\UART_RX/iBaudCount[3] ), .Z(n680)
         );
  notech_nand2 U461 ( .A(\UART_RX/RX_BRC/Q[1] ), .B(\UART_RX/RX_BRC/Q[0] ), 
        .Z(n681) );
  notech_nand2 U471 ( .A(\UART_BG16/n35 ), .B(n686), .Z(n682) );
  notech_nand2 U545 ( .A(N154), .B(\UART_ED_CTS/n1 ), .Z(n683) );
  notech_nand2 U546 ( .A(N155), .B(\UART_ED_DSR/n1 ), .Z(n684) );
  notech_nand2 U637 ( .A(N157), .B(\UART_ED_DCD/n1 ), .Z(n685) );
  notech_inv U672 ( .A(BAUDCE), .Z(n686) );
  notech_nand2 U756 ( .A(\UART_RX/n61 ), .B(n687), .Z(\UART_RX/RX_BRC/n6 ) );
  notech_inv U790 ( .A(iRCLK), .Z(n687) );
  notech_and2 U807 ( .A(\UART_RX/n61 ), .B(\UART_RX/n42 ), .Z(
        \UART_RX/RX_BRC/n23 ) );
  notech_xor2 U835 ( .A(n688), .B(\UART_RX/RX_BRC/n5 ), .Z(\UART_RX/RX_BRC/n9 ) );
  notech_inv U836 ( .A(\UART_RX/RX_BRC/Q[0] ), .Z(n688) );
  notech_xor2 U837 ( .A(n681), .B(\UART_RX/RX_BRC/Q[2] ), .Z(
        \UART_RX/RX_BRC/n13 ) );
  notech_xor2 U838 ( .A(n689), .B(\UART_RX/RX_BRC/n17 ), .Z(
        \UART_RX/RX_BRC/n18 ) );
  notech_inv U839 ( .A(\UART_RX/RX_BRC/n21 ), .Z(n689) );
  notech_nor2 U840 ( .A(\UART_RX/RX_BRC/n21 ), .B(\UART_RX/RX_BRC/n17 ), .Z(
        \UART_RX/RX_BRC/n22 ) );
  notech_or2 U841 ( .A(\UART_RX/RX_BRC/n12 ), .B(n681), .Z(
        \UART_RX/RX_BRC/n21 ) );
  notech_and2 U842 ( .A(\UART_RX/RX_MVF/n16 ), .B(\UART_RX/n43 ), .Z(
        \UART_RX/RX_MVF/n17 ) );
  notech_nand2 U843 ( .A(BAUDCE), .B(\UART_BG16/n35 ), .Z(\UART_BG16/n2 ) );
endmodule

