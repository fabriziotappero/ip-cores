package vcomponents is
end;
