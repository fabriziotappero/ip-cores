`timescale 1 ns/ 1 ps
package wb_ahb_pkg;
import global::*;
	`include "../avm_svtb/wb_ahb_stim_gen.svh"
	`include "../avm_svtb/wb_ahb_driver.svh"
	`include "../avm_svtb/wb_ahb_responder.svh"
	`include "../avm_svtb/wb_ahb_monitor.svh"
	`include "../avm_svtb/wb_ahb_scoreboard.svh"
	`include "../avm_svtb/wb_ahb_coverage.svh"
	`include "../avm_svtb/wb_ahb_env.svh"
endpackage

