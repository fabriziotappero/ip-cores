--------------------------------------------------------------------------------
--                                                                            --
--                          V H D L    F I L E                                --
--                          COPYRIGHT (C) 2006                                --
--                                                                            --
--------------------------------------------------------------------------------
--
-- Title       : DCT
-- Design      : MDCT Core
-- Author      : Michal Krepa
--
--------------------------------------------------------------------------------
--
-- File        : DCT_TROM.VHD
-- Created     : Sun Aug 27 18:09 2006
--
--------------------------------------------------------------------------------
--
--  Description : ROM for DCT quantizer matrix
--
--------------------------------------------------------------------------------

library IEEE; 
  use IEEE.STD_LOGIC_1164.all; 
  use ieee.numeric_std.all; 

entity DCT_TROM is 
  generic 
    ( 
      ROMADDR_W     : INTEGER := 9;
      ROMDATA_W     : INTEGER := 8
    );
  port( 
       addr         : in  STD_LOGIC_VECTOR(ROMADDR_W-1 downto 0);
       clk          : in  STD_LOGIC;  
       
       datao        : out STD_LOGIC_VECTOR(ROMDATA_W-1 downto 0) 
  );          
  
end DCT_TROM; 

architecture RTL of DCT_TROM is  

  type DCT_TROM_TYPE is array (0 to 2**ROMADDR_W-1) 
            of INTEGER;
  
  constant rom : DCT_TROM_TYPE := 
  -- (
  -- 16,11,10,16,24,40,51,61,
  -- 12,12,14,19,26,58,60,55,
  -- 14,13,16,24,40,57,69,56,
  -- 14,17,22,29,51,87,80,62,
  -- 18,22,37,56,68,109,103,77,
  -- 24,35,55,64,81,104,113,92,
  -- 49,64,78,87,103,121,120,101,
  -- 72,92,95,98,112,100,103,99);
                          (
    -280,    48,   -20,    16,   -26,    46,   -42,    27,
      45,    12,   -34,   -31,    11,    -1,    16,   -44,
      -5,   -63,   -34,    36,    24,   -27,     6,     1,
     -12,    12,    -8,    34,     5,     2,   -12,     5,
      22,   -18,    15,     9,    12,    -5,     1,   -11,
       1,    10,     6,    12,   -15,   -11,    -5,   -10,
       5,   -16,    -4,    10,    -1,   -11,    -5,   -11,
      -9,    11,     5,    -3,   -14,     4,     0,     0,
    -213,  -110,   -78,    38,    32,     2,    -1,    -9,
      28,    62,    -7,    -7,    22,   -11,     5,     7,
      85,   -21,    33,   -28,   -37,    36,   -11,     5,
     -34,   -18,     2,   -24,     8,   -12,   -11,    -8,
     -13,     8,    39,   -63,    27,     0,     1,    -4,
     -32,    -4,    -8,    24,   -22,    11,    20,    -4,
     -12,     8,    43,    41,   -16,   -12,     4,   -10,
     -11,    14,    15,     7,   -11,     9,   -32,     0,
    -225,    10,    25,    18,   -30,    18,   -14,     7,
      44,   -13,   -93,    -7,    20,    -7,     5,   -11,
     -88,   -53,     6,    36,     2,     1,    22,     2,
     -46,   -10,    17,    23,    16,    32,    -7,     8,
      66,    46,   -10,    -3,   -17,     4,    -5,    -5,
     -51,   -18,    -9,     6,    37,    15,    23,    -4,
     -21,    22,    44,    49,    25,    21,     1,   -12,
      25,    12,    -5,    -2,   -19,    -8,   -15,     0,
     390,   -97,   -41,   -15,    20,     6,     0,    12,
       4,   -62,    21,    -5,   -31,    -7,    -3,   -20,
    -352,    44,    27,    36,    35,     6,     5,    10,
      33,    48,    48,    14,    -8,    14,    10,    -9,
     -95,   108,     5,     1,   -11,   -23,   -20,     1,
      54,    -7,   -43,   -32,   -15,     3,     9,     3,
     -42,    57,   -32,   -19,    -4,     6,     5,    -3,
      23,   -31,   -22,    -1,    19,    24,    22,     1,
     -14,   148,    70,    67,    54,    30,     2,   -10,
      76,    20,    20,   -39,    14,   -10,    -8,   -11,
     -86,   -65,   -15,   -33,   -33,   -38,    -2,    10,
      61,    20,    50,    18,   -15,   -25,   -23,     2,
      11,    -3,    12,    12,    15,     8,   -18,    -5,
     -13,   -14,   -13,    16,    34,    15,   -22,   -18,
      -8,   -13,    -3,    11,    19,    26,     9,    -5,
       1,     1,     2,    -9,   -11,     2,     7,     0,
    -317,    -9,    63,    17,    10,   -26,     1,   -11,
     159,   -41,   -29,    42,    -3,    21,    11,     1,
      -6,   -13,   -18,     9,   -19,     5,    15,     7,
      -8,    -9,   -11,    16,    -4,    -1,   -12,    -3,
       1,    15,    -1,     3,   -13,    -8,     5,    -1,
      -9,     3,     2,     5,     7,    -6,    12,   -11,
      -3,     1,    -6,     1,    -5,    -4,     9,     6,
       3,     7,     7,     3,    -3,    -5,    -2,     0,


     -404,   148,    70,    67,    54,    30,     2,   -10,
      76,    20,    20,   -39,    14,   -10,    -8,   -11,
     -86,   -65,   -15,   -33,   -33,   -38,    -2,    10,
      61,    20,    50,    18,   -15,   -25,   -23,     2,
      11,    -3,    12,    12,    15,     8,   -18,    -5,
     -13,   -14,   -13,    16,    34,    15,   -22,   -18,
      -8,   -13,    -3,    11,    19,    26,     9,    -5,
       1,     1,     2,    -9,   -11,     2,     7,     0,
       -404,   148,    70,    67,    54,    30,     2,   -10,
      76,    20,    20,   -39,    14,   -10,    -8,   -11,
     -86,   -65,   -15,   -33,   -33,   -38,    -2,    10,
      61,    20,    50,    18,   -15,   -25,   -23,     2,
      11,    -3,    12,    12,    15,     8,   -18,    -5,
     -13,   -14,   -13,    16,    34,    15,   -22,   -18,
      -8,   -13,    -3,    11,    19,    26,     9,    -5,
       1,     1,     2,    -9,   -11,     2,     7,     0
       


                          );
            
 

  signal addr_reg : STD_LOGIC_VECTOR(ROMADDR_W-1 downto 0);
begin   
  
  datao <= STD_LOGIC_VECTOR(TO_SIGNED( rom( TO_INTEGER(UNSIGNED(addr_reg)) ), ROMDATA_W)); 
  
  process(clk)
  begin
   if clk = '1' and clk'event then
     addr_reg <= addr;
   end if;
  end process;
      
end RTL;    
