-- SPI_OC enable 
  constant CFG_SPI_OC  : integer := CONFIG_SPI_OC_ENABLE;

